VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO clkgate
  CLASS BLOCK ;
  FOREIGN clkgate ;
  ORIGIN 0.000 0.000 ;
  SIZE 60.000 BY 60.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 29.680 0.000 30.240 4.000 ;
    END
  END clk
  PIN gate
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 29.680 4.000 30.240 ;
    END
  END gate
  PIN gclk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 29.680 56.000 30.240 60.000 ;
    END
  END gclk
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 11.730 15.380 13.330 43.420 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 23.350 15.380 24.950 43.420 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 34.970 15.380 36.570 43.420 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 46.590 15.380 48.190 43.420 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 17.540 15.380 19.140 43.420 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 29.160 15.380 30.760 43.420 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 40.780 15.380 42.380 43.420 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 52.400 15.380 54.000 43.420 ;
    END
  END vss
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 54.000 43.420 ;
      LAYER Metal2 ;
        RECT 9.100 55.700 29.380 56.000 ;
        RECT 30.540 55.700 53.860 56.000 ;
        RECT 9.100 4.300 53.860 55.700 ;
        RECT 9.100 4.000 29.380 4.300 ;
        RECT 30.540 4.000 53.860 4.300 ;
      LAYER Metal3 ;
        RECT 4.000 30.540 53.910 43.260 ;
        RECT 4.300 29.380 53.910 30.540 ;
        RECT 4.000 15.540 53.910 29.380 ;
  END
END clkgate
END LIBRARY

