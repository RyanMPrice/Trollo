// This is the unpowered netlist.
module user_proj_example (wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    io_in,
    io_oeb,
    io_out,
    irq,
    la_data_in,
    la_data_out,
    la_oenb,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o,
    wbs_sel_i);
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;
 output [2:0] irq;
 input [63:0] la_data_in;
 output [63:0] la_data_out;
 input [63:0] la_oenb;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;
 input [3:0] wbs_sel_i;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire \dsynth.csTable.address[0] ;
 wire \dsynth.csTable.address[1] ;
 wire \dsynth.csTable.address[2] ;
 wire \dsynth.csTable.address[3] ;
 wire \dsynth.csTable.address[4] ;
 wire \dsynth.csTable.address[5] ;
 wire \dsynth.csTable.address[6] ;
 wire \dsynth.csTable.address[7] ;
 wire \dsynth.freeRunCntr[0] ;
 wire \dsynth.freeRunCntr[10] ;
 wire \dsynth.freeRunCntr[11] ;
 wire \dsynth.freeRunCntr[12] ;
 wire \dsynth.freeRunCntr[13] ;
 wire \dsynth.freeRunCntr[14] ;
 wire \dsynth.freeRunCntr[15] ;
 wire \dsynth.freeRunCntr[16] ;
 wire \dsynth.freeRunCntr[17] ;
 wire \dsynth.freeRunCntr[1] ;
 wire \dsynth.freeRunCntr[26] ;
 wire \dsynth.freeRunCntr[27] ;
 wire \dsynth.freeRunCntr[28] ;
 wire \dsynth.freeRunCntr[29] ;
 wire \dsynth.freeRunCntr[2] ;
 wire \dsynth.freeRunCntr[30] ;
 wire \dsynth.freeRunCntr[31] ;
 wire \dsynth.freeRunCntr[32] ;
 wire \dsynth.freeRunCntr[3] ;
 wire \dsynth.freeRunCntr[4] ;
 wire \dsynth.freeRunCntr[5] ;
 wire \dsynth.freeRunCntr[6] ;
 wire \dsynth.freeRunCntr[7] ;
 wire \dsynth.freeRunCntr[8] ;
 wire \dsynth.freeRunCntr[9] ;
 wire net196;
 wire net64;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net197;
 wire net70;
 wire net207;
 wire net208;
 wire net71;
 wire net72;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net73;
 wire net198;
 wire net74;
 wire net75;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net61;
 wire net62;
 wire net63;
 wire net76;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net77;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net78;
 wire net219;
 wire net220;
 wire net93;
 wire net94;
 wire net95;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net100;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net101;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net102;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net103;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net104;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire \tgate.clkp ;
 wire \tmux.clkapa ;
 wire \tmux.clkbpb ;
 wire \tmux.clkpaa ;
 wire \tmux.clkpab ;
 wire \tmux.clkpba ;
 wire \tmux.clkpbb ;
 wire net163;
 wire net164;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net165;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net166;
 wire net194;
 wire net195;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;

 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1920_ (.I(\dsynth.freeRunCntr[16] ),
    .ZN(_0063_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1921_ (.I(\dsynth.csTable.address[6] ),
    .Z(_0074_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1922_ (.I(_0074_),
    .Z(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1923_ (.I(\dsynth.csTable.address[7] ),
    .ZN(_0096_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1924_ (.A1(_0085_),
    .A2(_0096_),
    .Z(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1925_ (.I(_0107_),
    .Z(_0118_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1926_ (.I(_0118_),
    .Z(_0129_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1927_ (.A1(_0063_),
    .A2(_0129_),
    .ZN(_0140_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1928_ (.I(\dsynth.csTable.address[6] ),
    .Z(_0151_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1929_ (.A1(_0151_),
    .A2(\dsynth.csTable.address[4] ),
    .ZN(_0162_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1930_ (.I(_0162_),
    .Z(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1931_ (.I(_0173_),
    .Z(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1932_ (.I(_0184_),
    .Z(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1933_ (.I(_0195_),
    .Z(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1934_ (.A1(_0151_),
    .A2(\dsynth.csTable.address[2] ),
    .ZN(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1935_ (.I(_0217_),
    .Z(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1936_ (.I(_0228_),
    .Z(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1937_ (.I(\dsynth.csTable.address[0] ),
    .Z(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1938_ (.A1(_0151_),
    .A2(_0250_),
    .ZN(_0261_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1939_ (.I(_0261_),
    .Z(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1940_ (.I(_0272_),
    .Z(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1941_ (.A1(_0239_),
    .A2(_0283_),
    .ZN(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1942_ (.I(\dsynth.csTable.address[6] ),
    .Z(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1943_ (.A1(_0305_),
    .A2(\dsynth.csTable.address[1] ),
    .ZN(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1944_ (.I(_0316_),
    .Z(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1945_ (.I(_0217_),
    .Z(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1946_ (.I(\dsynth.csTable.address[3] ),
    .Z(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1947_ (.A1(_0151_),
    .A2(_0349_),
    .ZN(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1948_ (.I(_0360_),
    .Z(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1949_ (.A1(_0327_),
    .A2(_0338_),
    .B(_0371_),
    .ZN(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1950_ (.I(_0382_),
    .Z(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1951_ (.A1(_0294_),
    .A2(_0393_),
    .ZN(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1952_ (.A1(_0206_),
    .A2(_0404_),
    .ZN(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1953_ (.A1(_0305_),
    .A2(\dsynth.csTable.address[3] ),
    .Z(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1954_ (.I(_0426_),
    .Z(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1955_ (.I(_0437_),
    .Z(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1956_ (.I(_0448_),
    .Z(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1957_ (.I(_0459_),
    .Z(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1958_ (.I(_0316_),
    .Z(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1959_ (.I(_0481_),
    .Z(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1960_ (.I(_0492_),
    .Z(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1961_ (.I(_0338_),
    .Z(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1962_ (.A1(_0503_),
    .A2(_0514_),
    .ZN(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1963_ (.I(\dsynth.csTable.address[5] ),
    .Z(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1964_ (.A1(_0536_),
    .A2(_0074_),
    .Z(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1965_ (.I(_0547_),
    .Z(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1966_ (.I(_0558_),
    .Z(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1967_ (.I(_0569_),
    .Z(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1968_ (.A1(_0470_),
    .A2(_0525_),
    .B(_0580_),
    .ZN(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1969_ (.A1(\dsynth.csTable.address[6] ),
    .A2(\dsynth.csTable.address[1] ),
    .Z(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1970_ (.I(_0602_),
    .Z(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1971_ (.I(_0613_),
    .Z(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1972_ (.A1(_0305_),
    .A2(\dsynth.csTable.address[2] ),
    .Z(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1973_ (.I(_0635_),
    .Z(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1974_ (.I(_0646_),
    .Z(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1975_ (.A1(_0624_),
    .A2(_0657_),
    .ZN(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1976_ (.I(_0360_),
    .Z(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1977_ (.I(_0679_),
    .Z(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1978_ (.I(_0690_),
    .Z(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1979_ (.I(_0646_),
    .Z(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1980_ (.A1(_0305_),
    .A2(\dsynth.csTable.address[0] ),
    .Z(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1981_ (.I(_0723_),
    .Z(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1982_ (.I(_0734_),
    .Z(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1983_ (.A1(_0712_),
    .A2(_0745_),
    .ZN(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1984_ (.I(_0756_),
    .Z(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1985_ (.I(_0173_),
    .Z(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1986_ (.I(_0778_),
    .Z(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _1987_ (.A1(_0668_),
    .A2(_0701_),
    .A3(_0767_),
    .B(_0789_),
    .ZN(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1988_ (.I(_0437_),
    .Z(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1989_ (.I(_0217_),
    .Z(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1990_ (.A1(_0481_),
    .A2(_0272_),
    .B(_0822_),
    .ZN(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1991_ (.I(_0602_),
    .Z(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1992_ (.I(_0635_),
    .Z(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1993_ (.I(_0426_),
    .Z(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1994_ (.A1(_0844_),
    .A2(_0855_),
    .B(_0866_),
    .ZN(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1995_ (.I(_0316_),
    .Z(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1996_ (.I(_0261_),
    .Z(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1997_ (.A1(_0888_),
    .A2(_0338_),
    .A3(_0899_),
    .ZN(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _1998_ (.A1(_0811_),
    .A2(_0833_),
    .B1(_0877_),
    .B2(_0909_),
    .ZN(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1999_ (.I(_0173_),
    .Z(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2000_ (.I(_0931_),
    .Z(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2001_ (.A1(_0800_),
    .A2(_0404_),
    .B1(_0920_),
    .B2(_0942_),
    .ZN(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2002_ (.I(_0558_),
    .Z(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2003_ (.I(_0958_),
    .Z(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2004_ (.A1(_0415_),
    .A2(_0591_),
    .B1(_0952_),
    .B2(_0963_),
    .ZN(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2005_ (.A1(_0118_),
    .A2(_0971_),
    .Z(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2006_ (.I(_0981_),
    .Z(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2007_ (.I(\dsynth.csTable.address[7] ),
    .Z(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2008_ (.A1(_0085_),
    .A2(_1001_),
    .Z(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2009_ (.I(_1010_),
    .Z(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2010_ (.I(_1020_),
    .Z(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2011_ (.A1(_0074_),
    .A2(\dsynth.csTable.address[4] ),
    .Z(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2012_ (.I(_1040_),
    .Z(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2013_ (.I(_1049_),
    .Z(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2014_ (.I(_1059_),
    .Z(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2015_ (.A1(_1069_),
    .A2(_0393_),
    .ZN(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2016_ (.A1(_0800_),
    .A2(_1078_),
    .B(_0591_),
    .ZN(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _2017_ (.A1(_1030_),
    .A2(_1087_),
    .Z(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2018_ (.I(\dsynth.freeRunCntr[14] ),
    .Z(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2019_ (.A1(\dsynth.freeRunCntr[13] ),
    .A2(_0991_),
    .B1(_1095_),
    .B2(_1103_),
    .ZN(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2020_ (.I(\dsynth.freeRunCntr[15] ),
    .Z(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2021_ (.I(_1118_),
    .Z(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2022_ (.I(_0107_),
    .Z(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2023_ (.I(_0580_),
    .Z(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2024_ (.A1(_1125_),
    .A2(_0800_),
    .ZN(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2025_ (.A1(_1124_),
    .A2(_1126_),
    .Z(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2026_ (.I(_1127_),
    .Z(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2027_ (.I(_1128_),
    .Z(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2028_ (.A1(_1123_),
    .A2(_1129_),
    .B1(_1095_),
    .B2(_1103_),
    .ZN(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2029_ (.I(\dsynth.freeRunCntr[16] ),
    .Z(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2030_ (.I(_1030_),
    .Z(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2031_ (.A1(_1131_),
    .A2(_1132_),
    .B1(_1129_),
    .B2(_1123_),
    .ZN(_1133_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2032_ (.A1(_1110_),
    .A2(_1130_),
    .B(_1133_),
    .ZN(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2033_ (.I(\dsynth.freeRunCntr[13] ),
    .ZN(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2034_ (.I(_1135_),
    .Z(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2035_ (.A1(_1010_),
    .A2(_0971_),
    .Z(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2036_ (.A1(_1136_),
    .A2(_1137_),
    .B(_1130_),
    .ZN(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _2037_ (.A1(_0140_),
    .A2(_1133_),
    .A3(_1110_),
    .A4(_1138_),
    .Z(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2038_ (.I(_0613_),
    .Z(_1140_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2039_ (.I(_1140_),
    .Z(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2040_ (.I(_0712_),
    .Z(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2041_ (.A1(_1141_),
    .A2(_1142_),
    .ZN(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2042_ (.I(\dsynth.csTable.address[1] ),
    .Z(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2043_ (.I(_0250_),
    .Z(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2044_ (.A1(_1144_),
    .A2(_1145_),
    .Z(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2045_ (.A1(_0239_),
    .A2(_1146_),
    .B(_0690_),
    .ZN(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2046_ (.I(_1147_),
    .Z(_1148_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2047_ (.A1(_0481_),
    .A2(_0646_),
    .B(_0426_),
    .ZN(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2048_ (.I(_1149_),
    .Z(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2049_ (.A1(_1144_),
    .A2(_0250_),
    .ZN(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2050_ (.A1(_0338_),
    .A2(_1151_),
    .ZN(_1152_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2051_ (.A1(_0558_),
    .A2(_1049_),
    .ZN(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2052_ (.A1(_1143_),
    .A2(_1148_),
    .B1(_1150_),
    .B2(_1152_),
    .C(_1153_),
    .ZN(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2053_ (.I(_0899_),
    .Z(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2054_ (.A1(_0514_),
    .A2(_1155_),
    .B(_0690_),
    .ZN(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2055_ (.I(\dsynth.csTable.address[2] ),
    .Z(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2056_ (.A1(_1144_),
    .A2(_1157_),
    .Z(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2057_ (.I(_1158_),
    .Z(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2058_ (.A1(_0569_),
    .A2(_0931_),
    .ZN(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2059_ (.I(_1160_),
    .Z(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2060_ (.A1(_0822_),
    .A2(_0734_),
    .ZN(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2061_ (.I(_1162_),
    .Z(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2062_ (.I(_0855_),
    .Z(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2063_ (.A1(_0492_),
    .A2(_0283_),
    .B(_1164_),
    .ZN(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2064_ (.I(_0811_),
    .Z(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2065_ (.I(_1166_),
    .Z(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2066_ (.A1(_0503_),
    .A2(_1163_),
    .B(_1165_),
    .C(_1167_),
    .ZN(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2067_ (.A1(_1156_),
    .A2(_1159_),
    .B(_1161_),
    .C(_1168_),
    .ZN(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2068_ (.I(_0294_),
    .Z(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2069_ (.I(_0327_),
    .Z(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2070_ (.I(_0371_),
    .Z(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2071_ (.A1(_1171_),
    .A2(_1172_),
    .ZN(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2072_ (.A1(_1170_),
    .A2(_1173_),
    .ZN(_1174_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2073_ (.I(_1164_),
    .Z(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2074_ (.I(_0723_),
    .Z(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2075_ (.I(_1176_),
    .Z(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2076_ (.A1(_1175_),
    .A2(_1177_),
    .ZN(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2077_ (.I(_0877_),
    .Z(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2078_ (.I(_0778_),
    .Z(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2079_ (.A1(_1178_),
    .A2(_1179_),
    .B1(_1159_),
    .B2(_1167_),
    .C(_1180_),
    .ZN(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2080_ (.A1(_0206_),
    .A2(_1174_),
    .B(_1181_),
    .C(_0963_),
    .ZN(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2081_ (.A1(_1154_),
    .A2(_1169_),
    .A3(_1182_),
    .ZN(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2082_ (.A1(_1124_),
    .A2(_1183_),
    .Z(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2083_ (.I(_1184_),
    .Z(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2084_ (.I(_1185_),
    .Z(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2085_ (.A1(\dsynth.freeRunCntr[12] ),
    .A2(_1186_),
    .ZN(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2086_ (.I(_1010_),
    .Z(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2087_ (.A1(\dsynth.csTable.address[5] ),
    .A2(_0074_),
    .ZN(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2088_ (.I(_1189_),
    .Z(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2089_ (.I(_1190_),
    .Z(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2090_ (.I(_1049_),
    .Z(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2091_ (.A1(_1191_),
    .A2(_1192_),
    .ZN(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2092_ (.I(_1193_),
    .Z(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2093_ (.I(_0701_),
    .Z(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2094_ (.I(_0723_),
    .Z(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2095_ (.A1(\dsynth.csTable.address[1] ),
    .A2(\dsynth.csTable.address[2] ),
    .ZN(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2096_ (.A1(_1196_),
    .A2(_1197_),
    .ZN(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2097_ (.I(_1198_),
    .Z(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2098_ (.I(_1151_),
    .Z(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2099_ (.I(_1200_),
    .Z(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2100_ (.I(_0393_),
    .Z(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2101_ (.A1(_1195_),
    .A2(_1170_),
    .A3(_1199_),
    .B1(_1201_),
    .B2(_1202_),
    .ZN(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2102_ (.I(_0503_),
    .Z(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2103_ (.A1(_0327_),
    .A2(_0272_),
    .B(_0679_),
    .ZN(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2104_ (.I(_1192_),
    .Z(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2105_ (.I(_1206_),
    .Z(_1207_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _2106_ (.A1(_1204_),
    .A2(_1195_),
    .B1(_1199_),
    .B2(_1205_),
    .C(_1207_),
    .ZN(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2107_ (.A1(_0250_),
    .A2(_1157_),
    .Z(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2108_ (.I(_1209_),
    .Z(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2109_ (.I0(_0657_),
    .I1(_1210_),
    .S(_0844_),
    .Z(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2110_ (.I(_1059_),
    .Z(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2111_ (.I(_0371_),
    .Z(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2112_ (.I(_1213_),
    .Z(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2113_ (.A1(_1212_),
    .A2(_1214_),
    .ZN(_1215_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2114_ (.A1(_1211_),
    .A2(_1215_),
    .B(_0963_),
    .ZN(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2115_ (.I(_1191_),
    .Z(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2116_ (.I(_1217_),
    .Z(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2117_ (.I(_0844_),
    .Z(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2118_ (.I(_1219_),
    .Z(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2119_ (.I(_0239_),
    .Z(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2120_ (.A1(_1220_),
    .A2(_1221_),
    .A3(_1214_),
    .B(_1212_),
    .ZN(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2121_ (.A1(_1145_),
    .A2(_1157_),
    .ZN(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2122_ (.I(_1223_),
    .Z(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2123_ (.A1(_1218_),
    .A2(_1222_),
    .A3(_1224_),
    .ZN(_1225_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _2124_ (.A1(_1194_),
    .A2(_1203_),
    .B1(_1208_),
    .B2(_1216_),
    .C(_1225_),
    .ZN(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2125_ (.A1(_1188_),
    .A2(_1226_),
    .Z(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2126_ (.I(_1227_),
    .Z(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2127_ (.I(_1228_),
    .Z(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2128_ (.I(\dsynth.freeRunCntr[11] ),
    .Z(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2129_ (.A1(\dsynth.freeRunCntr[12] ),
    .A2(_1186_),
    .B1(_1229_),
    .B2(_1230_),
    .ZN(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2130_ (.I(_1230_),
    .Z(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2131_ (.I(\dsynth.freeRunCntr[10] ),
    .Z(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2132_ (.I(_1190_),
    .Z(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2133_ (.I(_1234_),
    .Z(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2134_ (.I(_1235_),
    .Z(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2135_ (.I(_0657_),
    .Z(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2136_ (.I(_1237_),
    .Z(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2137_ (.I(_0866_),
    .Z(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2138_ (.A1(_1239_),
    .A2(_1146_),
    .ZN(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2139_ (.A1(_1238_),
    .A2(_1240_),
    .B(_1069_),
    .ZN(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2140_ (.I(_0899_),
    .Z(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2141_ (.I(_1242_),
    .Z(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2142_ (.A1(_0503_),
    .A2(_1175_),
    .ZN(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2143_ (.I(_0624_),
    .Z(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2144_ (.I(_0283_),
    .Z(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2145_ (.A1(_1245_),
    .A2(_1246_),
    .ZN(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2146_ (.A1(_1243_),
    .A2(_1244_),
    .B1(_1247_),
    .B2(_0470_),
    .ZN(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2147_ (.A1(_1241_),
    .A2(_1248_),
    .Z(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2148_ (.A1(_1242_),
    .A2(_1158_),
    .ZN(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2149_ (.A1(_0613_),
    .A2(_0734_),
    .B(_0360_),
    .ZN(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2150_ (.I(_1251_),
    .Z(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2151_ (.A1(_1219_),
    .A2(_1166_),
    .B(_1192_),
    .ZN(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2152_ (.A1(_1250_),
    .A2(_1252_),
    .B(_1253_),
    .ZN(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _2153_ (.A1(_1214_),
    .A2(_1243_),
    .B1(_1224_),
    .B2(_1205_),
    .C(_1069_),
    .ZN(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2154_ (.A1(_0888_),
    .A2(_0899_),
    .B(_0866_),
    .ZN(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2155_ (.I(_1256_),
    .Z(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2156_ (.I(_1257_),
    .Z(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2157_ (.I(_0569_),
    .Z(_1259_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2158_ (.A1(_0942_),
    .A2(_1258_),
    .B(_1259_),
    .ZN(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2159_ (.A1(_0942_),
    .A2(_1204_),
    .A3(_1163_),
    .ZN(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2160_ (.A1(_1255_),
    .A2(_1260_),
    .A3(_1261_),
    .ZN(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2161_ (.A1(_1236_),
    .A2(_1249_),
    .A3(_1254_),
    .B(_1262_),
    .ZN(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2162_ (.A1(_1188_),
    .A2(_1263_),
    .Z(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2163_ (.I(_1264_),
    .Z(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2164_ (.I(_1265_),
    .Z(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2165_ (.A1(_1233_),
    .A2(_1266_),
    .ZN(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2166_ (.A1(_1187_),
    .A2(_1267_),
    .ZN(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _2167_ (.A1(_1232_),
    .A2(_1229_),
    .B(_1231_),
    .C(_1268_),
    .ZN(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2168_ (.I(_1223_),
    .Z(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2169_ (.I(_0679_),
    .Z(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2170_ (.A1(_1271_),
    .A2(_1176_),
    .B(_0184_),
    .ZN(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2171_ (.A1(_1270_),
    .A2(_1257_),
    .B(_1272_),
    .ZN(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2172_ (.A1(_0613_),
    .A2(_0734_),
    .B(_0822_),
    .ZN(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2173_ (.I(_0712_),
    .Z(_1275_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2174_ (.I(_0745_),
    .Z(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2175_ (.A1(_1275_),
    .A2(_1276_),
    .B(_1172_),
    .ZN(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2176_ (.A1(_1179_),
    .A2(_1274_),
    .B1(_1250_),
    .B2(_1277_),
    .ZN(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2177_ (.A1(_1142_),
    .A2(_1155_),
    .ZN(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2178_ (.A1(_1147_),
    .A2(_1279_),
    .B(_1059_),
    .C(_1179_),
    .ZN(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2179_ (.I(_1271_),
    .Z(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2180_ (.I0(_0624_),
    .I1(_1164_),
    .S(_1176_),
    .Z(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2181_ (.A1(_1281_),
    .A2(_1282_),
    .B(_0931_),
    .ZN(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2182_ (.A1(_1280_),
    .A2(_1283_),
    .B(_1217_),
    .ZN(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _2183_ (.A1(_1235_),
    .A2(_1273_),
    .B1(_1278_),
    .B2(_1160_),
    .C(_1284_),
    .ZN(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _2184_ (.A1(_1010_),
    .A2(_1285_),
    .Z(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2185_ (.I(_1286_),
    .Z(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2186_ (.I(\dsynth.freeRunCntr[9] ),
    .Z(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2187_ (.A1(_1233_),
    .A2(_1266_),
    .B1(_1287_),
    .B2(_1288_),
    .ZN(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2188_ (.I(\dsynth.freeRunCntr[9] ),
    .Z(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2189_ (.I(_1235_),
    .Z(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2190_ (.A1(_0437_),
    .A2(_0261_),
    .A3(_1197_),
    .ZN(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2191_ (.A1(_1167_),
    .A2(_1246_),
    .ZN(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2192_ (.I(_1197_),
    .Z(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2193_ (.A1(_0888_),
    .A2(_0745_),
    .B(_1294_),
    .ZN(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2194_ (.A1(_1293_),
    .A2(_1295_),
    .B(_1212_),
    .ZN(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2195_ (.I(_1196_),
    .Z(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2196_ (.A1(_1171_),
    .A2(_1297_),
    .B(_1164_),
    .ZN(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2197_ (.A1(_0942_),
    .A2(_1298_),
    .ZN(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2198_ (.A1(_1292_),
    .A2(_1296_),
    .B1(_1299_),
    .B2(_1173_),
    .ZN(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2199_ (.I(_1165_),
    .Z(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2200_ (.A1(_1219_),
    .A2(_0514_),
    .B(_1213_),
    .ZN(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2201_ (.I(_0371_),
    .Z(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2202_ (.I(_1303_),
    .Z(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _2203_ (.A1(_1301_),
    .A2(_1302_),
    .B1(_1211_),
    .B2(_1304_),
    .C(_1069_),
    .ZN(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2204_ (.A1(_1221_),
    .A2(_0701_),
    .A3(_1200_),
    .ZN(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2205_ (.A1(_1304_),
    .A2(_1201_),
    .B(_1306_),
    .C(_1178_),
    .ZN(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2206_ (.A1(_1218_),
    .A2(_1305_),
    .B1(_1307_),
    .B2(_1161_),
    .ZN(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2207_ (.A1(_1291_),
    .A2(_1300_),
    .B(_1308_),
    .ZN(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2208_ (.A1(_1020_),
    .A2(_1309_),
    .Z(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2209_ (.I(_1310_),
    .Z(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2210_ (.I(_1311_),
    .Z(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2211_ (.I(\dsynth.freeRunCntr[8] ),
    .Z(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2212_ (.I(_1313_),
    .Z(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2213_ (.A1(_1195_),
    .A2(_1201_),
    .ZN(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2214_ (.A1(_0624_),
    .A2(_0657_),
    .A3(_1297_),
    .ZN(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2215_ (.I(_1040_),
    .Z(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2216_ (.I(_1317_),
    .Z(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2217_ (.I(_1318_),
    .Z(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2218_ (.A1(_0393_),
    .A2(_1316_),
    .B(_1319_),
    .ZN(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2219_ (.I(_0448_),
    .Z(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2220_ (.A1(_1237_),
    .A2(_1321_),
    .A3(_1177_),
    .B(_0195_),
    .ZN(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2221_ (.I(_1175_),
    .Z(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2222_ (.A1(_0481_),
    .A2(_0855_),
    .A3(_1196_),
    .B(_0866_),
    .ZN(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2223_ (.A1(_1323_),
    .A2(_1201_),
    .B(_1324_),
    .ZN(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2224_ (.A1(_1315_),
    .A2(_1320_),
    .B1(_1322_),
    .B2(_1325_),
    .ZN(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2225_ (.A1(_0492_),
    .A2(_0283_),
    .B(_1239_),
    .ZN(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2226_ (.I(_1297_),
    .Z(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2227_ (.A1(_1238_),
    .A2(_1304_),
    .A3(_1328_),
    .B(_1180_),
    .ZN(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2228_ (.A1(_0833_),
    .A2(_1327_),
    .B(_1329_),
    .C(_0963_),
    .ZN(_1330_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2229_ (.A1(_1141_),
    .A2(_1297_),
    .ZN(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2230_ (.A1(_1214_),
    .A2(_1331_),
    .ZN(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _2231_ (.A1(_1245_),
    .A2(_1237_),
    .A3(_0459_),
    .A4(_1177_),
    .ZN(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2232_ (.A1(_1189_),
    .A2(_1049_),
    .ZN(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2233_ (.A1(_1332_),
    .A2(_1295_),
    .B(_1333_),
    .C(_1334_),
    .ZN(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2234_ (.A1(_1125_),
    .A2(_1326_),
    .B(_1330_),
    .C(_1335_),
    .ZN(_1336_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2235_ (.A1(_1188_),
    .A2(_1336_),
    .Z(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2236_ (.I(_1337_),
    .Z(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2237_ (.I(_1338_),
    .Z(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2238_ (.I(\dsynth.freeRunCntr[7] ),
    .Z(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2239_ (.A1(_1313_),
    .A2(_1312_),
    .B1(_1339_),
    .B2(_1340_),
    .ZN(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2240_ (.A1(_1271_),
    .A2(_1294_),
    .ZN(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2241_ (.A1(_1328_),
    .A2(_1222_),
    .ZN(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2242_ (.I(_0811_),
    .Z(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2243_ (.A1(_1275_),
    .A2(_1344_),
    .ZN(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2244_ (.A1(_1141_),
    .A2(_1155_),
    .ZN(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2245_ (.A1(_0327_),
    .A2(_0228_),
    .ZN(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2246_ (.A1(_1345_),
    .A2(_1346_),
    .B1(_1252_),
    .B2(_1347_),
    .ZN(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2247_ (.I(_0206_),
    .Z(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2248_ (.A1(_1342_),
    .A2(_1343_),
    .B1(_1348_),
    .B2(_1349_),
    .ZN(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2249_ (.I(_1146_),
    .Z(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2250_ (.A1(_1221_),
    .A2(_1351_),
    .ZN(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2251_ (.A1(_1352_),
    .A2(_1298_),
    .B(_1195_),
    .ZN(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2252_ (.I(_1321_),
    .Z(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2253_ (.I(_0789_),
    .Z(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2254_ (.A1(_1354_),
    .A2(_0767_),
    .A3(_1247_),
    .B(_1355_),
    .ZN(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2255_ (.A1(_1175_),
    .A2(_1246_),
    .ZN(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2256_ (.A1(_1220_),
    .A2(_1246_),
    .B(_1167_),
    .ZN(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2257_ (.A1(_1357_),
    .A2(_1358_),
    .ZN(_1359_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2258_ (.I(_0958_),
    .Z(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _2259_ (.A1(_1353_),
    .A2(_1356_),
    .B1(_1359_),
    .B2(_1320_),
    .C(_1360_),
    .ZN(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2260_ (.A1(_1125_),
    .A2(_1350_),
    .B(_1361_),
    .ZN(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2261_ (.A1(_1188_),
    .A2(_1362_),
    .Z(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2262_ (.I(_1363_),
    .Z(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2263_ (.I(_1364_),
    .Z(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2264_ (.A1(_1357_),
    .A2(_1358_),
    .Z(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2265_ (.A1(_1245_),
    .A2(_1221_),
    .ZN(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2266_ (.A1(_1275_),
    .A2(_1276_),
    .B(_1166_),
    .ZN(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2267_ (.A1(_1367_),
    .A2(_1368_),
    .ZN(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2268_ (.I(_1212_),
    .Z(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2269_ (.A1(_1366_),
    .A2(_1369_),
    .B(_1370_),
    .ZN(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2270_ (.A1(_1301_),
    .A2(_1258_),
    .B(_1272_),
    .C(_1202_),
    .ZN(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2271_ (.A1(_1125_),
    .A2(_1372_),
    .ZN(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2272_ (.I(_0888_),
    .Z(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2273_ (.A1(_1374_),
    .A2(_1237_),
    .B(_1344_),
    .C(_1223_),
    .ZN(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2274_ (.A1(_1207_),
    .A2(_1369_),
    .A3(_1375_),
    .Z(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2275_ (.A1(_1292_),
    .A2(_1329_),
    .B(_1291_),
    .ZN(_1377_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2276_ (.A1(_1371_),
    .A2(_1373_),
    .B1(_1376_),
    .B2(_1377_),
    .ZN(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2277_ (.A1(_0118_),
    .A2(_1378_),
    .Z(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2278_ (.I(_1379_),
    .Z(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2279_ (.I(_1380_),
    .ZN(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2280_ (.I(\dsynth.freeRunCntr[5] ),
    .Z(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2281_ (.A1(\dsynth.freeRunCntr[6] ),
    .A2(_1365_),
    .B1(_1381_),
    .B2(_1382_),
    .ZN(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2282_ (.I(_1383_),
    .ZN(_1384_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2283_ (.I(\dsynth.freeRunCntr[4] ),
    .Z(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2284_ (.A1(_0844_),
    .A2(_0228_),
    .B(_0272_),
    .ZN(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2285_ (.I(_0525_),
    .Z(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2286_ (.A1(_1218_),
    .A2(_1387_),
    .ZN(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2287_ (.I(_1304_),
    .Z(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2288_ (.A1(_1291_),
    .A2(_1386_),
    .B1(_1388_),
    .B2(_1152_),
    .C(_1389_),
    .ZN(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2289_ (.A1(_1331_),
    .A2(_1202_),
    .B(_1349_),
    .ZN(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2290_ (.A1(_1323_),
    .A2(_1243_),
    .B(_1354_),
    .ZN(_1392_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2291_ (.A1(_1374_),
    .A2(_1242_),
    .ZN(_1393_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2292_ (.I(_1393_),
    .Z(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2293_ (.A1(_1394_),
    .A2(_1277_),
    .B1(_1327_),
    .B2(_1367_),
    .C(_0206_),
    .ZN(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2294_ (.A1(_0558_),
    .A2(_0184_),
    .ZN(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2295_ (.A1(_1360_),
    .A2(_1392_),
    .A3(_1353_),
    .B1(_1395_),
    .B2(_1396_),
    .ZN(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2296_ (.A1(_1390_),
    .A2(_1391_),
    .B(_1397_),
    .ZN(_1398_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _2297_ (.A1(_0129_),
    .A2(_1398_),
    .Z(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _2298_ (.A1(_1344_),
    .A2(_1198_),
    .A3(_1386_),
    .B(_1059_),
    .ZN(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2299_ (.A1(_0712_),
    .A2(_0811_),
    .ZN(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2300_ (.I(_1401_),
    .Z(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2301_ (.I(_1351_),
    .Z(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2302_ (.I(_1360_),
    .Z(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2303_ (.A1(_1402_),
    .A2(_1403_),
    .B(_1404_),
    .ZN(_1405_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2304_ (.I(_0470_),
    .Z(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2305_ (.A1(_1406_),
    .A2(_1301_),
    .B(_1358_),
    .ZN(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2306_ (.A1(_1143_),
    .A2(_1194_),
    .A3(_1407_),
    .ZN(_1408_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2307_ (.A1(_1250_),
    .A2(_1252_),
    .B(_1370_),
    .C(_1179_),
    .ZN(_1409_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2308_ (.A1(_1253_),
    .A2(_1282_),
    .ZN(_1410_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2309_ (.I(_1218_),
    .Z(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2310_ (.A1(_1409_),
    .A2(_1410_),
    .B(_1411_),
    .ZN(_1412_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2311_ (.A1(_1400_),
    .A2(_1405_),
    .B(_1408_),
    .C(_1412_),
    .ZN(_1413_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2312_ (.A1(_1020_),
    .A2(_1413_),
    .Z(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2313_ (.I(_1414_),
    .Z(_1415_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2314_ (.I(_1415_),
    .Z(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2315_ (.I(\dsynth.freeRunCntr[3] ),
    .Z(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2316_ (.A1(_1385_),
    .A2(_1399_),
    .B1(_1416_),
    .B2(_1417_),
    .ZN(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2317_ (.I(\dsynth.freeRunCntr[2] ),
    .Z(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2318_ (.A1(_1347_),
    .A2(_1252_),
    .B(_1349_),
    .ZN(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _2319_ (.A1(_1319_),
    .A2(_1204_),
    .A3(_1323_),
    .A4(_1328_),
    .ZN(_1421_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2320_ (.A1(_1215_),
    .A2(_1421_),
    .Z(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2321_ (.A1(_1394_),
    .A2(_1420_),
    .B1(_1422_),
    .B2(_1366_),
    .ZN(_1423_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2322_ (.A1(_1345_),
    .A2(_1403_),
    .B(_1148_),
    .ZN(_1424_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2323_ (.A1(_1404_),
    .A2(_0767_),
    .A3(_1302_),
    .ZN(_1425_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2324_ (.A1(_1349_),
    .A2(_1199_),
    .A3(_1424_),
    .B1(_1425_),
    .B2(_1260_),
    .ZN(_1426_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2325_ (.A1(_1411_),
    .A2(_1423_),
    .B(_1426_),
    .ZN(_1427_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2326_ (.A1(_1030_),
    .A2(_1427_),
    .Z(_1428_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2327_ (.I(_1428_),
    .Z(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2328_ (.I(_1429_),
    .Z(_1430_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2329_ (.A1(_1419_),
    .A2(_1430_),
    .ZN(_1431_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2330_ (.A1(_0261_),
    .A2(_1197_),
    .Z(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2331_ (.A1(_1239_),
    .A2(_1432_),
    .ZN(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2332_ (.I(_1370_),
    .Z(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _2333_ (.A1(_1359_),
    .A2(_1432_),
    .B1(_1433_),
    .B2(_1247_),
    .C(_1434_),
    .ZN(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2334_ (.A1(_1434_),
    .A2(_1199_),
    .A3(_1368_),
    .ZN(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2335_ (.A1(_1404_),
    .A2(_1436_),
    .ZN(_1437_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2336_ (.A1(_1142_),
    .A2(_1155_),
    .B(_1239_),
    .C(_1141_),
    .ZN(_1438_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2337_ (.A1(_1434_),
    .A2(_1438_),
    .Z(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _2338_ (.A1(_1224_),
    .A2(_1205_),
    .B1(_1258_),
    .B2(_1387_),
    .C(_1434_),
    .ZN(_1440_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2339_ (.A1(_1387_),
    .A2(_1357_),
    .A3(_1439_),
    .B(_1440_),
    .ZN(_1441_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2340_ (.A1(_1435_),
    .A2(_1437_),
    .B1(_1441_),
    .B2(_1404_),
    .ZN(_1442_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2341_ (.A1(_1030_),
    .A2(_1442_),
    .Z(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2342_ (.I(_1443_),
    .Z(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2343_ (.I(\dsynth.freeRunCntr[1] ),
    .Z(_1445_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2344_ (.A1(_1419_),
    .A2(_1430_),
    .B1(_1444_),
    .B2(_1445_),
    .ZN(_1446_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2345_ (.A1(_1431_),
    .A2(_1446_),
    .ZN(_1447_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2346_ (.A1(_1417_),
    .A2(_1416_),
    .B(_1447_),
    .ZN(_1448_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2347_ (.A1(\dsynth.freeRunCntr[4] ),
    .A2(_1399_),
    .B1(_1381_),
    .B2(_1382_),
    .ZN(_1449_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2348_ (.A1(_1418_),
    .A2(_1448_),
    .B(_1449_),
    .ZN(_1450_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2349_ (.I(\dsynth.freeRunCntr[6] ),
    .Z(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _2350_ (.A1(_1340_),
    .A2(_1339_),
    .B1(_1384_),
    .B2(_1450_),
    .C1(_1365_),
    .C2(_1451_),
    .ZN(_1452_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2351_ (.A1(_1341_),
    .A2(_1452_),
    .ZN(_1453_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2352_ (.A1(_1290_),
    .A2(_1287_),
    .B1(_1312_),
    .B2(_1314_),
    .C(_1453_),
    .ZN(_1454_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2353_ (.A1(_1289_),
    .A2(_1454_),
    .Z(_1455_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2354_ (.A1(_1187_),
    .A2(_1231_),
    .B1(_1269_),
    .B2(_1455_),
    .ZN(_1456_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2355_ (.A1(_0140_),
    .A2(_1134_),
    .B1(_1139_),
    .B2(_1456_),
    .ZN(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2356_ (.A1(_1290_),
    .A2(_1287_),
    .B(_1289_),
    .C(_1139_),
    .ZN(_1458_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2357_ (.I(_1314_),
    .Z(_1459_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2358_ (.A1(_1459_),
    .A2(_1312_),
    .B(_1431_),
    .C(_1383_),
    .ZN(_1460_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2359_ (.I(_1340_),
    .Z(_1461_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2360_ (.A1(_1461_),
    .A2(_1339_),
    .B1(_1365_),
    .B2(_1451_),
    .C(_1418_),
    .ZN(_1462_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2361_ (.I(_1417_),
    .Z(_1463_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2362_ (.I(_1463_),
    .Z(_1464_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2363_ (.I(_1445_),
    .Z(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2364_ (.A1(_1465_),
    .A2(_1444_),
    .B(_1449_),
    .ZN(_1466_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2365_ (.A1(_1464_),
    .A2(_1416_),
    .B(_1466_),
    .C(_1341_),
    .ZN(_1467_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2366_ (.A1(_1446_),
    .A2(_1460_),
    .A3(_1462_),
    .A4(_1467_),
    .Z(_1468_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2367_ (.A1(_1269_),
    .A2(_1458_),
    .A3(_1468_),
    .ZN(_1469_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2368_ (.A1(_1457_),
    .A2(_1469_),
    .Z(_1470_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2369_ (.I(_1470_),
    .Z(net27));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2370_ (.I(\dsynth.freeRunCntr[32] ),
    .ZN(_1471_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2371_ (.I(_1471_),
    .Z(_1472_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2372_ (.I(_1472_),
    .Z(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2373_ (.I(\dsynth.freeRunCntr[31] ),
    .Z(_1474_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2374_ (.I(_1474_),
    .Z(_1475_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2375_ (.I(_1475_),
    .Z(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2376_ (.I(\dsynth.freeRunCntr[29] ),
    .Z(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2377_ (.A1(_1476_),
    .A2(_1477_),
    .ZN(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2378_ (.A1(_1473_),
    .A2(_1478_),
    .Z(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2379_ (.A1(_1286_),
    .A2(_1479_),
    .ZN(_1480_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2380_ (.I(\dsynth.freeRunCntr[32] ),
    .Z(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2381_ (.I(\dsynth.freeRunCntr[29] ),
    .ZN(_1482_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2382_ (.A1(_1481_),
    .A2(_1482_),
    .ZN(_1483_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2383_ (.I(_1483_),
    .Z(_1484_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2384_ (.A1(\dsynth.freeRunCntr[30] ),
    .A2(_1474_),
    .Z(_1485_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2385_ (.I(\dsynth.freeRunCntr[30] ),
    .Z(_1486_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2386_ (.A1(_1486_),
    .A2(_1474_),
    .A3(\dsynth.freeRunCntr[29] ),
    .B(_1481_),
    .ZN(_1487_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2387_ (.A1(_1481_),
    .A2(_1485_),
    .B(_1487_),
    .ZN(_1488_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2388_ (.A1(_1484_),
    .A2(_1488_),
    .Z(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2389_ (.I(_1489_),
    .Z(_1490_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2390_ (.A1(_1475_),
    .A2(_1472_),
    .A3(_1482_),
    .ZN(_1491_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2391_ (.I(_1491_),
    .Z(_1492_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2392_ (.I(_1492_),
    .Z(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2393_ (.A1(_0118_),
    .A2(_1493_),
    .ZN(_1494_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2394_ (.A1(_1228_),
    .A2(_1490_),
    .B(_1494_),
    .ZN(_1495_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2395_ (.A1(_1480_),
    .A2(_1495_),
    .ZN(_1496_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2396_ (.I(_1496_),
    .ZN(_1497_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2397_ (.I(_1494_),
    .Z(_1498_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2398_ (.A1(\dsynth.freeRunCntr[31] ),
    .A2(_1471_),
    .ZN(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2399_ (.A1(_1477_),
    .A2(_1499_),
    .ZN(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2400_ (.I(_1500_),
    .Z(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2401_ (.A1(_1127_),
    .A2(_1501_),
    .ZN(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2402_ (.I(_1502_),
    .Z(_1503_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2403_ (.I(_1500_),
    .Z(_1504_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2404_ (.A1(_1227_),
    .A2(_1504_),
    .ZN(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2405_ (.I(_1505_),
    .Z(_1506_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2406_ (.A1(_1228_),
    .A2(_1504_),
    .Z(_1507_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2407_ (.A1(_1128_),
    .A2(_1507_),
    .Z(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2408_ (.A1(_1503_),
    .A2(_1506_),
    .B(_1508_),
    .ZN(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2409_ (.A1(_1498_),
    .A2(_1509_),
    .B(_1508_),
    .ZN(_1510_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2410_ (.A1(_1497_),
    .A2(_1510_),
    .ZN(_1511_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2411_ (.A1(_1496_),
    .A2(_1510_),
    .Z(_1512_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2412_ (.I(\dsynth.freeRunCntr[30] ),
    .ZN(_1513_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _2413_ (.A1(_1513_),
    .A2(_1476_),
    .A3(_1473_),
    .ZN(_1514_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2414_ (.I(_1514_),
    .Z(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2415_ (.I(_0096_),
    .Z(_1516_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2416_ (.A1(_1171_),
    .A2(_1172_),
    .ZN(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2417_ (.A1(_0756_),
    .A2(_1517_),
    .B1(_1211_),
    .B2(_1281_),
    .ZN(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2418_ (.A1(_1374_),
    .A2(_0459_),
    .B1(_1159_),
    .B2(_1327_),
    .C(_0778_),
    .ZN(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2419_ (.A1(_0789_),
    .A2(_1518_),
    .B(_1519_),
    .ZN(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2420_ (.A1(_1351_),
    .A2(_1210_),
    .B(_1213_),
    .ZN(_1521_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2421_ (.A1(_1303_),
    .A2(_1295_),
    .Z(_1522_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2422_ (.A1(_0492_),
    .A2(_0239_),
    .B(_0448_),
    .ZN(_1523_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _2423_ (.A1(_0382_),
    .A2(_1316_),
    .B1(_1523_),
    .B2(_1163_),
    .C(_1272_),
    .ZN(_1524_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2424_ (.A1(_1318_),
    .A2(_1521_),
    .A3(_1522_),
    .B(_1524_),
    .ZN(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2425_ (.I0(_1520_),
    .I1(_1525_),
    .S(_0958_),
    .Z(_1526_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2426_ (.A1(_1516_),
    .A2(_1526_),
    .Z(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2427_ (.I(_1527_),
    .Z(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2428_ (.A1(_1513_),
    .A2(_1483_),
    .Z(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2429_ (.A1(_1475_),
    .A2(_1529_),
    .ZN(_1530_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2430_ (.I(_1530_),
    .Z(_1531_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2431_ (.I(_1531_),
    .ZN(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2432_ (.I(_1001_),
    .Z(_1533_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _2433_ (.A1(_1198_),
    .A2(_1205_),
    .B1(_1324_),
    .B2(_1386_),
    .C(_1317_),
    .ZN(_1534_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2434_ (.A1(_0184_),
    .A2(_1271_),
    .A3(_1274_),
    .ZN(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2435_ (.A1(_1191_),
    .A2(_1534_),
    .A3(_1535_),
    .Z(_1536_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2436_ (.A1(_0690_),
    .A2(_1295_),
    .B(_1317_),
    .ZN(_1537_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2437_ (.A1(_1140_),
    .A2(_0855_),
    .B(_0679_),
    .ZN(_1538_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2438_ (.A1(_1274_),
    .A2(_1150_),
    .B1(_1209_),
    .B2(_1538_),
    .ZN(_1539_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _2439_ (.A1(_1433_),
    .A2(_1537_),
    .B1(_1539_),
    .B2(_1192_),
    .C(_1191_),
    .ZN(_1540_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _2440_ (.A1(_1533_),
    .A2(_1536_),
    .A3(_1540_),
    .Z(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2441_ (.A1(_1536_),
    .A2(_1540_),
    .B(_1533_),
    .ZN(_1542_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2442_ (.A1(_1541_),
    .A2(_1542_),
    .Z(_1543_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2443_ (.I(_1543_),
    .Z(_1544_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2444_ (.A1(\dsynth.freeRunCntr[29] ),
    .A2(_1485_),
    .ZN(_1545_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2445_ (.A1(_1472_),
    .A2(_1545_),
    .ZN(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2446_ (.A1(_1487_),
    .A2(_1546_),
    .ZN(_1547_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2447_ (.I(_1547_),
    .Z(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2448_ (.I(_1548_),
    .Z(_1549_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2449_ (.A1(_1176_),
    .A2(_1294_),
    .Z(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2450_ (.A1(_0701_),
    .A2(_1550_),
    .ZN(_1551_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2451_ (.A1(_1140_),
    .A2(_0646_),
    .A3(_0437_),
    .ZN(_1552_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2452_ (.A1(_1240_),
    .A2(_1552_),
    .Z(_1553_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2453_ (.A1(_1551_),
    .A2(_1553_),
    .B(_1396_),
    .ZN(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2454_ (.I(_0745_),
    .Z(_1555_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2455_ (.A1(_1172_),
    .A2(_1555_),
    .ZN(_1556_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2456_ (.A1(_1555_),
    .A2(_1294_),
    .ZN(_1557_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2457_ (.A1(_1402_),
    .A2(_1393_),
    .B(_1556_),
    .C(_1557_),
    .ZN(_1558_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2458_ (.A1(_1156_),
    .A2(_1173_),
    .A3(_1253_),
    .B(_0569_),
    .ZN(_1559_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2459_ (.A1(_1303_),
    .A2(_1555_),
    .B(_1171_),
    .ZN(_1560_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2460_ (.A1(_1318_),
    .A2(_1438_),
    .A3(_1560_),
    .B(_1217_),
    .ZN(_1561_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2461_ (.A1(_1194_),
    .A2(_1558_),
    .B1(_1559_),
    .B2(_1561_),
    .ZN(_1562_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2462_ (.A1(_1554_),
    .A2(_1562_),
    .B(_1516_),
    .ZN(_1563_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2463_ (.I(_0096_),
    .Z(_1564_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2464_ (.A1(_1564_),
    .A2(_1554_),
    .A3(_1562_),
    .Z(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2465_ (.A1(_1563_),
    .A2(_1565_),
    .ZN(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _2466_ (.A1(_1515_),
    .A2(_1528_),
    .B1(_1532_),
    .B2(_1544_),
    .C1(_1549_),
    .C2(_1566_),
    .ZN(_1567_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2467_ (.I(_1567_),
    .ZN(_1568_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2468_ (.I(_1533_),
    .Z(_1569_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2469_ (.A1(_1354_),
    .A2(_0833_),
    .A3(_1161_),
    .ZN(_1570_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _2470_ (.A1(_0800_),
    .A2(_1078_),
    .B(_1333_),
    .C(_0580_),
    .ZN(_1571_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _2471_ (.A1(_1569_),
    .A2(_1570_),
    .A3(_1571_),
    .Z(_1572_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2472_ (.I(_1001_),
    .Z(_1573_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2473_ (.I(_1573_),
    .Z(_1574_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2474_ (.A1(_1570_),
    .A2(_1571_),
    .B(_1574_),
    .ZN(_1575_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2475_ (.A1(_1572_),
    .A2(_1575_),
    .ZN(_1576_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2476_ (.A1(\dsynth.freeRunCntr[30] ),
    .A2(_1499_),
    .ZN(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2477_ (.I(_1577_),
    .Z(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2478_ (.I(_1578_),
    .Z(_1579_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2479_ (.I(_1579_),
    .Z(_1580_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2480_ (.A1(_1566_),
    .A2(_1580_),
    .ZN(_1581_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2481_ (.A1(_1180_),
    .A2(_1333_),
    .ZN(_1582_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2482_ (.A1(_1235_),
    .A2(_1078_),
    .A3(_1582_),
    .ZN(_1583_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2483_ (.A1(_1516_),
    .A2(_1583_),
    .Z(_1584_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2484_ (.A1(_1579_),
    .A2(_1584_),
    .ZN(_1585_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2485_ (.A1(_1572_),
    .A2(_1575_),
    .Z(_1586_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2486_ (.I(_1578_),
    .Z(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2487_ (.A1(_1572_),
    .A2(_1575_),
    .B(_1587_),
    .ZN(_1588_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2488_ (.A1(_1513_),
    .A2(_1474_),
    .A3(_1471_),
    .ZN(_1589_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2489_ (.I(_1589_),
    .Z(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2490_ (.A1(_1563_),
    .A2(_1565_),
    .B(_1590_),
    .ZN(_1591_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2491_ (.I0(_1586_),
    .I1(_1588_),
    .S(_1591_),
    .Z(_1592_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2492_ (.A1(_1576_),
    .A2(_1581_),
    .B1(_1585_),
    .B2(_1592_),
    .ZN(_1593_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2493_ (.I(_1590_),
    .Z(_1594_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2494_ (.A1(_1236_),
    .A2(_1355_),
    .A3(_1333_),
    .ZN(_1595_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _2495_ (.A1(_1569_),
    .A2(_1595_),
    .Z(_1596_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2496_ (.A1(_1594_),
    .A2(_1596_),
    .ZN(_1597_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2497_ (.A1(_1374_),
    .A2(_1555_),
    .ZN(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2498_ (.A1(_1298_),
    .A2(_1598_),
    .B(_1281_),
    .ZN(_1599_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2499_ (.A1(_1281_),
    .A2(_1432_),
    .ZN(_1600_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2500_ (.A1(_0459_),
    .A2(_1331_),
    .A3(_1270_),
    .B(_0931_),
    .ZN(_1601_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _2501_ (.A1(_1400_),
    .A2(_1599_),
    .B1(_1600_),
    .B2(_1601_),
    .C(_1217_),
    .ZN(_1602_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2502_ (.A1(_1234_),
    .A2(_0195_),
    .A3(_1321_),
    .ZN(_1603_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2503_ (.A1(_1303_),
    .A2(_1200_),
    .ZN(_1604_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2504_ (.A1(_1165_),
    .A2(_1257_),
    .B(_1604_),
    .ZN(_1605_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2505_ (.A1(_1159_),
    .A2(_1603_),
    .B1(_1605_),
    .B2(_1193_),
    .ZN(_1606_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2506_ (.A1(_1573_),
    .A2(_1602_),
    .A3(_1606_),
    .Z(_1607_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2507_ (.A1(_1602_),
    .A2(_1606_),
    .B(_1573_),
    .ZN(_1608_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2508_ (.A1(_1578_),
    .A2(_1607_),
    .A3(_1608_),
    .ZN(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2509_ (.I0(_1585_),
    .I1(_1584_),
    .S(_1609_),
    .Z(_1610_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2510_ (.A1(_1597_),
    .A2(_1610_),
    .Z(_1611_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2511_ (.A1(_1593_),
    .A2(_1611_),
    .ZN(_1612_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2512_ (.A1(_1593_),
    .A2(_1611_),
    .Z(_1613_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2513_ (.A1(_1568_),
    .A2(_1612_),
    .B(_1613_),
    .ZN(_1614_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2514_ (.A1(_1184_),
    .A2(_1500_),
    .Z(_1615_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2515_ (.A1(_1513_),
    .A2(_1475_),
    .A3(_1472_),
    .Z(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2516_ (.I(_1616_),
    .Z(_1617_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2517_ (.A1(_1541_),
    .A2(_1542_),
    .ZN(_1618_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2518_ (.A1(_1142_),
    .A2(_1200_),
    .B(_1166_),
    .ZN(_1619_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2519_ (.A1(_1256_),
    .A2(_1342_),
    .B(_1163_),
    .ZN(_1620_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _2520_ (.A1(_1619_),
    .A2(_1272_),
    .B1(_1620_),
    .B2(_0195_),
    .C(_1234_),
    .ZN(_1621_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2521_ (.A1(_1517_),
    .A2(_1270_),
    .ZN(_1622_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2522_ (.A1(_1143_),
    .A2(_1346_),
    .A3(_1396_),
    .ZN(_1623_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2523_ (.A1(_0668_),
    .A2(_1344_),
    .A3(_1276_),
    .B(_0778_),
    .ZN(_1624_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2524_ (.A1(_1213_),
    .A2(_1242_),
    .B(_1234_),
    .ZN(_1625_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2525_ (.A1(_1622_),
    .A2(_1623_),
    .B1(_1624_),
    .B2(_1625_),
    .ZN(_1626_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _2526_ (.A1(_1564_),
    .A2(_1621_),
    .A3(_1626_),
    .Z(_1627_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2527_ (.A1(_1621_),
    .A2(_1626_),
    .B(_1564_),
    .ZN(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2528_ (.A1(_1627_),
    .A2(_1628_),
    .ZN(_1629_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2529_ (.I(_1530_),
    .Z(_1630_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2530_ (.A1(_1617_),
    .A2(_1618_),
    .B1(_1629_),
    .B2(_1630_),
    .ZN(_1631_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2531_ (.A1(_1615_),
    .A2(_1631_),
    .Z(_1632_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2532_ (.I(_1533_),
    .Z(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2533_ (.A1(_1633_),
    .A2(_1583_),
    .Z(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2534_ (.I(_1609_),
    .Z(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2535_ (.I(_1564_),
    .Z(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2536_ (.A1(_1636_),
    .A2(_1595_),
    .Z(_1637_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2537_ (.A1(_1580_),
    .A2(_1637_),
    .ZN(_1638_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2538_ (.A1(_1634_),
    .A2(_1635_),
    .B1(_1610_),
    .B2(_1638_),
    .ZN(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2539_ (.A1(_1607_),
    .A2(_1608_),
    .ZN(_1640_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2540_ (.I(_1487_),
    .ZN(_1641_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2541_ (.A1(_1473_),
    .A2(_1545_),
    .B(_1641_),
    .ZN(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2542_ (.A1(_1347_),
    .A2(_1538_),
    .A3(_1209_),
    .ZN(_1643_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2543_ (.A1(_1190_),
    .A2(_0173_),
    .ZN(_1644_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2544_ (.A1(_1149_),
    .A2(_1152_),
    .B(_1644_),
    .ZN(_1645_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _2545_ (.A1(_0822_),
    .A2(_0360_),
    .B(_0547_),
    .C(_0162_),
    .ZN(_1646_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2546_ (.A1(_1162_),
    .A2(_1292_),
    .A3(_1646_),
    .B1(_1552_),
    .B2(_1153_),
    .ZN(_1647_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2547_ (.A1(_1140_),
    .A2(_0228_),
    .A3(_1196_),
    .ZN(_1648_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2548_ (.A1(_1149_),
    .A2(_1648_),
    .B1(_1251_),
    .B2(_1274_),
    .C(_1334_),
    .ZN(_1649_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2549_ (.A1(_1643_),
    .A2(_1645_),
    .B(_1647_),
    .C(_1649_),
    .ZN(_1650_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2550_ (.A1(_0096_),
    .A2(_1650_),
    .Z(_1651_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2551_ (.A1(_1589_),
    .A2(_1651_),
    .ZN(_1652_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2552_ (.I(_1652_),
    .Z(_1653_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2553_ (.A1(_1597_),
    .A2(_1653_),
    .ZN(_1654_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2554_ (.I(_1651_),
    .Z(_1655_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2555_ (.A1(_1638_),
    .A2(_1655_),
    .ZN(_1656_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2556_ (.A1(_1640_),
    .A2(_1642_),
    .B1(_1654_),
    .B2(_1656_),
    .ZN(_1657_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2557_ (.A1(_1639_),
    .A2(_1657_),
    .Z(_1658_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2558_ (.A1(_1632_),
    .A2(_1658_),
    .Z(_1659_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2559_ (.A1(_1614_),
    .A2(_1659_),
    .ZN(_1660_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2560_ (.A1(_1614_),
    .A2(_1659_),
    .ZN(_1661_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2561_ (.A1(_1512_),
    .A2(_1660_),
    .B(_1661_),
    .ZN(_1662_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2562_ (.A1(_1480_),
    .A2(_1495_),
    .ZN(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2563_ (.I(_1615_),
    .Z(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2564_ (.A1(_1664_),
    .A2(_1631_),
    .ZN(_1665_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2565_ (.I(_1479_),
    .Z(_1666_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2566_ (.I(_1666_),
    .Z(_1667_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2567_ (.I(_1667_),
    .Z(_1668_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2568_ (.A1(_1486_),
    .A2(_1476_),
    .Z(_1669_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _2569_ (.A1(_1484_),
    .A2(_1669_),
    .ZN(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _2570_ (.A1(_1266_),
    .A2(_1668_),
    .B1(_1670_),
    .B2(_1287_),
    .ZN(_1671_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2571_ (.A1(_1663_),
    .A2(_1665_),
    .A3(_1671_),
    .Z(_1672_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2572_ (.A1(_1639_),
    .A2(_1657_),
    .ZN(_1673_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2573_ (.A1(_1632_),
    .A2(_1658_),
    .B(_1673_),
    .ZN(_1674_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2574_ (.I(_1490_),
    .Z(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2575_ (.I(_1675_),
    .Z(_1676_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2576_ (.I(_1629_),
    .ZN(_1677_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2577_ (.I(_1677_),
    .Z(_1678_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2578_ (.A1(_1137_),
    .A2(_1491_),
    .ZN(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _2579_ (.A1(_1185_),
    .A2(_1676_),
    .B1(_1515_),
    .B2(_1678_),
    .C(_1679_),
    .ZN(_1680_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2580_ (.I(_1637_),
    .Z(_1681_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2581_ (.A1(_1681_),
    .A2(_1653_),
    .ZN(_1682_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2582_ (.I(_1566_),
    .Z(_1683_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2583_ (.A1(_1683_),
    .A2(_1532_),
    .ZN(_1684_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2584_ (.I(_1642_),
    .Z(_1685_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2585_ (.A1(_1685_),
    .A2(_1655_),
    .ZN(_1686_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2586_ (.I(_1594_),
    .Z(_1687_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2587_ (.A1(_0448_),
    .A2(_0833_),
    .ZN(_1688_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2588_ (.A1(_1190_),
    .A2(_1317_),
    .A3(_1401_),
    .A4(_0382_),
    .ZN(_1689_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _2589_ (.A1(_0920_),
    .A2(_1644_),
    .B1(_1646_),
    .B2(_1688_),
    .C(_1689_),
    .ZN(_1690_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2590_ (.A1(_1636_),
    .A2(_1690_),
    .Z(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2591_ (.A1(_1687_),
    .A2(_1691_),
    .ZN(_1692_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2592_ (.A1(_1686_),
    .A2(_1692_),
    .ZN(_1693_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2593_ (.A1(_1684_),
    .A2(_1693_),
    .Z(_1694_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2594_ (.A1(_1682_),
    .A2(_1694_),
    .Z(_1695_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2595_ (.A1(_1680_),
    .A2(_1695_),
    .ZN(_1696_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2596_ (.A1(_1674_),
    .A2(_1696_),
    .ZN(_1697_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2597_ (.A1(_1672_),
    .A2(_1697_),
    .Z(_1698_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _2598_ (.A1(_1511_),
    .A2(_1662_),
    .A3(_1698_),
    .ZN(_1699_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2599_ (.I(_1670_),
    .Z(_1700_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2600_ (.A1(_1124_),
    .A2(_1087_),
    .Z(_1701_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2601_ (.I(_1701_),
    .Z(_1702_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2602_ (.A1(_1264_),
    .A2(_1501_),
    .ZN(_1703_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2603_ (.I(_1703_),
    .Z(_1704_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2604_ (.A1(_1701_),
    .A2(_1491_),
    .ZN(_1705_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2605_ (.I(_1705_),
    .Z(_1706_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2606_ (.I(_1703_),
    .ZN(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2607_ (.A1(_1706_),
    .A2(_1707_),
    .ZN(_1708_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2608_ (.A1(_1702_),
    .A2(_1704_),
    .B1(_1708_),
    .B2(_1503_),
    .ZN(_1709_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2609_ (.A1(_1498_),
    .A2(_1509_),
    .ZN(_1710_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2610_ (.A1(_1312_),
    .A2(_1700_),
    .B1(_1709_),
    .B2(_1710_),
    .ZN(_1711_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2611_ (.A1(_1709_),
    .A2(_1710_),
    .ZN(_1712_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2612_ (.A1(_1633_),
    .A2(_1526_),
    .Z(_1713_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2613_ (.I(_1713_),
    .Z(_1714_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2614_ (.I(_1531_),
    .Z(_1715_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2615_ (.A1(_1321_),
    .A2(_1177_),
    .ZN(_1716_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2616_ (.A1(_1347_),
    .A2(_1716_),
    .B(_1206_),
    .ZN(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2617_ (.A1(_1219_),
    .A2(_1275_),
    .A3(_1276_),
    .ZN(_1718_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2618_ (.A1(_1148_),
    .A2(_1718_),
    .ZN(_1719_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2619_ (.I0(_1150_),
    .I1(_1251_),
    .S(_1210_),
    .Z(_1720_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _2620_ (.A1(_1717_),
    .A2(_1719_),
    .B1(_1720_),
    .B2(_1319_),
    .C(_1259_),
    .ZN(_1721_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2621_ (.A1(_1243_),
    .A2(_1150_),
    .B1(_1282_),
    .B2(_1538_),
    .ZN(_1722_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2622_ (.A1(_0958_),
    .A2(_1206_),
    .A3(_1402_),
    .A4(_1257_),
    .ZN(_1723_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2623_ (.A1(_1161_),
    .A2(_1722_),
    .B1(_1723_),
    .B2(_0404_),
    .ZN(_1724_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2624_ (.A1(_1721_),
    .A2(_1724_),
    .B(_1569_),
    .ZN(_1725_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _2625_ (.A1(_1633_),
    .A2(_1721_),
    .A3(_1724_),
    .Z(_1726_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2626_ (.A1(_1725_),
    .A2(_1726_),
    .ZN(_1727_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2627_ (.I(_1727_),
    .Z(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _2628_ (.A1(_1714_),
    .A2(_1715_),
    .B1(_1629_),
    .B2(_1685_),
    .C1(_1728_),
    .C2(_1617_),
    .ZN(_1729_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2629_ (.A1(_1001_),
    .A2(_1690_),
    .Z(_1730_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2630_ (.A1(_1577_),
    .A2(_1730_),
    .ZN(_1731_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2631_ (.I(_1731_),
    .Z(_1732_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2632_ (.A1(_1627_),
    .A2(_1628_),
    .B(_1578_),
    .ZN(_1733_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2633_ (.I(_1733_),
    .Z(_1734_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2634_ (.A1(_1732_),
    .A2(_1734_),
    .ZN(_1735_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2635_ (.I(_1594_),
    .Z(_1736_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2636_ (.A1(_1576_),
    .A2(_1736_),
    .ZN(_1737_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2637_ (.A1(_1677_),
    .A2(_1692_),
    .B1(_1735_),
    .B2(_1737_),
    .ZN(_1738_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2638_ (.A1(_1585_),
    .A2(_1592_),
    .Z(_1739_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2639_ (.A1(_1738_),
    .A2(_1739_),
    .ZN(_1740_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2640_ (.A1(_1738_),
    .A2(_1739_),
    .ZN(_1741_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2641_ (.A1(_1729_),
    .A2(_1740_),
    .B(_1741_),
    .ZN(_1742_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2642_ (.A1(_1568_),
    .A2(_1612_),
    .Z(_1743_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2643_ (.A1(_1742_),
    .A2(_1743_),
    .ZN(_1744_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2644_ (.A1(_1742_),
    .A2(_1743_),
    .ZN(_1745_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2645_ (.A1(_1712_),
    .A2(_1744_),
    .B(_1745_),
    .ZN(_1746_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2646_ (.A1(_1512_),
    .A2(_1660_),
    .Z(_1747_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2647_ (.A1(_1746_),
    .A2(_1747_),
    .Z(_1748_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2648_ (.A1(_1746_),
    .A2(_1747_),
    .Z(_1749_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2649_ (.A1(_1711_),
    .A2(_1748_),
    .B(_1749_),
    .ZN(_1750_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2650_ (.A1(_1699_),
    .A2(_1750_),
    .Z(_1751_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2651_ (.A1(_1328_),
    .A2(_1302_),
    .ZN(_1752_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _2652_ (.A1(_1244_),
    .A2(_1153_),
    .A3(_1599_),
    .A4(_1752_),
    .ZN(_1753_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2653_ (.A1(_1345_),
    .A2(_1351_),
    .B1(_1718_),
    .B2(_1156_),
    .C(_1318_),
    .ZN(_1754_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2654_ (.A1(_1173_),
    .A2(_1279_),
    .B(_1368_),
    .C(_0789_),
    .ZN(_1755_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2655_ (.A1(_1245_),
    .A2(_0514_),
    .B(_1210_),
    .ZN(_1756_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2656_ (.A1(_1538_),
    .A2(_1756_),
    .B(_1375_),
    .C(_1193_),
    .ZN(_1757_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2657_ (.A1(_1259_),
    .A2(_1754_),
    .A3(_1755_),
    .B(_1757_),
    .ZN(_1758_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _2658_ (.A1(_1573_),
    .A2(_1753_),
    .A3(_1758_),
    .Z(_1759_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2659_ (.A1(_1753_),
    .A2(_1758_),
    .B(_1633_),
    .ZN(_1760_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2660_ (.A1(_1759_),
    .A2(_1760_),
    .ZN(_1761_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2661_ (.A1(_1286_),
    .A2(_1500_),
    .ZN(_1762_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2662_ (.A1(_1616_),
    .A2(_1761_),
    .B(_1762_),
    .ZN(_1763_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2663_ (.A1(_1679_),
    .A2(_1763_),
    .Z(_1764_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2664_ (.I(_1715_),
    .Z(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2665_ (.A1(_1547_),
    .A2(_1544_),
    .B(_1597_),
    .ZN(_1766_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2666_ (.A1(_1765_),
    .A2(_1728_),
    .A3(_1766_),
    .ZN(_1767_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2667_ (.I0(_1705_),
    .I1(_1702_),
    .S(_1703_),
    .Z(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2668_ (.A1(_1503_),
    .A2(_1768_),
    .Z(_1769_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2669_ (.A1(_1767_),
    .A2(_1769_),
    .ZN(_1770_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2670_ (.A1(_1767_),
    .A2(_1769_),
    .Z(_1771_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2671_ (.A1(_1764_),
    .A2(_1770_),
    .B(_1771_),
    .ZN(_1772_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_4 _2672_ (.A1(_1311_),
    .A2(_1667_),
    .B1(_1670_),
    .B2(_1339_),
    .C1(_1676_),
    .C2(_1265_),
    .ZN(_1773_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2673_ (.A1(_1772_),
    .A2(_1773_),
    .ZN(_1774_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_4 _2674_ (.A1(_1338_),
    .A2(_1666_),
    .B1(_1670_),
    .B2(_1364_),
    .C1(_1675_),
    .C2(_1286_),
    .ZN(_1775_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2675_ (.A1(_1087_),
    .A2(_1498_),
    .ZN(_1776_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2676_ (.A1(_1775_),
    .A2(_1776_),
    .ZN(_1777_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2677_ (.A1(_1772_),
    .A2(_1773_),
    .ZN(_1778_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2678_ (.A1(_1774_),
    .A2(_1777_),
    .B(_1778_),
    .ZN(_1779_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2679_ (.A1(_1774_),
    .A2(_1777_),
    .Z(_1780_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2680_ (.A1(_1764_),
    .A2(_1770_),
    .ZN(_1781_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2681_ (.I(_1588_),
    .Z(_1782_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2682_ (.I0(_1732_),
    .I1(_1730_),
    .S(_1733_),
    .Z(_1783_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2683_ (.A1(_1782_),
    .A2(_1783_),
    .Z(_1784_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2684_ (.A1(_1594_),
    .A2(_1651_),
    .Z(_1785_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2685_ (.A1(_1541_),
    .A2(_1542_),
    .B(_1577_),
    .ZN(_1786_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2686_ (.I0(_1543_),
    .I1(_1786_),
    .S(_1652_),
    .Z(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2687_ (.A1(_1618_),
    .A2(_1785_),
    .B1(_1732_),
    .B2(_1787_),
    .ZN(_1788_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2688_ (.A1(_1782_),
    .A2(_1783_),
    .ZN(_1789_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2689_ (.A1(_1531_),
    .A2(_1727_),
    .ZN(_1790_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2690_ (.A1(_1790_),
    .A2(_1766_),
    .Z(_1791_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2691_ (.A1(_1588_),
    .A2(_1783_),
    .Z(_1792_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2692_ (.A1(_1788_),
    .A2(_1792_),
    .Z(_1793_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2693_ (.A1(_1784_),
    .A2(_1788_),
    .A3(_1789_),
    .B1(_1791_),
    .B2(_1793_),
    .ZN(_1794_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2694_ (.A1(_1729_),
    .A2(_1740_),
    .Z(_1795_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2695_ (.A1(_1794_),
    .A2(_1795_),
    .ZN(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2696_ (.A1(_1794_),
    .A2(_1795_),
    .ZN(_1797_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2697_ (.A1(_1781_),
    .A2(_1796_),
    .B(_1797_),
    .ZN(_1798_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2698_ (.A1(_1712_),
    .A2(_1744_),
    .Z(_1799_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2699_ (.A1(_1798_),
    .A2(_1799_),
    .Z(_1800_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2700_ (.A1(_1798_),
    .A2(_1799_),
    .Z(_1801_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2701_ (.A1(_1780_),
    .A2(_1800_),
    .B(_1801_),
    .ZN(_1802_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2702_ (.A1(_1711_),
    .A2(_1748_),
    .ZN(_1803_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2703_ (.A1(_1802_),
    .A2(_1803_),
    .Z(_1804_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2704_ (.A1(_1802_),
    .A2(_1803_),
    .ZN(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2705_ (.A1(_1779_),
    .A2(_1804_),
    .B(_1805_),
    .ZN(_1806_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2706_ (.A1(_1751_),
    .A2(_1806_),
    .ZN(_1807_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2707_ (.A1(_1662_),
    .A2(_1698_),
    .ZN(_1808_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2708_ (.A1(_1662_),
    .A2(_1698_),
    .ZN(_1809_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2709_ (.A1(_1511_),
    .A2(_1808_),
    .B(_1809_),
    .ZN(_1810_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2710_ (.I(_1810_),
    .ZN(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2711_ (.A1(_1665_),
    .A2(_1671_),
    .ZN(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2712_ (.A1(_1665_),
    .A2(_1671_),
    .ZN(_1813_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2713_ (.A1(_1663_),
    .A2(_1812_),
    .B(_1813_),
    .ZN(_1814_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2714_ (.A1(_1674_),
    .A2(_1696_),
    .Z(_1815_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2715_ (.A1(_1672_),
    .A2(_1697_),
    .B(_1815_),
    .ZN(_1816_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2716_ (.I(_1668_),
    .Z(_1817_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2717_ (.A1(_1229_),
    .A2(_1817_),
    .B1(_1700_),
    .B2(_1266_),
    .ZN(_1818_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2718_ (.A1(_1682_),
    .A2(_1694_),
    .Z(_1819_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2719_ (.A1(_1680_),
    .A2(_1695_),
    .B(_1819_),
    .ZN(_1820_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _2720_ (.A1(_0991_),
    .A2(_1676_),
    .B1(_1683_),
    .B2(_1515_),
    .C(_1706_),
    .ZN(_1821_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2721_ (.A1(_1684_),
    .A2(_1693_),
    .Z(_1822_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2722_ (.A1(_1640_),
    .A2(_1765_),
    .ZN(_1823_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2723_ (.I(_1691_),
    .Z(_1824_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2724_ (.A1(_1685_),
    .A2(_1824_),
    .B(_1782_),
    .ZN(_1825_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2725_ (.A1(_1823_),
    .A2(_1825_),
    .Z(_1826_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2726_ (.A1(_1822_),
    .A2(_1826_),
    .Z(_1827_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2727_ (.A1(_1821_),
    .A2(_1827_),
    .ZN(_1828_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2728_ (.A1(_1820_),
    .A2(_1828_),
    .Z(_1829_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2729_ (.A1(_1818_),
    .A2(_1829_),
    .Z(_1830_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _2730_ (.A1(_1814_),
    .A2(_1816_),
    .A3(_1830_),
    .ZN(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2731_ (.A1(_1811_),
    .A2(_1831_),
    .Z(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2732_ (.I(_1699_),
    .ZN(_1833_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2733_ (.A1(_1833_),
    .A2(_1750_),
    .ZN(_1834_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2734_ (.A1(_1834_),
    .A2(_1832_),
    .Z(_1835_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2735_ (.A1(_1807_),
    .A2(_1835_),
    .ZN(_1836_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2736_ (.I(_1836_),
    .ZN(_1837_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2737_ (.A1(_1124_),
    .A2(_1309_),
    .Z(_1838_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2738_ (.A1(_1148_),
    .A2(_1718_),
    .Z(_1839_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2739_ (.A1(_1204_),
    .A2(_1224_),
    .B(_1180_),
    .ZN(_1840_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _2740_ (.A1(_0668_),
    .A2(_1258_),
    .B1(_1342_),
    .B2(_1270_),
    .C(_1206_),
    .ZN(_1841_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _2741_ (.A1(_1839_),
    .A2(_1840_),
    .B(_1841_),
    .C(_0580_),
    .ZN(_1842_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2742_ (.A1(_1170_),
    .A2(_1316_),
    .A3(_1523_),
    .B1(_1556_),
    .B2(_0668_),
    .ZN(_1843_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2743_ (.A1(_1238_),
    .A2(_1604_),
    .B(_1322_),
    .C(_1259_),
    .ZN(_1844_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2744_ (.A1(_1396_),
    .A2(_1843_),
    .B(_1844_),
    .ZN(_1845_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2745_ (.A1(_1569_),
    .A2(_1842_),
    .A3(_1845_),
    .Z(_1846_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2746_ (.A1(_1842_),
    .A2(_1845_),
    .B(_1574_),
    .ZN(_1847_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2747_ (.A1(_1846_),
    .A2(_1847_),
    .ZN(_1848_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2748_ (.A1(_1838_),
    .A2(_1491_),
    .B1(_1616_),
    .B2(_1848_),
    .ZN(_1849_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2749_ (.A1(_1664_),
    .A2(_1849_),
    .Z(_1850_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2750_ (.I(_1761_),
    .Z(_1851_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2751_ (.A1(_1590_),
    .A2(_1634_),
    .ZN(_1852_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2752_ (.A1(_1527_),
    .A2(_1547_),
    .B(_1852_),
    .ZN(_1853_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2753_ (.A1(_1630_),
    .A2(_1851_),
    .A3(_1853_),
    .ZN(_1854_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2754_ (.A1(_1679_),
    .A2(_1763_),
    .Z(_1855_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2755_ (.A1(_1854_),
    .A2(_1855_),
    .Z(_1856_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2756_ (.I(_1765_),
    .Z(_1857_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2757_ (.I(_1851_),
    .Z(_1858_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2758_ (.A1(_1857_),
    .A2(_1858_),
    .A3(_1853_),
    .A4(_1855_),
    .ZN(_1859_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2759_ (.A1(_1850_),
    .A2(_1856_),
    .B(_1859_),
    .ZN(_1860_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2760_ (.A1(_1775_),
    .A2(_1776_),
    .Z(_1861_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2761_ (.A1(_1860_),
    .A2(_1861_),
    .ZN(_1862_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2762_ (.A1(_1484_),
    .A2(_1488_),
    .ZN(_1863_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2763_ (.A1(_1087_),
    .A2(_1492_),
    .B1(_1863_),
    .B2(_1838_),
    .ZN(_1864_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2764_ (.A1(_1137_),
    .A2(_1502_),
    .ZN(_1865_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2765_ (.A1(_1364_),
    .A2(_1479_),
    .ZN(_1866_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2766_ (.A1(_1864_),
    .A2(_1865_),
    .Z(_1867_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2767_ (.A1(_1866_),
    .A2(_1867_),
    .ZN(_1868_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2768_ (.A1(_1864_),
    .A2(_1865_),
    .B(_1868_),
    .ZN(_1869_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2769_ (.A1(_1860_),
    .A2(_1861_),
    .Z(_1870_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2770_ (.A1(_1869_),
    .A2(_1870_),
    .ZN(_1871_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2771_ (.A1(_1862_),
    .A2(_1871_),
    .ZN(_1872_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2772_ (.A1(_1869_),
    .A2(_1870_),
    .Z(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2773_ (.A1(_1850_),
    .A2(_1856_),
    .ZN(_1874_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2774_ (.A1(_1530_),
    .A2(_1851_),
    .ZN(_1875_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2775_ (.A1(_1875_),
    .A2(_1853_),
    .Z(_1876_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2776_ (.A1(_1590_),
    .A2(_1713_),
    .B(_1609_),
    .ZN(_1877_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2777_ (.A1(_1609_),
    .A2(_1713_),
    .ZN(_1878_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2778_ (.A1(_1653_),
    .A2(_1877_),
    .B(_1878_),
    .ZN(_1879_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2779_ (.A1(_1731_),
    .A2(_1787_),
    .Z(_1880_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2780_ (.A1(_1879_),
    .A2(_1880_),
    .ZN(_1881_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2781_ (.A1(_1879_),
    .A2(_1880_),
    .ZN(_1882_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2782_ (.A1(_1876_),
    .A2(_1881_),
    .B(_1882_),
    .ZN(_1883_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2783_ (.A1(_1791_),
    .A2(_1793_),
    .Z(_1884_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2784_ (.A1(_1883_),
    .A2(_1884_),
    .ZN(_1885_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2785_ (.A1(_1883_),
    .A2(_1884_),
    .ZN(_1886_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2786_ (.A1(_1874_),
    .A2(_1885_),
    .B(_1886_),
    .ZN(_1887_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2787_ (.A1(_1781_),
    .A2(_1796_),
    .Z(_1888_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2788_ (.A1(_1887_),
    .A2(_1888_),
    .Z(_1889_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2789_ (.A1(_1887_),
    .A2(_1888_),
    .Z(_1890_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2790_ (.A1(_1873_),
    .A2(_1889_),
    .B(_1890_),
    .ZN(_1891_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2791_ (.A1(_1780_),
    .A2(_1800_),
    .ZN(_1892_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2792_ (.A1(_1891_),
    .A2(_1892_),
    .Z(_1893_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2793_ (.A1(_1891_),
    .A2(_1892_),
    .ZN(_1894_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2794_ (.A1(_1872_),
    .A2(_1893_),
    .B(_1894_),
    .ZN(_1895_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2795_ (.A1(_1779_),
    .A2(_1804_),
    .ZN(_1896_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2796_ (.A1(_1895_),
    .A2(_1896_),
    .ZN(_1897_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2797_ (.I(_1501_),
    .Z(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2798_ (.A1(_1127_),
    .A2(_0981_),
    .B(_1898_),
    .ZN(_1899_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2799_ (.A1(_1337_),
    .A2(_1489_),
    .ZN(_1900_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2800_ (.A1(_1865_),
    .A2(_1899_),
    .B(_1900_),
    .ZN(_1901_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2801_ (.A1(_1481_),
    .A2(_1478_),
    .Z(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2802_ (.A1(_1185_),
    .A2(_1705_),
    .ZN(_1903_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2803_ (.A1(_1901_),
    .A2(_1903_),
    .ZN(_1904_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2804_ (.A1(_1380_),
    .A2(_1902_),
    .A3(_1904_),
    .ZN(_1905_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2805_ (.A1(_1185_),
    .A2(_1706_),
    .A3(_1901_),
    .B(_1905_),
    .ZN(_1906_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2806_ (.A1(_0525_),
    .A2(_1619_),
    .B(_1211_),
    .C(_1393_),
    .ZN(_1907_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2807_ (.A1(_1389_),
    .A2(_1394_),
    .B(_1907_),
    .C(_1355_),
    .ZN(_1908_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2808_ (.A1(_1220_),
    .A2(_1402_),
    .B1(_1550_),
    .B2(_0470_),
    .ZN(_1909_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2809_ (.A1(_1207_),
    .A2(_1909_),
    .B(_1360_),
    .ZN(_1910_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2810_ (.A1(_1207_),
    .A2(_1354_),
    .A3(_1244_),
    .ZN(_1911_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2811_ (.A1(_1178_),
    .A2(_1346_),
    .B1(_1251_),
    .B2(_1238_),
    .C(_1319_),
    .ZN(_1912_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2812_ (.A1(_1236_),
    .A2(_1912_),
    .ZN(_1913_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2813_ (.A1(_1908_),
    .A2(_1910_),
    .B1(_1911_),
    .B2(_1913_),
    .ZN(_1914_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2814_ (.A1(_1636_),
    .A2(_1914_),
    .Z(_1915_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2815_ (.A1(_1337_),
    .A2(_1501_),
    .Z(_1916_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2816_ (.A1(_1514_),
    .A2(_1915_),
    .B(_1916_),
    .ZN(_1917_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2817_ (.A1(_1506_),
    .A2(_1917_),
    .Z(_1918_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2818_ (.A1(_1725_),
    .A2(_1726_),
    .Z(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2819_ (.A1(_1547_),
    .A2(_0033_),
    .ZN(_0034_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _2820_ (.A1(_1782_),
    .A2(_0034_),
    .B(_1848_),
    .C(_1531_),
    .ZN(_0035_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2821_ (.A1(_1615_),
    .A2(_1849_),
    .ZN(_0036_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2822_ (.A1(_0035_),
    .A2(_0036_),
    .Z(_0037_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2823_ (.A1(_0035_),
    .A2(_0036_),
    .ZN(_0038_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2824_ (.A1(_1918_),
    .A2(_0037_),
    .B(_0038_),
    .ZN(_0039_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2825_ (.A1(_1866_),
    .A2(_1867_),
    .ZN(_0040_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2826_ (.A1(_0039_),
    .A2(_0040_),
    .Z(_0041_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2827_ (.A1(_1906_),
    .A2(_0041_),
    .ZN(_0042_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2828_ (.A1(_1918_),
    .A2(_0037_),
    .Z(_0043_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2829_ (.I(_0043_),
    .ZN(_0044_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2830_ (.A1(_1846_),
    .A2(_1847_),
    .Z(_0045_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _2831_ (.A1(_1548_),
    .A2(_0033_),
    .B1(_0045_),
    .B2(_1532_),
    .C(_1737_),
    .ZN(_0046_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2832_ (.A1(_0035_),
    .A2(_0046_),
    .Z(_0047_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2833_ (.A1(_1607_),
    .A2(_1608_),
    .Z(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2834_ (.A1(_0048_),
    .A2(_1527_),
    .B(_1579_),
    .ZN(_0049_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2835_ (.A1(_1785_),
    .A2(_1878_),
    .A3(_0049_),
    .Z(_0050_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2836_ (.A1(_1878_),
    .A2(_0049_),
    .B(_1785_),
    .ZN(_0051_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2837_ (.A1(_1563_),
    .A2(_1565_),
    .Z(_0052_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2838_ (.A1(_1725_),
    .A2(_1726_),
    .B(_1587_),
    .ZN(_0053_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2839_ (.I(_0053_),
    .Z(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2840_ (.I(_1591_),
    .Z(_0055_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2841_ (.A1(_1580_),
    .A2(_0033_),
    .B(_0055_),
    .ZN(_0056_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2842_ (.A1(_0052_),
    .A2(_0054_),
    .B1(_0056_),
    .B2(_1635_),
    .ZN(_0057_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2843_ (.A1(_0050_),
    .A2(_0051_),
    .B(_0057_),
    .ZN(_0058_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2844_ (.A1(_0050_),
    .A2(_0057_),
    .A3(_0051_),
    .ZN(_0059_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2845_ (.A1(_0047_),
    .A2(_0058_),
    .B(_0059_),
    .ZN(_0060_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2846_ (.A1(_1876_),
    .A2(_1881_),
    .ZN(_0061_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2847_ (.A1(_0060_),
    .A2(_0061_),
    .ZN(_0062_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2848_ (.A1(_0060_),
    .A2(_0061_),
    .Z(_0064_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2849_ (.A1(_0044_),
    .A2(_0062_),
    .B(_0064_),
    .ZN(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _2850_ (.A1(_1883_),
    .A2(_1884_),
    .A3(_1874_),
    .ZN(_0066_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2851_ (.A1(_0065_),
    .A2(_0066_),
    .ZN(_0067_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2852_ (.A1(_0065_),
    .A2(_0066_),
    .ZN(_0068_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2853_ (.A1(_0042_),
    .A2(_0067_),
    .B(_0068_),
    .ZN(_0069_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2854_ (.A1(_1873_),
    .A2(_1889_),
    .Z(_0070_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2855_ (.A1(_0069_),
    .A2(_0070_),
    .Z(_0071_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2856_ (.A1(_0039_),
    .A2(_0040_),
    .ZN(_0072_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2857_ (.A1(_1906_),
    .A2(_0041_),
    .B(_0072_),
    .ZN(_0073_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2858_ (.A1(_0069_),
    .A2(_0070_),
    .ZN(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2859_ (.A1(_0073_),
    .A2(_0075_),
    .ZN(_0076_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2860_ (.A1(_1872_),
    .A2(_1893_),
    .Z(_0077_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2861_ (.A1(_0071_),
    .A2(_0076_),
    .B(_0077_),
    .ZN(_0078_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2862_ (.A1(_1897_),
    .A2(_0078_),
    .ZN(_0079_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2863_ (.A1(_1751_),
    .A2(_1806_),
    .Z(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2864_ (.A1(_1895_),
    .A2(_1896_),
    .ZN(_0081_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2865_ (.A1(_0080_),
    .A2(_0081_),
    .ZN(_0082_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2866_ (.A1(_0079_),
    .A2(_0082_),
    .Z(_0083_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2867_ (.A1(_1137_),
    .A2(_1506_),
    .ZN(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2868_ (.A1(_1615_),
    .A2(_1706_),
    .B(_1903_),
    .ZN(_0086_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2869_ (.A1(_1363_),
    .A2(_1490_),
    .ZN(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2870_ (.A1(_0086_),
    .A2(_0087_),
    .ZN(_0088_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2871_ (.A1(_1020_),
    .A2(_1398_),
    .Z(_0089_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2872_ (.I(_0089_),
    .Z(_0090_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2873_ (.A1(_0090_),
    .A2(_1902_),
    .ZN(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2874_ (.I(_0091_),
    .ZN(_0092_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2875_ (.A1(_0084_),
    .A2(_0088_),
    .Z(_0093_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2876_ (.A1(_0092_),
    .A2(_0093_),
    .ZN(_0094_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2877_ (.A1(_0084_),
    .A2(_0088_),
    .B(_0094_),
    .ZN(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2878_ (.A1(_1642_),
    .A2(_1851_),
    .B(_1732_),
    .ZN(_0097_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2879_ (.A1(_1574_),
    .A2(_1914_),
    .Z(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2880_ (.A1(_1630_),
    .A2(_0098_),
    .ZN(_0099_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2881_ (.A1(_0097_),
    .A2(_0099_),
    .Z(_0100_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2882_ (.A1(_1506_),
    .A2(_1917_),
    .ZN(_0101_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2883_ (.A1(_1918_),
    .A2(_0100_),
    .A3(_0101_),
    .ZN(_0102_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2884_ (.A1(_1619_),
    .A2(_1557_),
    .ZN(_0103_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2885_ (.A1(_1174_),
    .A2(_0103_),
    .B(_1334_),
    .ZN(_0104_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2886_ (.A1(_1323_),
    .A2(_1403_),
    .ZN(_0105_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2887_ (.A1(_1170_),
    .A2(_1523_),
    .A3(_0105_),
    .B1(_1215_),
    .B2(_1421_),
    .ZN(_0106_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2888_ (.A1(_1406_),
    .A2(_1387_),
    .B(_1236_),
    .ZN(_0108_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2889_ (.A1(_1331_),
    .A2(_1202_),
    .B1(_1301_),
    .B2(_1389_),
    .ZN(_0109_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _2890_ (.A1(_1411_),
    .A2(_0106_),
    .B1(_0108_),
    .B2(_1283_),
    .C1(_0109_),
    .C2(_1194_),
    .ZN(_0110_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _2891_ (.A1(_1636_),
    .A2(_0104_),
    .A3(_0110_),
    .Z(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2892_ (.I(_1516_),
    .Z(_0112_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2893_ (.A1(_0104_),
    .A2(_0110_),
    .B(_0112_),
    .ZN(_0113_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2894_ (.A1(_0111_),
    .A2(_0113_),
    .ZN(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2895_ (.A1(_1363_),
    .A2(_1504_),
    .Z(_0115_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2896_ (.A1(_1514_),
    .A2(_0114_),
    .B(_0115_),
    .ZN(_0116_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2897_ (.A1(_1704_),
    .A2(_0116_),
    .ZN(_0117_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2898_ (.A1(_1505_),
    .A2(_1917_),
    .A3(_0100_),
    .Z(_0119_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2899_ (.A1(_0117_),
    .A2(_0119_),
    .ZN(_0120_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2900_ (.A1(_0102_),
    .A2(_0120_),
    .ZN(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2901_ (.A1(_1380_),
    .A2(_1902_),
    .ZN(_0122_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2902_ (.A1(_0122_),
    .A2(_1904_),
    .Z(_0123_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2903_ (.A1(_0121_),
    .A2(_0123_),
    .Z(_0124_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2904_ (.A1(_0121_),
    .A2(_0123_),
    .ZN(_0125_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2905_ (.A1(_0095_),
    .A2(_0124_),
    .B(_0125_),
    .ZN(_0126_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2906_ (.A1(_0097_),
    .A2(_0099_),
    .ZN(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2907_ (.A1(_0100_),
    .A2(_0127_),
    .ZN(_0128_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2908_ (.A1(_1759_),
    .A2(_1760_),
    .B(_1587_),
    .ZN(_0130_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2909_ (.A1(_1759_),
    .A2(_1760_),
    .Z(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2910_ (.I0(_0130_),
    .I1(_0131_),
    .S(_1733_),
    .Z(_0132_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2911_ (.A1(_1734_),
    .A2(_1858_),
    .B1(_0132_),
    .B2(_1581_),
    .ZN(_0133_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2912_ (.I0(_0055_),
    .I1(_0052_),
    .S(_0053_),
    .Z(_0134_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2913_ (.A1(_1635_),
    .A2(_0134_),
    .Z(_0135_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2914_ (.A1(_0133_),
    .A2(_0135_),
    .ZN(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2915_ (.A1(_0133_),
    .A2(_0135_),
    .Z(_0137_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2916_ (.A1(_0128_),
    .A2(_0136_),
    .B(_0137_),
    .ZN(_0138_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2917_ (.A1(_0050_),
    .A2(_0051_),
    .ZN(_0139_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2918_ (.A1(_0057_),
    .A2(_0139_),
    .A3(_0047_),
    .Z(_0141_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2919_ (.A1(_0138_),
    .A2(_0141_),
    .ZN(_0142_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2920_ (.A1(_0117_),
    .A2(_0119_),
    .Z(_0143_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2921_ (.A1(_0128_),
    .A2(_0136_),
    .Z(_0144_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2922_ (.A1(_0137_),
    .A2(_0144_),
    .B(_0141_),
    .ZN(_0145_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2923_ (.A1(_0142_),
    .A2(_0143_),
    .B(_0145_),
    .ZN(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2924_ (.A1(_0043_),
    .A2(_0062_),
    .Z(_0147_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2925_ (.A1(_0146_),
    .A2(_0147_),
    .Z(_0148_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2926_ (.A1(_0095_),
    .A2(_0124_),
    .Z(_0149_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2927_ (.A1(_0146_),
    .A2(_0147_),
    .ZN(_0150_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2928_ (.A1(_0148_),
    .A2(_0149_),
    .B(_0150_),
    .ZN(_0152_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2929_ (.A1(_0042_),
    .A2(_0067_),
    .ZN(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2930_ (.A1(_0152_),
    .A2(_0153_),
    .ZN(_0154_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2931_ (.A1(_0152_),
    .A2(_0153_),
    .Z(_0155_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2932_ (.A1(_0126_),
    .A2(_0154_),
    .B(_0155_),
    .ZN(_0156_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2933_ (.A1(_0073_),
    .A2(_0075_),
    .Z(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2934_ (.A1(_0156_),
    .A2(_0157_),
    .Z(_0158_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2935_ (.A1(_1484_),
    .A2(_1669_),
    .Z(_0159_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2936_ (.A1(_1380_),
    .A2(_0159_),
    .ZN(_0160_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2937_ (.A1(_1265_),
    .A2(_1664_),
    .ZN(_0161_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2938_ (.A1(_0981_),
    .A2(_1228_),
    .B(_1898_),
    .ZN(_0163_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2939_ (.A1(_0084_),
    .A2(_0163_),
    .ZN(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2940_ (.A1(_1381_),
    .A2(_1490_),
    .B(_0164_),
    .ZN(_0165_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2941_ (.A1(_1415_),
    .A2(_1666_),
    .ZN(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2942_ (.A1(_0161_),
    .A2(_0165_),
    .Z(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2943_ (.A1(_0166_),
    .A2(_0167_),
    .Z(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2944_ (.A1(_0161_),
    .A2(_0165_),
    .B(_0168_),
    .ZN(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2945_ (.A1(_0111_),
    .A2(_0113_),
    .Z(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2946_ (.A1(_1548_),
    .A2(_0045_),
    .B(_1653_),
    .ZN(_0171_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2947_ (.A1(_1715_),
    .A2(_0170_),
    .A3(_0171_),
    .ZN(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2948_ (.A1(_1707_),
    .A2(_0116_),
    .Z(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2949_ (.I(_1762_),
    .Z(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2950_ (.A1(_1406_),
    .A2(_0767_),
    .A3(_1247_),
    .B(_1298_),
    .ZN(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2951_ (.A1(_1394_),
    .A2(_1277_),
    .B1(_1392_),
    .B2(_1648_),
    .C(_1355_),
    .ZN(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2952_ (.A1(_1241_),
    .A2(_0176_),
    .B(_0177_),
    .C(_1411_),
    .ZN(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2953_ (.A1(_1220_),
    .A2(_1389_),
    .B(_1291_),
    .C(_1370_),
    .ZN(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2954_ (.A1(_1403_),
    .A2(_1367_),
    .B1(_1250_),
    .B2(_1406_),
    .ZN(_0180_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2955_ (.A1(_1553_),
    .A2(_0179_),
    .B1(_0180_),
    .B2(_1644_),
    .ZN(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _2956_ (.A1(_0112_),
    .A2(_0178_),
    .A3(_0181_),
    .Z(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2957_ (.A1(_0178_),
    .A2(_0181_),
    .B(_0112_),
    .ZN(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2958_ (.A1(_0182_),
    .A2(_0183_),
    .ZN(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2959_ (.A1(_1379_),
    .A2(_1492_),
    .ZN(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2960_ (.A1(_1514_),
    .A2(_0185_),
    .B(_0186_),
    .ZN(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2961_ (.A1(_0175_),
    .A2(_0187_),
    .Z(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2962_ (.A1(_1707_),
    .A2(_0116_),
    .A3(_0172_),
    .Z(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2963_ (.A1(_0188_),
    .A2(_0189_),
    .ZN(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2964_ (.A1(_0172_),
    .A2(_0174_),
    .B(_0190_),
    .ZN(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2965_ (.A1(_0092_),
    .A2(_0093_),
    .Z(_0192_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2966_ (.A1(_0191_),
    .A2(_0192_),
    .ZN(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2967_ (.A1(_0191_),
    .A2(_0192_),
    .ZN(_0194_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2968_ (.A1(_0169_),
    .A2(_0193_),
    .B(_0194_),
    .ZN(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2969_ (.I(_0196_),
    .ZN(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2970_ (.A1(_1630_),
    .A2(_0170_),
    .ZN(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2971_ (.A1(_0171_),
    .A2(_0198_),
    .Z(_0199_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2972_ (.I(_0199_),
    .ZN(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2973_ (.A1(_1587_),
    .A2(_1846_),
    .A3(_1847_),
    .ZN(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2974_ (.I0(_1786_),
    .I1(_1543_),
    .S(_0201_),
    .Z(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2975_ (.A1(_1618_),
    .A2(_0201_),
    .B1(_0202_),
    .B2(_1734_),
    .ZN(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2976_ (.A1(_0055_),
    .A2(_0132_),
    .Z(_0204_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2977_ (.A1(_0203_),
    .A2(_0204_),
    .Z(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2978_ (.A1(_0203_),
    .A2(_0204_),
    .ZN(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2979_ (.A1(_0200_),
    .A2(_0205_),
    .B(_0207_),
    .ZN(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2980_ (.A1(_0128_),
    .A2(_0136_),
    .ZN(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2981_ (.A1(_0208_),
    .A2(_0209_),
    .Z(_0210_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2982_ (.A1(_0188_),
    .A2(_0189_),
    .Z(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2983_ (.A1(_0208_),
    .A2(_0209_),
    .ZN(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2984_ (.A1(_0210_),
    .A2(_0211_),
    .B(_0212_),
    .ZN(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2985_ (.A1(_0142_),
    .A2(_0143_),
    .Z(_0214_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2986_ (.A1(_0213_),
    .A2(_0214_),
    .Z(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2987_ (.A1(_0169_),
    .A2(_0193_),
    .ZN(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2988_ (.A1(_0210_),
    .A2(_0211_),
    .Z(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2989_ (.A1(_0212_),
    .A2(_0218_),
    .B(_0214_),
    .ZN(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2990_ (.A1(_0215_),
    .A2(_0216_),
    .B(_0219_),
    .ZN(_0220_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2991_ (.A1(_0148_),
    .A2(_0149_),
    .Z(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2992_ (.A1(_0220_),
    .A2(_0221_),
    .ZN(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2993_ (.A1(_0220_),
    .A2(_0221_),
    .ZN(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2994_ (.A1(_0197_),
    .A2(_0222_),
    .B(_0223_),
    .ZN(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2995_ (.A1(_0126_),
    .A2(_0154_),
    .Z(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2996_ (.A1(_0224_),
    .A2(_0225_),
    .ZN(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2997_ (.A1(_0224_),
    .A2(_0225_),
    .ZN(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2998_ (.A1(_0160_),
    .A2(_0226_),
    .B(_0227_),
    .ZN(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2999_ (.A1(_0158_),
    .A2(_0229_),
    .Z(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3000_ (.I(_0230_),
    .Z(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3001_ (.A1(_0071_),
    .A2(_0076_),
    .ZN(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3002_ (.A1(_0232_),
    .A2(_0077_),
    .ZN(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3003_ (.A1(_0156_),
    .A2(_0157_),
    .Z(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3004_ (.A1(_0233_),
    .A2(_0234_),
    .Z(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3005_ (.I(_0233_),
    .ZN(_0236_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3006_ (.A1(_0158_),
    .A2(_0229_),
    .B(_0234_),
    .ZN(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3007_ (.A1(_0236_),
    .A2(_0237_),
    .ZN(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3008_ (.A1(_0231_),
    .A2(_0235_),
    .B(_0238_),
    .ZN(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3009_ (.I(_0115_),
    .Z(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3010_ (.A1(_1311_),
    .A2(_0241_),
    .ZN(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3011_ (.I(_0186_),
    .Z(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3012_ (.A1(_0129_),
    .A2(_1442_),
    .Z(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3013_ (.A1(_0244_),
    .A2(_1493_),
    .ZN(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3014_ (.A1(_1786_),
    .A2(_0245_),
    .Z(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3015_ (.A1(_0244_),
    .A2(_1493_),
    .A3(_1786_),
    .ZN(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3016_ (.A1(_0243_),
    .A2(_0246_),
    .B(_0247_),
    .ZN(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3017_ (.I(_1898_),
    .Z(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3018_ (.A1(_1364_),
    .A2(_0249_),
    .ZN(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3019_ (.I(_1916_),
    .Z(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3020_ (.I0(_1365_),
    .I1(_0251_),
    .S(_0252_),
    .Z(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3021_ (.A1(_0175_),
    .A2(_0253_),
    .Z(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3022_ (.A1(_0248_),
    .A2(_0254_),
    .Z(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3023_ (.I(_1676_),
    .Z(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3024_ (.A1(_0248_),
    .A2(_0254_),
    .ZN(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3025_ (.A1(_1429_),
    .A2(_0256_),
    .B(_0257_),
    .ZN(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3026_ (.A1(_0242_),
    .A2(_0255_),
    .B(_0258_),
    .ZN(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3027_ (.I(_0201_),
    .Z(_0260_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3028_ (.I(_0130_),
    .Z(_0262_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3029_ (.I0(_0262_),
    .I1(_0131_),
    .S(_0260_),
    .Z(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3030_ (.A1(_1580_),
    .A2(_1528_),
    .ZN(_0264_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3031_ (.A1(_1858_),
    .A2(_0260_),
    .B1(_0263_),
    .B2(_0264_),
    .ZN(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3032_ (.I(_1736_),
    .Z(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3033_ (.A1(_0266_),
    .A2(_1728_),
    .ZN(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _3034_ (.A1(_1736_),
    .A2(_0182_),
    .A3(_0183_),
    .ZN(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3035_ (.I0(_0131_),
    .I1(_0130_),
    .S(_0268_),
    .Z(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3036_ (.A1(_0267_),
    .A2(_0269_),
    .Z(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3037_ (.A1(_0265_),
    .A2(_0270_),
    .ZN(_0271_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3038_ (.A1(_0186_),
    .A2(_0246_),
    .Z(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3039_ (.A1(_0265_),
    .A2(_0270_),
    .ZN(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3040_ (.A1(_0271_),
    .A2(_0273_),
    .B(_0274_),
    .ZN(_0275_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3041_ (.A1(_0182_),
    .A2(_0183_),
    .Z(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3042_ (.A1(_0262_),
    .A2(_0276_),
    .B1(_0269_),
    .B2(_0054_),
    .ZN(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3043_ (.A1(_1736_),
    .A2(_0111_),
    .A3(_0113_),
    .ZN(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3044_ (.I0(_0278_),
    .I1(_0170_),
    .S(_0054_),
    .Z(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3045_ (.A1(_0264_),
    .A2(_0279_),
    .Z(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3046_ (.A1(_0277_),
    .A2(_0280_),
    .ZN(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3047_ (.I(_1579_),
    .Z(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3048_ (.A1(_0282_),
    .A2(_1678_),
    .B1(_0185_),
    .B2(_1549_),
    .ZN(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3049_ (.A1(_1428_),
    .A2(_0249_),
    .ZN(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3050_ (.A1(_0281_),
    .A2(_0284_),
    .A3(_0285_),
    .Z(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3051_ (.A1(_0275_),
    .A2(_0286_),
    .Z(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3052_ (.A1(_0242_),
    .A2(_0255_),
    .Z(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3053_ (.A1(_0275_),
    .A2(_0286_),
    .ZN(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3054_ (.A1(_0287_),
    .A2(_0288_),
    .B(_0289_),
    .ZN(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3055_ (.A1(_0284_),
    .A2(_0285_),
    .Z(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3056_ (.A1(_0284_),
    .A2(_0285_),
    .ZN(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _3057_ (.A1(_0281_),
    .A2(_0291_),
    .A3(_0292_),
    .B1(_0280_),
    .B2(_0277_),
    .ZN(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3058_ (.I(_0114_),
    .Z(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _3059_ (.A1(_0282_),
    .A2(_1528_),
    .A3(_0279_),
    .B1(_0295_),
    .B2(_0267_),
    .ZN(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3060_ (.A1(_1687_),
    .A2(_1618_),
    .ZN(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3061_ (.A1(_0282_),
    .A2(_1527_),
    .A3(_1915_),
    .ZN(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3062_ (.A1(_1714_),
    .A2(_0098_),
    .B(_1687_),
    .ZN(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _3063_ (.A1(_0297_),
    .A2(_0298_),
    .A3(_0299_),
    .Z(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3064_ (.A1(_0298_),
    .A2(_0299_),
    .B(_0297_),
    .ZN(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3065_ (.A1(_0300_),
    .A2(_0301_),
    .Z(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3066_ (.A1(_1548_),
    .A2(_0114_),
    .B(_0055_),
    .ZN(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3067_ (.A1(_1414_),
    .A2(_1898_),
    .ZN(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3068_ (.I(_0304_),
    .ZN(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3069_ (.A1(_0303_),
    .A2(_0306_),
    .Z(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _3070_ (.A1(_0296_),
    .A2(_0302_),
    .A3(_0307_),
    .ZN(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3071_ (.A1(_0293_),
    .A2(_0308_),
    .ZN(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3072_ (.A1(_1338_),
    .A2(_0241_),
    .ZN(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3073_ (.A1(_0175_),
    .A2(_0253_),
    .B(_0310_),
    .ZN(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3074_ (.A1(_1310_),
    .A2(_1504_),
    .ZN(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3075_ (.I0(_1311_),
    .I1(_0312_),
    .S(_0252_),
    .Z(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3076_ (.A1(_1707_),
    .A2(_0313_),
    .Z(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3077_ (.A1(_0291_),
    .A2(_0314_),
    .ZN(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3078_ (.A1(_0311_),
    .A2(_0315_),
    .Z(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3079_ (.A1(_0309_),
    .A2(_0317_),
    .ZN(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3080_ (.A1(_0290_),
    .A2(_0318_),
    .ZN(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3081_ (.A1(_0290_),
    .A2(_0318_),
    .Z(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3082_ (.A1(_0259_),
    .A2(_0319_),
    .B(_0320_),
    .ZN(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3083_ (.I(_0311_),
    .ZN(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3084_ (.I(_0291_),
    .ZN(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3085_ (.A1(_0323_),
    .A2(_0314_),
    .ZN(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3086_ (.A1(_0322_),
    .A2(_0315_),
    .B(_0324_),
    .ZN(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3087_ (.A1(_1443_),
    .A2(_1666_),
    .ZN(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3088_ (.A1(_1414_),
    .A2(_1675_),
    .B(_1507_),
    .ZN(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3089_ (.A1(_0326_),
    .A2(_0328_),
    .ZN(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3090_ (.A1(_0325_),
    .A2(_0329_),
    .Z(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3091_ (.A1(_0293_),
    .A2(_0308_),
    .ZN(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3092_ (.A1(_0309_),
    .A2(_0317_),
    .B(_0331_),
    .ZN(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3093_ (.A1(_0300_),
    .A2(_0301_),
    .B(_0296_),
    .ZN(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3094_ (.A1(_0296_),
    .A2(_0300_),
    .A3(_0301_),
    .ZN(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3095_ (.A1(_0333_),
    .A2(_0307_),
    .B(_0334_),
    .ZN(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3096_ (.I(_0098_),
    .Z(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3097_ (.A1(_1642_),
    .A2(_0336_),
    .B(_1635_),
    .ZN(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3098_ (.A1(_1715_),
    .A2(_0276_),
    .ZN(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3099_ (.A1(_0337_),
    .A2(_0339_),
    .Z(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3100_ (.A1(_1687_),
    .A2(_1714_),
    .A3(_0098_),
    .ZN(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3101_ (.A1(_0297_),
    .A2(_0299_),
    .B(_0341_),
    .ZN(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3102_ (.A1(_1734_),
    .A2(_0202_),
    .Z(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3103_ (.A1(_0342_),
    .A2(_0343_),
    .Z(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3104_ (.A1(_0340_),
    .A2(_0344_),
    .Z(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3105_ (.A1(_0335_),
    .A2(_0345_),
    .ZN(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3106_ (.A1(_1338_),
    .A2(_0249_),
    .ZN(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3107_ (.A1(_1838_),
    .A2(_0347_),
    .B1(_0313_),
    .B2(_1704_),
    .ZN(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3108_ (.A1(_0303_),
    .A2(_0304_),
    .ZN(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3109_ (.A1(_0089_),
    .A2(_1492_),
    .ZN(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3110_ (.I0(_1310_),
    .I1(_0312_),
    .S(_0351_),
    .Z(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3111_ (.A1(_1762_),
    .A2(_0352_),
    .ZN(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3112_ (.A1(_0350_),
    .A2(_0353_),
    .Z(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3113_ (.A1(_0348_),
    .A2(_0354_),
    .Z(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3114_ (.A1(_0346_),
    .A2(_0355_),
    .Z(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3115_ (.A1(_0332_),
    .A2(_0356_),
    .Z(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3116_ (.A1(_0330_),
    .A2(_0357_),
    .Z(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3117_ (.A1(_0325_),
    .A2(_0329_),
    .ZN(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3118_ (.A1(_0332_),
    .A2(_0356_),
    .Z(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3119_ (.A1(_0330_),
    .A2(_0357_),
    .B(_0361_),
    .ZN(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3120_ (.I(_0348_),
    .ZN(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3121_ (.A1(_0350_),
    .A2(_0353_),
    .ZN(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3122_ (.A1(_0363_),
    .A2(_0354_),
    .B(_0364_),
    .ZN(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3123_ (.A1(_1428_),
    .A2(_1667_),
    .ZN(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3124_ (.A1(_0326_),
    .A2(_0328_),
    .Z(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3125_ (.I0(_1265_),
    .I1(_1704_),
    .S(_1664_),
    .Z(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3126_ (.A1(_1399_),
    .A2(_1675_),
    .ZN(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3127_ (.A1(_0368_),
    .A2(_0369_),
    .Z(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3128_ (.A1(_0367_),
    .A2(_0370_),
    .ZN(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3129_ (.A1(_0366_),
    .A2(_0372_),
    .Z(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3130_ (.A1(_0365_),
    .A2(_0373_),
    .Z(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3131_ (.A1(_0365_),
    .A2(_0373_),
    .ZN(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3132_ (.A1(_0374_),
    .A2(_0375_),
    .ZN(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3133_ (.A1(_0335_),
    .A2(_0345_),
    .ZN(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3134_ (.A1(_0346_),
    .A2(_0355_),
    .B(_0377_),
    .ZN(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3135_ (.A1(_0342_),
    .A2(_0343_),
    .Z(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3136_ (.A1(_0340_),
    .A2(_0344_),
    .B(_0379_),
    .ZN(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3137_ (.A1(_0199_),
    .A2(_0205_),
    .Z(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3138_ (.A1(_0380_),
    .A2(_0381_),
    .Z(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3139_ (.A1(_0090_),
    .A2(_0312_),
    .B1(_0352_),
    .B2(_0175_),
    .ZN(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3140_ (.A1(_0337_),
    .A2(_0339_),
    .ZN(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3141_ (.A1(_1762_),
    .A2(_0187_),
    .Z(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3142_ (.A1(_0385_),
    .A2(_0386_),
    .ZN(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3143_ (.A1(_0384_),
    .A2(_0387_),
    .Z(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3144_ (.A1(_0383_),
    .A2(_0388_),
    .Z(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3145_ (.A1(_0378_),
    .A2(_0389_),
    .ZN(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3146_ (.A1(_0376_),
    .A2(_0390_),
    .ZN(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3147_ (.A1(_0359_),
    .A2(_0362_),
    .A3(_0391_),
    .Z(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3148_ (.A1(_0321_),
    .A2(_0358_),
    .A3(_0392_),
    .ZN(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3149_ (.I(_1700_),
    .Z(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3150_ (.I(_0395_),
    .Z(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3151_ (.A1(_1444_),
    .A2(_0396_),
    .ZN(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3152_ (.A1(_0321_),
    .A2(_0358_),
    .ZN(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3153_ (.A1(_0398_),
    .A2(_0392_),
    .ZN(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3154_ (.A1(_0397_),
    .A2(_0399_),
    .ZN(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3155_ (.A1(_0394_),
    .A2(_0400_),
    .ZN(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3156_ (.I(_0396_),
    .Z(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3157_ (.A1(_1430_),
    .A2(_0402_),
    .ZN(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3158_ (.A1(_0362_),
    .A2(_0391_),
    .ZN(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _3159_ (.A1(_0325_),
    .A2(_0329_),
    .A3(_0405_),
    .B1(_0391_),
    .B2(_0362_),
    .ZN(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3160_ (.I(_0374_),
    .ZN(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3161_ (.A1(_0378_),
    .A2(_0389_),
    .ZN(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3162_ (.A1(_0376_),
    .A2(_0390_),
    .B(_0408_),
    .ZN(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3163_ (.A1(_0380_),
    .A2(_0381_),
    .ZN(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3164_ (.A1(_0383_),
    .A2(_0388_),
    .B(_0410_),
    .ZN(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3165_ (.A1(_0210_),
    .A2(_0211_),
    .A3(_0411_),
    .Z(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3166_ (.A1(_1428_),
    .A2(_1667_),
    .A3(_0372_),
    .ZN(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3167_ (.A1(_0367_),
    .A2(_0370_),
    .B(_0413_),
    .ZN(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3168_ (.A1(_0385_),
    .A2(_0386_),
    .ZN(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3169_ (.A1(_0384_),
    .A2(_0387_),
    .B(_0416_),
    .ZN(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3170_ (.A1(_0166_),
    .A2(_0167_),
    .Z(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3171_ (.A1(_0417_),
    .A2(_0418_),
    .Z(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3172_ (.A1(_0414_),
    .A2(_0419_),
    .Z(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3173_ (.A1(_0412_),
    .A2(_0420_),
    .Z(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3174_ (.A1(_0409_),
    .A2(_0421_),
    .Z(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3175_ (.A1(_0407_),
    .A2(_0422_),
    .Z(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _3176_ (.A1(_0406_),
    .A2(_0423_),
    .Z(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3177_ (.A1(_0403_),
    .A2(_0424_),
    .Z(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3178_ (.A1(_1430_),
    .A2(_0402_),
    .Z(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3179_ (.A1(_0406_),
    .A2(_0423_),
    .ZN(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3180_ (.A1(_0406_),
    .A2(_0423_),
    .ZN(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3181_ (.A1(_0427_),
    .A2(_0428_),
    .B(_0429_),
    .ZN(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3182_ (.A1(_1416_),
    .A2(_0396_),
    .ZN(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3183_ (.A1(_0409_),
    .A2(_0421_),
    .Z(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3184_ (.A1(_0407_),
    .A2(_0422_),
    .B(_0432_),
    .ZN(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3185_ (.A1(_0417_),
    .A2(_0418_),
    .ZN(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3186_ (.A1(_0417_),
    .A2(_0418_),
    .ZN(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3187_ (.A1(_0414_),
    .A2(_0434_),
    .B(_0435_),
    .ZN(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3188_ (.A1(_0210_),
    .A2(_0211_),
    .ZN(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _3189_ (.A1(_0218_),
    .A2(_0411_),
    .A3(_0438_),
    .B1(_0412_),
    .B2(_0420_),
    .ZN(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3190_ (.A1(_0215_),
    .A2(_0216_),
    .Z(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3191_ (.A1(_0439_),
    .A2(_0440_),
    .Z(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3192_ (.A1(_0436_),
    .A2(_0441_),
    .ZN(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3193_ (.A1(_0431_),
    .A2(_0433_),
    .A3(_0442_),
    .Z(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3194_ (.A1(_0401_),
    .A2(_0425_),
    .B1(_0430_),
    .B2(_0443_),
    .ZN(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3195_ (.A1(_0406_),
    .A2(_0423_),
    .Z(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _3196_ (.A1(_0403_),
    .A2(_0424_),
    .B(_0443_),
    .C(_0445_),
    .ZN(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _3197_ (.A1(_0431_),
    .A2(_0433_),
    .A3(_0442_),
    .ZN(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3198_ (.A1(_0427_),
    .A2(_0428_),
    .B(_0447_),
    .C(_0429_),
    .ZN(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3199_ (.A1(_0401_),
    .A2(_0425_),
    .B(_0449_),
    .ZN(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3200_ (.I(_0243_),
    .ZN(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3201_ (.I(_0351_),
    .Z(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3202_ (.I0(_0090_),
    .I1(_0452_),
    .S(_0243_),
    .Z(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3203_ (.A1(_0252_),
    .A2(_0453_),
    .ZN(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3204_ (.A1(_0090_),
    .A2(_0451_),
    .B(_0454_),
    .ZN(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3205_ (.A1(_1838_),
    .A2(_1493_),
    .ZN(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3206_ (.A1(_0456_),
    .A2(_0241_),
    .B(_0242_),
    .ZN(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3207_ (.I(_0457_),
    .ZN(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3208_ (.A1(_0455_),
    .A2(_0458_),
    .Z(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3209_ (.I(_1915_),
    .Z(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3210_ (.A1(_0266_),
    .A2(_1848_),
    .ZN(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3211_ (.A1(_0266_),
    .A2(_0336_),
    .B(_0260_),
    .ZN(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3212_ (.A1(_0461_),
    .A2(_0462_),
    .B1(_0463_),
    .B2(_0267_),
    .ZN(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3213_ (.A1(_0264_),
    .A2(_0263_),
    .Z(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3214_ (.A1(_0464_),
    .A2(_0465_),
    .Z(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3215_ (.A1(_0252_),
    .A2(_0453_),
    .Z(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3216_ (.A1(_0464_),
    .A2(_0465_),
    .Z(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3217_ (.A1(_0466_),
    .A2(_0467_),
    .B(_0468_),
    .ZN(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _3218_ (.A1(_0265_),
    .A2(_0270_),
    .A3(_0273_),
    .ZN(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3219_ (.A1(_0469_),
    .A2(_0471_),
    .ZN(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3220_ (.A1(_0469_),
    .A2(_0471_),
    .ZN(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3221_ (.A1(_0460_),
    .A2(_0472_),
    .B(_0473_),
    .ZN(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3222_ (.A1(_0287_),
    .A2(_0288_),
    .ZN(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3223_ (.A1(_0474_),
    .A2(_0475_),
    .Z(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3224_ (.A1(_1444_),
    .A2(_0256_),
    .B1(_0455_),
    .B2(_0458_),
    .ZN(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3225_ (.A1(_0474_),
    .A2(_0475_),
    .ZN(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3226_ (.A1(_0476_),
    .A2(_0477_),
    .B(_0478_),
    .ZN(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3227_ (.A1(_0259_),
    .A2(_0319_),
    .ZN(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3228_ (.A1(_0479_),
    .A2(_0480_),
    .ZN(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3229_ (.A1(_0321_),
    .A2(_0358_),
    .B(_0482_),
    .ZN(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3230_ (.A1(_0398_),
    .A2(_0392_),
    .A3(_0397_),
    .Z(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3231_ (.A1(_0483_),
    .A2(_0484_),
    .ZN(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3232_ (.A1(_1415_),
    .A2(_0351_),
    .ZN(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3233_ (.A1(_0306_),
    .A2(_0452_),
    .B(_0486_),
    .ZN(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3234_ (.A1(_0241_),
    .A2(_0487_),
    .Z(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3235_ (.I(_0461_),
    .Z(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3236_ (.I(_0278_),
    .Z(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3237_ (.I(_0490_),
    .Z(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3238_ (.A1(_0282_),
    .A2(_0461_),
    .ZN(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3239_ (.I0(_0461_),
    .I1(_0493_),
    .S(_0490_),
    .Z(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3240_ (.A1(_0262_),
    .A2(_0494_),
    .ZN(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3241_ (.A1(_0489_),
    .A2(_0491_),
    .B(_0495_),
    .ZN(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3242_ (.A1(_0336_),
    .A2(_0260_),
    .B(_0463_),
    .ZN(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3243_ (.A1(_0054_),
    .A2(_0497_),
    .Z(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3244_ (.A1(_0496_),
    .A2(_0498_),
    .ZN(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3245_ (.A1(_0496_),
    .A2(_0498_),
    .ZN(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3246_ (.A1(_0488_),
    .A2(_0499_),
    .B(_0500_),
    .ZN(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3247_ (.A1(_0466_),
    .A2(_0467_),
    .Z(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3248_ (.A1(_0501_),
    .A2(_0502_),
    .ZN(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3249_ (.A1(_0251_),
    .A2(_0487_),
    .B(_0486_),
    .ZN(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3250_ (.A1(_0501_),
    .A2(_0502_),
    .ZN(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3251_ (.A1(_0505_),
    .A2(_0506_),
    .Z(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _3252_ (.A1(_0469_),
    .A2(_0471_),
    .A3(_0460_),
    .ZN(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3253_ (.A1(_0504_),
    .A2(_0507_),
    .B(_0508_),
    .ZN(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3254_ (.A1(_0321_),
    .A2(_0358_),
    .ZN(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3255_ (.A1(_0479_),
    .A2(_0480_),
    .Z(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3256_ (.A1(_0476_),
    .A2(_0477_),
    .ZN(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _3257_ (.A1(_0482_),
    .A2(_0510_),
    .A3(_0511_),
    .A4(_0512_),
    .ZN(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3258_ (.A1(_0509_),
    .A2(_0513_),
    .Z(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3259_ (.A1(_0483_),
    .A2(_0484_),
    .ZN(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3260_ (.A1(_0485_),
    .A2(_0515_),
    .B(_0516_),
    .ZN(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3261_ (.I(_0185_),
    .Z(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3262_ (.A1(_0268_),
    .A2(_0490_),
    .ZN(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3263_ (.A1(_0518_),
    .A2(_0490_),
    .B(_0519_),
    .ZN(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3264_ (.A1(_0518_),
    .A2(_0491_),
    .B1(_0520_),
    .B2(_0462_),
    .ZN(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3265_ (.A1(_0262_),
    .A2(_0494_),
    .Z(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3266_ (.A1(_0521_),
    .A2(_0522_),
    .ZN(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3267_ (.I(_1415_),
    .ZN(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3268_ (.I(_0285_),
    .Z(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3269_ (.A1(_0526_),
    .A2(_0304_),
    .ZN(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3270_ (.A1(_0524_),
    .A2(_0526_),
    .B(_0527_),
    .ZN(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3271_ (.A1(_0243_),
    .A2(_0528_),
    .Z(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3272_ (.A1(_0521_),
    .A2(_0522_),
    .ZN(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3273_ (.A1(_0529_),
    .A2(_0530_),
    .Z(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3274_ (.A1(_0496_),
    .A2(_0498_),
    .A3(_0488_),
    .Z(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3275_ (.A1(_0523_),
    .A2(_0531_),
    .B(_0532_),
    .ZN(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3276_ (.A1(_0524_),
    .A2(_0526_),
    .B1(_0528_),
    .B2(_0451_),
    .ZN(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3277_ (.A1(_0523_),
    .A2(_0531_),
    .ZN(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3278_ (.A1(_0532_),
    .A2(_0535_),
    .Z(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3279_ (.A1(_0534_),
    .A2(_0537_),
    .ZN(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3280_ (.A1(_0505_),
    .A2(_0506_),
    .Z(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3281_ (.A1(_0533_),
    .A2(_0538_),
    .A3(_0539_),
    .ZN(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3282_ (.A1(_0529_),
    .A2(_0530_),
    .Z(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3283_ (.I(_0245_),
    .Z(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3284_ (.A1(_1429_),
    .A2(_0249_),
    .Z(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3285_ (.A1(_0245_),
    .A2(_0543_),
    .ZN(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3286_ (.A1(_1429_),
    .A2(_0542_),
    .B(_0544_),
    .ZN(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3287_ (.A1(_0452_),
    .A2(_0545_),
    .ZN(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3288_ (.A1(_0336_),
    .A2(_0276_),
    .B(_0266_),
    .ZN(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3289_ (.A1(_0489_),
    .A2(_0268_),
    .B1(_0542_),
    .B2(_0548_),
    .ZN(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3290_ (.A1(_0462_),
    .A2(_0520_),
    .Z(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3291_ (.A1(_0549_),
    .A2(_0550_),
    .ZN(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3292_ (.A1(_0549_),
    .A2(_0550_),
    .ZN(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3293_ (.A1(_0546_),
    .A2(_0551_),
    .B(_0552_),
    .ZN(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3294_ (.A1(_0541_),
    .A2(_0553_),
    .Z(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3295_ (.A1(_0534_),
    .A2(_0537_),
    .Z(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3296_ (.A1(_0452_),
    .A2(_0545_),
    .ZN(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3297_ (.A1(_0244_),
    .A2(_0526_),
    .B(_0556_),
    .ZN(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3298_ (.A1(_0541_),
    .A2(_0553_),
    .ZN(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3299_ (.A1(_0557_),
    .A2(_0559_),
    .ZN(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3300_ (.A1(_0491_),
    .A2(_0543_),
    .ZN(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3301_ (.A1(_0268_),
    .A2(_0542_),
    .A3(_0561_),
    .ZN(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3302_ (.A1(_0276_),
    .A2(_0493_),
    .B(_0548_),
    .ZN(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3303_ (.A1(_0542_),
    .A2(_0563_),
    .ZN(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3304_ (.A1(_0561_),
    .A2(_0564_),
    .ZN(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3305_ (.A1(_0306_),
    .A2(_0565_),
    .ZN(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3306_ (.A1(_0306_),
    .A2(_0565_),
    .ZN(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3307_ (.A1(_0491_),
    .A2(_0543_),
    .B(_0567_),
    .ZN(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3308_ (.A1(_0562_),
    .A2(_0566_),
    .A3(_0568_),
    .Z(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3309_ (.A1(_0546_),
    .A2(_0551_),
    .Z(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3310_ (.A1(_0557_),
    .A2(_0559_),
    .ZN(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3311_ (.A1(_0570_),
    .A2(_0571_),
    .B(_0572_),
    .ZN(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3312_ (.A1(_0560_),
    .A2(_0573_),
    .ZN(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3313_ (.A1(_0561_),
    .A2(_0564_),
    .B1(_0570_),
    .B2(_0571_),
    .C(_0567_),
    .ZN(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3314_ (.A1(_0554_),
    .A2(_0555_),
    .B(_0575_),
    .ZN(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3315_ (.A1(_0554_),
    .A2(_0555_),
    .B(_0574_),
    .C(_0576_),
    .ZN(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3316_ (.A1(_0533_),
    .A2(_0538_),
    .B(_0539_),
    .ZN(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _3317_ (.A1(_0554_),
    .A2(_0560_),
    .B1(_0539_),
    .B2(_0533_),
    .C(_0555_),
    .ZN(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3318_ (.A1(_0578_),
    .A2(_0579_),
    .Z(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3319_ (.A1(_0540_),
    .A2(_0577_),
    .B(_0581_),
    .ZN(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3320_ (.A1(_0504_),
    .A2(_0507_),
    .ZN(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3321_ (.A1(_0508_),
    .A2(_0583_),
    .ZN(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3322_ (.A1(_0485_),
    .A2(_0513_),
    .A3(_0582_),
    .A4(_0584_),
    .ZN(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3323_ (.A1(_0517_),
    .A2(_0585_),
    .Z(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _3324_ (.A1(_0444_),
    .A2(_0446_),
    .B1(_0450_),
    .B2(_0586_),
    .ZN(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3325_ (.A1(_0224_),
    .A2(_0225_),
    .Z(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3326_ (.A1(_0160_),
    .A2(_0588_),
    .Z(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _3327_ (.A1(_1399_),
    .A2(_0402_),
    .ZN(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3328_ (.A1(_0439_),
    .A2(_0440_),
    .Z(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3329_ (.A1(_0436_),
    .A2(_0441_),
    .B(_0592_),
    .ZN(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3330_ (.A1(_0196_),
    .A2(_0222_),
    .Z(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _3331_ (.A1(_0593_),
    .A2(_0594_),
    .Z(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3332_ (.A1(_0593_),
    .A2(_0594_),
    .ZN(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _3333_ (.A1(_0590_),
    .A2(_0595_),
    .B(_0596_),
    .ZN(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3334_ (.A1(_0589_),
    .A2(_0597_),
    .Z(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _3335_ (.A1(_0590_),
    .A2(_0595_),
    .ZN(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3336_ (.A1(_0433_),
    .A2(_0442_),
    .ZN(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3337_ (.A1(_0433_),
    .A2(_0442_),
    .ZN(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3338_ (.A1(_0431_),
    .A2(_0600_),
    .B(_0601_),
    .ZN(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3339_ (.A1(_0599_),
    .A2(_0603_),
    .Z(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3340_ (.A1(_0598_),
    .A2(_0604_),
    .Z(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3341_ (.A1(_1381_),
    .A2(_0402_),
    .ZN(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3342_ (.A1(_0606_),
    .A2(_0588_),
    .Z(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3343_ (.A1(_0606_),
    .A2(_0588_),
    .ZN(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3344_ (.A1(_0224_),
    .A2(_0225_),
    .A3(_0606_),
    .Z(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _3345_ (.A1(_0590_),
    .A2(_0595_),
    .B(_0609_),
    .C(_0596_),
    .ZN(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__oai33_4 _3346_ (.A1(_0607_),
    .A2(_0608_),
    .A3(_0597_),
    .B1(_0610_),
    .B2(_0599_),
    .B3(_0603_),
    .ZN(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _3347_ (.A1(_0587_),
    .A2(_0605_),
    .B(_0611_),
    .C(_0238_),
    .ZN(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3348_ (.A1(_1897_),
    .A2(_0078_),
    .ZN(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3349_ (.A1(_0081_),
    .A2(_0614_),
    .B(_0080_),
    .ZN(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _3350_ (.A1(_0083_),
    .A2(_0240_),
    .A3(_0612_),
    .B(_0615_),
    .ZN(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3351_ (.A1(_1807_),
    .A2(_1832_),
    .B1(_1837_),
    .B2(_0616_),
    .ZN(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3352_ (.A1(_1811_),
    .A2(_1831_),
    .ZN(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3353_ (.A1(_1834_),
    .A2(_1832_),
    .B(_0618_),
    .ZN(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3354_ (.A1(_1186_),
    .A2(_1817_),
    .B1(_0395_),
    .B2(_1229_),
    .ZN(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3355_ (.A1(_1822_),
    .A2(_1826_),
    .Z(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3356_ (.A1(_1821_),
    .A2(_1827_),
    .B(_0621_),
    .ZN(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3357_ (.I(_1617_),
    .Z(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _3358_ (.A1(_1702_),
    .A2(_1863_),
    .B1(_1640_),
    .B2(_0623_),
    .C(_1503_),
    .ZN(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3359_ (.A1(_1823_),
    .A2(_1825_),
    .ZN(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3360_ (.A1(_1857_),
    .A2(_1655_),
    .ZN(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3361_ (.A1(_1586_),
    .A2(_1549_),
    .B(_1852_),
    .ZN(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3362_ (.A1(_0627_),
    .A2(_0628_),
    .Z(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3363_ (.A1(_0626_),
    .A2(_0629_),
    .Z(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3364_ (.A1(_0625_),
    .A2(_0630_),
    .ZN(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _3365_ (.A1(_0620_),
    .A2(_0622_),
    .A3(_0631_),
    .ZN(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3366_ (.A1(_1820_),
    .A2(_1828_),
    .ZN(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3367_ (.A1(_1818_),
    .A2(_1829_),
    .B(_0633_),
    .ZN(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3368_ (.A1(_0632_),
    .A2(_0634_),
    .Z(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3369_ (.A1(_0632_),
    .A2(_0634_),
    .ZN(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3370_ (.A1(_0636_),
    .A2(_0637_),
    .ZN(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3371_ (.A1(_1816_),
    .A2(_1830_),
    .Z(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3372_ (.A1(_1816_),
    .A2(_1830_),
    .Z(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3373_ (.A1(_1814_),
    .A2(_0639_),
    .B(_0640_),
    .ZN(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3374_ (.A1(_0638_),
    .A2(_0641_),
    .Z(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3375_ (.A1(_0619_),
    .A2(_0642_),
    .Z(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3376_ (.A1(_0617_),
    .A2(_0643_),
    .ZN(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3377_ (.A1(_1459_),
    .A2(_0644_),
    .ZN(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3378_ (.I(_1340_),
    .ZN(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3379_ (.A1(_1837_),
    .A2(_0616_),
    .Z(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _3380_ (.A1(_0079_),
    .A2(_0240_),
    .A3(_0612_),
    .B1(_0078_),
    .B2(_1897_),
    .ZN(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3381_ (.A1(_0082_),
    .A2(_0649_),
    .ZN(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3382_ (.I(\dsynth.freeRunCntr[6] ),
    .ZN(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3383_ (.A1(_0647_),
    .A2(_0648_),
    .B1(_0650_),
    .B2(_0651_),
    .ZN(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3384_ (.A1(_0240_),
    .A2(_0612_),
    .ZN(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3385_ (.A1(_0079_),
    .A2(_0653_),
    .ZN(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3386_ (.I(_1382_),
    .ZN(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3387_ (.A1(_0651_),
    .A2(_0650_),
    .B1(_0654_),
    .B2(_0655_),
    .ZN(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3388_ (.A1(_1836_),
    .A2(_0616_),
    .Z(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _3389_ (.A1(_1459_),
    .A2(_0644_),
    .B1(_0652_),
    .B2(_0656_),
    .C1(_0658_),
    .C2(_1461_),
    .ZN(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3390_ (.A1(_0645_),
    .A2(_0659_),
    .Z(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3391_ (.A1(_1314_),
    .A2(_0644_),
    .Z(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3392_ (.A1(_1459_),
    .A2(_0644_),
    .B1(_0658_),
    .B2(_1461_),
    .ZN(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3393_ (.A1(_0082_),
    .A2(_0649_),
    .Z(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3394_ (.A1(_1461_),
    .A2(_0658_),
    .B1(_0663_),
    .B2(_1451_),
    .ZN(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3395_ (.A1(_0655_),
    .A2(_0654_),
    .B(_0656_),
    .C(_0664_),
    .ZN(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3396_ (.A1(_0394_),
    .A2(_0400_),
    .Z(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3397_ (.A1(_0427_),
    .A2(_0424_),
    .Z(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3398_ (.A1(_0403_),
    .A2(_0424_),
    .B(_0445_),
    .ZN(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3399_ (.A1(_0666_),
    .A2(_0667_),
    .B1(_0669_),
    .B2(_0447_),
    .ZN(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3400_ (.A1(_0666_),
    .A2(_0667_),
    .B1(_0517_),
    .B2(_0585_),
    .C(_0446_),
    .ZN(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3401_ (.A1(_0670_),
    .A2(_0449_),
    .B(_0671_),
    .ZN(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3402_ (.A1(_0598_),
    .A2(_0604_),
    .ZN(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3403_ (.A1(_0589_),
    .A2(_0597_),
    .ZN(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3404_ (.A1(_0599_),
    .A2(_0603_),
    .ZN(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3405_ (.A1(_0674_),
    .A2(_0675_),
    .ZN(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3406_ (.A1(_0672_),
    .A2(_0673_),
    .B1(_0676_),
    .B2(_0610_),
    .ZN(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3407_ (.A1(_0158_),
    .A2(_0229_),
    .Z(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3408_ (.A1(_0231_),
    .A2(_0677_),
    .B(_0678_),
    .ZN(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3409_ (.A1(_0235_),
    .A2(_0680_),
    .Z(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3410_ (.A1(_0231_),
    .A2(_0677_),
    .ZN(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3411_ (.A1(_1385_),
    .A2(_0681_),
    .B1(_0682_),
    .B2(_1463_),
    .ZN(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3412_ (.I(_1419_),
    .Z(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3413_ (.I(_0684_),
    .ZN(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3414_ (.A1(_0587_),
    .A2(_0604_),
    .B(_0675_),
    .ZN(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3415_ (.A1(_0598_),
    .A2(_0686_),
    .ZN(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3416_ (.A1(_0685_),
    .A2(_0687_),
    .ZN(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3417_ (.A1(_0672_),
    .A2(_0604_),
    .Z(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3418_ (.A1(_1465_),
    .A2(_0689_),
    .ZN(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3419_ (.A1(_0685_),
    .A2(_0687_),
    .B(_0691_),
    .ZN(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3420_ (.A1(_1464_),
    .A2(_0682_),
    .B1(_0688_),
    .B2(_0692_),
    .ZN(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3421_ (.A1(_1385_),
    .A2(_0681_),
    .ZN(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3422_ (.A1(_0683_),
    .A2(_0693_),
    .B(_0694_),
    .ZN(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _3423_ (.A1(_0661_),
    .A2(_0662_),
    .A3(_0665_),
    .A4(_0695_),
    .ZN(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3424_ (.I(\dsynth.freeRunCntr[12] ),
    .ZN(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3425_ (.I(_0697_),
    .Z(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3426_ (.I(_1857_),
    .Z(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _3427_ (.A1(_1596_),
    .A2(_1685_),
    .B1(_1824_),
    .B2(_0623_),
    .C1(_0699_),
    .C2(_1576_),
    .ZN(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3428_ (.I(_1584_),
    .Z(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3429_ (.A1(_0702_),
    .A2(_1549_),
    .B(_1597_),
    .ZN(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3430_ (.A1(_0699_),
    .A2(_1824_),
    .A3(_0703_),
    .ZN(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_4 _3431_ (.A1(_1132_),
    .A2(_0256_),
    .B1(_1700_),
    .B2(_0991_),
    .C1(_1095_),
    .C2(_1668_),
    .ZN(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _3432_ (.A1(_0700_),
    .A2(_0704_),
    .A3(_0705_),
    .ZN(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3433_ (.I(_1655_),
    .Z(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3434_ (.A1(_1617_),
    .A2(_0707_),
    .ZN(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _3435_ (.A1(_1128_),
    .A2(_0256_),
    .B(_0708_),
    .C(_1498_),
    .ZN(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3436_ (.A1(_1857_),
    .A2(_0707_),
    .A3(_0628_),
    .ZN(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3437_ (.A1(_1765_),
    .A2(_1824_),
    .ZN(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3438_ (.A1(_0711_),
    .A2(_0703_),
    .Z(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3439_ (.A1(_0710_),
    .A2(_0713_),
    .Z(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3440_ (.A1(_0710_),
    .A2(_0713_),
    .ZN(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3441_ (.A1(_0709_),
    .A2(_0714_),
    .B(_0715_),
    .ZN(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3442_ (.A1(_0706_),
    .A2(_0716_),
    .Z(_0717_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _3443_ (.A1(_1823_),
    .A2(_1825_),
    .A3(_0629_),
    .B1(_0630_),
    .B2(_0625_),
    .ZN(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3444_ (.A1(_0709_),
    .A2(_0714_),
    .Z(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3445_ (.A1(_0718_),
    .A2(_0719_),
    .ZN(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3446_ (.A1(_0991_),
    .A2(_1817_),
    .B1(_0395_),
    .B2(_1186_),
    .ZN(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3447_ (.A1(_0718_),
    .A2(_0719_),
    .Z(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3448_ (.A1(_0721_),
    .A2(_0722_),
    .ZN(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3449_ (.A1(_0720_),
    .A2(_0724_),
    .ZN(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3450_ (.A1(_0717_),
    .A2(_0725_),
    .ZN(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3451_ (.A1(_0706_),
    .A2(_0716_),
    .Z(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3452_ (.A1(_1702_),
    .A2(_0159_),
    .ZN(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3453_ (.A1(_1128_),
    .A2(_1668_),
    .ZN(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3454_ (.A1(_1576_),
    .A2(_0623_),
    .B1(_0699_),
    .B2(_1634_),
    .ZN(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3455_ (.A1(_0729_),
    .A2(_0730_),
    .Z(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3456_ (.A1(_0728_),
    .A2(_0731_),
    .ZN(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3457_ (.A1(_0700_),
    .A2(_0704_),
    .ZN(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3458_ (.A1(_0700_),
    .A2(_0704_),
    .ZN(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3459_ (.A1(_0733_),
    .A2(_0705_),
    .B(_0735_),
    .ZN(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3460_ (.A1(_0732_),
    .A2(_0736_),
    .Z(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3461_ (.A1(_0727_),
    .A2(_0737_),
    .Z(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3462_ (.A1(_0726_),
    .A2(_0738_),
    .Z(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3463_ (.A1(_0717_),
    .A2(_0725_),
    .Z(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3464_ (.A1(_0721_),
    .A2(_0722_),
    .ZN(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3465_ (.A1(_0622_),
    .A2(_0631_),
    .ZN(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3466_ (.A1(_0622_),
    .A2(_0631_),
    .ZN(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3467_ (.A1(_0620_),
    .A2(_0742_),
    .B(_0743_),
    .ZN(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3468_ (.A1(_0741_),
    .A2(_0744_),
    .ZN(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3469_ (.A1(_0740_),
    .A2(_0746_),
    .Z(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3470_ (.A1(_0741_),
    .A2(_0744_),
    .ZN(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3471_ (.A1(_0636_),
    .A2(_0748_),
    .ZN(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3472_ (.A1(_0747_),
    .A2(_0749_),
    .Z(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3473_ (.A1(_0739_),
    .A2(_0750_),
    .ZN(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3474_ (.A1(_0230_),
    .A2(_0235_),
    .A3(_0611_),
    .Z(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3475_ (.A1(_1836_),
    .A2(_0643_),
    .Z(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3476_ (.A1(_0083_),
    .A2(_0753_),
    .ZN(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3477_ (.A1(_0238_),
    .A2(_0752_),
    .B(_0754_),
    .ZN(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3478_ (.A1(_1834_),
    .A2(_1832_),
    .A3(_0642_),
    .Z(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3479_ (.A1(_1807_),
    .A2(_1835_),
    .ZN(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3480_ (.A1(_0758_),
    .A2(_0643_),
    .ZN(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3481_ (.A1(_0615_),
    .A2(_0753_),
    .ZN(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3482_ (.A1(_0757_),
    .A2(_0759_),
    .A3(_0760_),
    .ZN(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3483_ (.A1(_0638_),
    .A2(_0641_),
    .ZN(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3484_ (.A1(_0636_),
    .A2(_0748_),
    .Z(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3485_ (.A1(_0762_),
    .A2(_0763_),
    .Z(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3486_ (.A1(_0749_),
    .A2(_0764_),
    .ZN(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3487_ (.A1(_0747_),
    .A2(_0765_),
    .ZN(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3488_ (.A1(_0618_),
    .A2(_0642_),
    .B(_0762_),
    .ZN(_0768_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3489_ (.A1(_0763_),
    .A2(_0768_),
    .ZN(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3490_ (.A1(_0766_),
    .A2(_0769_),
    .ZN(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3491_ (.A1(_0755_),
    .A2(_0761_),
    .B(_0770_),
    .ZN(_0771_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3492_ (.A1(_0618_),
    .A2(_0642_),
    .A3(_0763_),
    .Z(_0772_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3493_ (.A1(_0747_),
    .A2(_0764_),
    .B1(_0766_),
    .B2(_0772_),
    .ZN(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3494_ (.I(_0773_),
    .ZN(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3495_ (.A1(_0740_),
    .A2(_0746_),
    .Z(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3496_ (.A1(_0775_),
    .A2(_0750_),
    .ZN(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3497_ (.A1(_0739_),
    .A2(_0776_),
    .Z(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3498_ (.I(_0777_),
    .Z(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3499_ (.I(_0779_),
    .ZN(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3500_ (.A1(_0771_),
    .A2(_0774_),
    .B(_0780_),
    .ZN(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3501_ (.A1(_1129_),
    .A2(_0395_),
    .ZN(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3502_ (.A1(_1129_),
    .A2(_1817_),
    .A3(_0730_),
    .ZN(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3503_ (.A1(_0129_),
    .A2(_1902_),
    .ZN(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3504_ (.A1(_1634_),
    .A2(_0623_),
    .B1(_0699_),
    .B2(_1596_),
    .ZN(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3505_ (.A1(_0784_),
    .A2(_0785_),
    .Z(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3506_ (.A1(_0783_),
    .A2(_0786_),
    .Z(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _3507_ (.A1(_0782_),
    .A2(_0787_),
    .Z(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3508_ (.A1(_0728_),
    .A2(_0731_),
    .ZN(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3509_ (.A1(_0732_),
    .A2(_0736_),
    .ZN(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3510_ (.A1(_0790_),
    .A2(_0791_),
    .ZN(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3511_ (.A1(_0788_),
    .A2(_0792_),
    .Z(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3512_ (.I(_0727_),
    .ZN(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3513_ (.A1(_0794_),
    .A2(_0737_),
    .ZN(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3514_ (.A1(_0726_),
    .A2(_0738_),
    .Z(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3515_ (.A1(_0795_),
    .A2(_0796_),
    .ZN(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3516_ (.A1(_0793_),
    .A2(_0797_),
    .Z(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3517_ (.I(_0798_),
    .Z(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3518_ (.A1(_0739_),
    .A2(_0775_),
    .ZN(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3519_ (.A1(_0799_),
    .A2(_0801_),
    .Z(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3520_ (.I(_0802_),
    .ZN(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3521_ (.A1(_0798_),
    .A2(_0801_),
    .Z(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3522_ (.A1(_0803_),
    .A2(_0804_),
    .ZN(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3523_ (.A1(_0751_),
    .A2(_0781_),
    .B(_0805_),
    .ZN(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3524_ (.I(_0751_),
    .ZN(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3525_ (.I(_0805_),
    .ZN(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3526_ (.A1(_0236_),
    .A2(_0237_),
    .Z(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3527_ (.A1(_0231_),
    .A2(_0235_),
    .A3(_0611_),
    .ZN(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _3528_ (.A1(_0809_),
    .A2(_0810_),
    .B(_0753_),
    .C(_0083_),
    .ZN(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _3529_ (.A1(_0757_),
    .A2(_0759_),
    .A3(_0760_),
    .Z(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3530_ (.I(_0766_),
    .Z(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3531_ (.A1(_0812_),
    .A2(_0813_),
    .B(_0814_),
    .C(_0769_),
    .ZN(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3532_ (.A1(_0815_),
    .A2(_0773_),
    .B(_0779_),
    .ZN(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3533_ (.A1(_0807_),
    .A2(_0808_),
    .A3(_0816_),
    .ZN(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3534_ (.A1(_0698_),
    .A2(_0806_),
    .A3(_0817_),
    .ZN(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _3535_ (.A1(_0799_),
    .A2(_0777_),
    .A3(_0770_),
    .Z(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3536_ (.A1(_0755_),
    .A2(_0761_),
    .B(_0819_),
    .ZN(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _3537_ (.A1(_0799_),
    .A2(_0777_),
    .A3(_0773_),
    .Z(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3538_ (.A1(_0804_),
    .A2(_0751_),
    .Z(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3539_ (.A1(_0821_),
    .A2(_0802_),
    .A3(_0823_),
    .ZN(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3540_ (.A1(_0793_),
    .A2(_0796_),
    .Z(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3541_ (.A1(_0793_),
    .A2(_0795_),
    .ZN(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3542_ (.A1(_0788_),
    .A2(_0790_),
    .ZN(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3543_ (.A1(_0783_),
    .A2(_0786_),
    .ZN(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3544_ (.A1(_0782_),
    .A2(_0787_),
    .ZN(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3545_ (.A1(_0828_),
    .A2(_0829_),
    .ZN(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3546_ (.A1(_0784_),
    .A2(_0785_),
    .ZN(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3547_ (.A1(_1681_),
    .A2(_1515_),
    .ZN(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3548_ (.A1(_1132_),
    .A2(_0396_),
    .ZN(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3549_ (.A1(_0832_),
    .A2(_0834_),
    .Z(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3550_ (.A1(_0831_),
    .A2(_0835_),
    .ZN(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3551_ (.A1(_0830_),
    .A2(_0836_),
    .Z(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3552_ (.A1(_0827_),
    .A2(_0837_),
    .Z(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _3553_ (.A1(_0788_),
    .A2(_0791_),
    .B(_0826_),
    .C(_0838_),
    .ZN(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3554_ (.A1(_0825_),
    .A2(_0839_),
    .Z(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3555_ (.A1(_0820_),
    .A2(_0824_),
    .B(_0840_),
    .ZN(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3556_ (.A1(_0799_),
    .A2(_0779_),
    .A3(_0770_),
    .ZN(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3557_ (.A1(_0812_),
    .A2(_0813_),
    .B(_0842_),
    .ZN(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3558_ (.A1(_0821_),
    .A2(_0802_),
    .A3(_0823_),
    .Z(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3559_ (.I(_0840_),
    .ZN(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3560_ (.A1(_0843_),
    .A2(_0845_),
    .A3(_0846_),
    .ZN(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3561_ (.A1(_0841_),
    .A2(_0847_),
    .B(_1136_),
    .ZN(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3562_ (.I(\dsynth.freeRunCntr[14] ),
    .ZN(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3563_ (.A1(_0843_),
    .A2(_0845_),
    .B(_0846_),
    .ZN(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3564_ (.A1(_0828_),
    .A2(_0829_),
    .B(_0836_),
    .ZN(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3565_ (.A1(_0832_),
    .A2(_0834_),
    .B(_0851_),
    .ZN(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _3566_ (.A1(_0827_),
    .A2(_0837_),
    .B1(_0839_),
    .B2(_0825_),
    .C(_0852_),
    .ZN(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3567_ (.A1(\dsynth.freeRunCntr[16] ),
    .A2(_1118_),
    .ZN(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _3568_ (.A1(_0849_),
    .A2(_0850_),
    .A3(_0853_),
    .B(_0854_),
    .ZN(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3569_ (.A1(_1136_),
    .A2(_0841_),
    .A3(_0847_),
    .Z(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3570_ (.I(_0853_),
    .ZN(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3571_ (.A1(_0841_),
    .A2(_0858_),
    .B(_1103_),
    .ZN(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _3572_ (.A1(_0848_),
    .A2(_0856_),
    .A3(_0857_),
    .A4(_0859_),
    .Z(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3573_ (.A1(_0807_),
    .A2(_0805_),
    .A3(_0816_),
    .ZN(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3574_ (.A1(_0751_),
    .A2(_0781_),
    .B(_0808_),
    .ZN(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3575_ (.A1(_0779_),
    .A2(_0771_),
    .A3(_0774_),
    .ZN(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3576_ (.A1(_0815_),
    .A2(_0773_),
    .B(_0780_),
    .ZN(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3577_ (.A1(_0863_),
    .A2(_0864_),
    .ZN(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _3578_ (.A1(\dsynth.freeRunCntr[12] ),
    .A2(_0861_),
    .A3(_0862_),
    .B1(_0865_),
    .B2(_1232_),
    .ZN(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3579_ (.I(_1230_),
    .ZN(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3580_ (.I(_0772_),
    .ZN(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3581_ (.A1(_0812_),
    .A2(_0813_),
    .B(_0769_),
    .ZN(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3582_ (.A1(_0814_),
    .A2(_0869_),
    .A3(_0870_),
    .Z(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3583_ (.A1(_0869_),
    .A2(_0870_),
    .B(_0814_),
    .ZN(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3584_ (.I(\dsynth.freeRunCntr[10] ),
    .ZN(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__oai33_1 _3585_ (.A1(_0868_),
    .A2(_0863_),
    .A3(_0864_),
    .B1(_0871_),
    .B2(_0872_),
    .B3(_0873_),
    .ZN(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3586_ (.I(_0814_),
    .ZN(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3587_ (.A1(_0875_),
    .A2(_0869_),
    .A3(_0870_),
    .Z(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3588_ (.A1(_0869_),
    .A2(_0870_),
    .B(_0875_),
    .ZN(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3589_ (.A1(\dsynth.freeRunCntr[10] ),
    .A2(_0876_),
    .A3(_0878_),
    .ZN(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3590_ (.A1(_0755_),
    .A2(_0761_),
    .ZN(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3591_ (.A1(_0880_),
    .A2(_0769_),
    .ZN(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3592_ (.A1(_1288_),
    .A2(_0881_),
    .ZN(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3593_ (.A1(_1288_),
    .A2(_0881_),
    .Z(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _3594_ (.A1(_0874_),
    .A2(_0879_),
    .A3(_0882_),
    .A4(_0883_),
    .Z(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _3595_ (.A1(_0818_),
    .A2(_0860_),
    .A3(_0867_),
    .A4(_0884_),
    .ZN(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3596_ (.A1(_0660_),
    .A2(_0696_),
    .B(_0885_),
    .ZN(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3597_ (.A1(_0818_),
    .A2(_0860_),
    .ZN(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3598_ (.A1(_0879_),
    .A2(_0882_),
    .ZN(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3599_ (.A1(_0806_),
    .A2(_0817_),
    .B(_0698_),
    .ZN(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _3600_ (.A1(_1232_),
    .A2(_0865_),
    .B1(_0874_),
    .B2(_0889_),
    .C(_0890_),
    .ZN(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3601_ (.A1(_0857_),
    .A2(_0859_),
    .ZN(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3602_ (.A1(_0856_),
    .A2(_0892_),
    .ZN(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3603_ (.A1(_0887_),
    .A2(_0891_),
    .B(_0893_),
    .ZN(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _3604_ (.A1(_0661_),
    .A2(_0662_),
    .A3(_0665_),
    .Z(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3605_ (.A1(_1465_),
    .A2(_0689_),
    .B(_0694_),
    .ZN(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3606_ (.A1(_0685_),
    .A2(_0687_),
    .B(_0692_),
    .ZN(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3607_ (.A1(_1464_),
    .A2(_0682_),
    .ZN(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3608_ (.A1(_0897_),
    .A2(_0898_),
    .ZN(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _3609_ (.A1(_0895_),
    .A2(_0683_),
    .A3(_0896_),
    .A4(_0900_),
    .ZN(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3610_ (.A1(_0886_),
    .A2(_0894_),
    .B1(_0901_),
    .B2(_0885_),
    .ZN(net25));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3611_ (.A1(_1463_),
    .A2(_0489_),
    .ZN(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3612_ (.A1(_0684_),
    .A2(_0295_),
    .B1(_0518_),
    .B2(_1445_),
    .ZN(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3613_ (.A1(_0684_),
    .A2(_0295_),
    .B(_0903_),
    .ZN(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3614_ (.I(\dsynth.freeRunCntr[4] ),
    .ZN(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3615_ (.A1(_0905_),
    .A2(_1848_),
    .ZN(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3616_ (.A1(_1385_),
    .A2(_0045_),
    .ZN(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3617_ (.A1(_1465_),
    .A2(_0518_),
    .Z(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3618_ (.A1(_0651_),
    .A2(_1728_),
    .B1(_1858_),
    .B2(_0655_),
    .ZN(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3619_ (.A1(_1382_),
    .A2(_0131_),
    .ZN(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3620_ (.A1(_1451_),
    .A2(_0033_),
    .ZN(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3621_ (.A1(_0910_),
    .A2(_0911_),
    .A3(_0912_),
    .Z(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3622_ (.A1(_0906_),
    .A2(_0907_),
    .A3(_0908_),
    .A4(_0913_),
    .ZN(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3623_ (.A1(_1131_),
    .A2(_1681_),
    .ZN(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3624_ (.A1(_1103_),
    .A2(_1586_),
    .B1(_1730_),
    .B2(\dsynth.freeRunCntr[13] ),
    .ZN(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3625_ (.A1(\dsynth.freeRunCntr[14] ),
    .A2(_1586_),
    .B1(_0702_),
    .B2(_1118_),
    .ZN(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3626_ (.A1(_1118_),
    .A2(_0702_),
    .ZN(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3627_ (.A1(_0063_),
    .A2(_1596_),
    .B1(_1730_),
    .B2(\dsynth.freeRunCntr[13] ),
    .C(_0918_),
    .ZN(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3628_ (.A1(_0917_),
    .A2(_0919_),
    .ZN(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3629_ (.A1(_0916_),
    .A2(_0921_),
    .ZN(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3630_ (.A1(_0698_),
    .A2(_0707_),
    .B(_0915_),
    .C(_0922_),
    .ZN(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3631_ (.I(_0923_),
    .ZN(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3632_ (.A1(_1463_),
    .A2(_0489_),
    .ZN(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3633_ (.A1(_0924_),
    .A2(_0925_),
    .ZN(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _3634_ (.A1(_0902_),
    .A2(_0904_),
    .A3(_0914_),
    .A4(_0926_),
    .ZN(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3635_ (.A1(\dsynth.freeRunCntr[7] ),
    .A2(_1528_),
    .B1(_1544_),
    .B2(_1313_),
    .ZN(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3636_ (.I(_0928_),
    .ZN(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3637_ (.A1(_1314_),
    .A2(_1544_),
    .ZN(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3638_ (.A1(_0647_),
    .A2(_1714_),
    .B(_0929_),
    .C(_0930_),
    .ZN(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3639_ (.A1(_0868_),
    .A2(_1640_),
    .B1(_0707_),
    .B2(_0698_),
    .ZN(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3640_ (.A1(_1233_),
    .A2(_1683_),
    .B1(_0048_),
    .B2(_1230_),
    .ZN(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3641_ (.A1(_1233_),
    .A2(_1683_),
    .B1(_1678_),
    .B2(_1288_),
    .ZN(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3642_ (.A1(_1290_),
    .A2(_1678_),
    .B(_0935_),
    .ZN(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3643_ (.A1(_0933_),
    .A2(_0934_),
    .A3(_0936_),
    .ZN(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3644_ (.A1(_0932_),
    .A2(_0937_),
    .ZN(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3645_ (.A1(_0916_),
    .A2(_0917_),
    .ZN(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _3646_ (.A1(_1123_),
    .A2(_0702_),
    .B1(_1681_),
    .B2(_1131_),
    .C(_0939_),
    .ZN(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3647_ (.A1(_0684_),
    .A2(_0295_),
    .ZN(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _3648_ (.A1(_0902_),
    .A2(_0941_),
    .A3(_0903_),
    .B(_0925_),
    .ZN(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3649_ (.A1(_0906_),
    .A2(_0943_),
    .ZN(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3650_ (.A1(_0944_),
    .A2(_0911_),
    .A3(_0907_),
    .ZN(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3651_ (.A1(_0910_),
    .A2(_0945_),
    .B(_0932_),
    .ZN(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3652_ (.A1(_0928_),
    .A2(_0930_),
    .B1(_0912_),
    .B2(_0946_),
    .ZN(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3653_ (.A1(_0935_),
    .A2(_0934_),
    .ZN(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3654_ (.A1(_0947_),
    .A2(_0937_),
    .B(_0933_),
    .C(_0948_),
    .ZN(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3655_ (.A1(_0915_),
    .A2(_0940_),
    .B1(_0924_),
    .B2(_0949_),
    .ZN(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3656_ (.A1(_0927_),
    .A2(_0938_),
    .B(_0950_),
    .ZN(net26));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3657_ (.I(net11),
    .Z(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3658_ (.I(net14),
    .ZN(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3659_ (.A1(_0951_),
    .A2(_0953_),
    .A3(net15),
    .ZN(net28));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3660_ (.I(net11),
    .ZN(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3661_ (.A1(_0954_),
    .A2(_0953_),
    .A3(net15),
    .ZN(net29));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3662_ (.A1(_0954_),
    .A2(net14),
    .A3(net15),
    .ZN(net16));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3663_ (.A1(_0951_),
    .A2(net14),
    .A3(net15),
    .ZN(net30));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3664_ (.I(net2),
    .Z(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3665_ (.A1(net3),
    .A2(net4),
    .B(net1),
    .ZN(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3666_ (.A1(_0955_),
    .A2(_0956_),
    .B(_0951_),
    .ZN(net20));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3667_ (.A1(net3),
    .A2(net4),
    .B(net1),
    .ZN(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3668_ (.A1(_0951_),
    .A2(_0955_),
    .A3(_0957_),
    .ZN(net19));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3669_ (.A1(_0954_),
    .A2(net1),
    .Z(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3670_ (.A1(net3),
    .A2(net4),
    .B(net2),
    .ZN(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3671_ (.A1(_0959_),
    .A2(_0960_),
    .ZN(net18));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3672_ (.A1(net3),
    .A2(net4),
    .B(net11),
    .C(net2),
    .ZN(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3673_ (.A1(_0959_),
    .A2(_0961_),
    .ZN(net17));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3674_ (.A1(_0955_),
    .A2(_0959_),
    .ZN(net22));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3675_ (.A1(net11),
    .A2(_0955_),
    .A3(net1),
    .ZN(net21));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3676_ (.A1(net43),
    .A2(\tmux.clkpab ),
    .B1(net5),
    .B2(\tmux.clkpbb ),
    .ZN(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3677_ (.I(_0962_),
    .ZN(net23));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3678_ (.I(net6),
    .ZN(_0964_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3679_ (.A1(\tmux.clkpab ),
    .A2(_0964_),
    .ZN(\tmux.clkbpb ));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3680_ (.A1(\tmux.clkpbb ),
    .A2(net6),
    .ZN(\tmux.clkapa ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3681_ (.A1(net43),
    .A2(\tgate.clkp ),
    .Z(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3682_ (.I(_0965_),
    .Z(net24));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3683_ (.I(net10),
    .Z(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3684_ (.I(_0966_),
    .ZN(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3685_ (.I(net7),
    .Z(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3686_ (.I(net9),
    .Z(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3687_ (.A1(net8),
    .A2(_0968_),
    .A3(_0969_),
    .ZN(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3688_ (.A1(_0967_),
    .A2(_0970_),
    .Z(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3689_ (.A1(\dsynth.freeRunCntr[0] ),
    .A2(_0972_),
    .ZN(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3690_ (.I(net7),
    .ZN(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _3691_ (.A1(net8),
    .A2(_0974_),
    .A3(net9),
    .A4(net10),
    .ZN(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3692_ (.A1(\dsynth.freeRunCntr[1] ),
    .A2(_0975_),
    .ZN(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3693_ (.A1(_0973_),
    .A2(_0976_),
    .Z(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3694_ (.I(_0977_),
    .Z(_0011_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3695_ (.I(net8),
    .Z(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3696_ (.I(_0974_),
    .Z(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3697_ (.A1(_0978_),
    .A2(_0979_),
    .ZN(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3698_ (.A1(_0969_),
    .A2(_0966_),
    .A3(_0980_),
    .ZN(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3699_ (.A1(\dsynth.freeRunCntr[2] ),
    .A2(_0982_),
    .Z(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3700_ (.A1(_1445_),
    .A2(_0975_),
    .ZN(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3701_ (.A1(_0973_),
    .A2(_0976_),
    .B(_0984_),
    .ZN(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3702_ (.A1(_0983_),
    .A2(_0985_),
    .Z(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3703_ (.I(_0986_),
    .Z(_0022_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3704_ (.I(_0969_),
    .Z(_0987_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3705_ (.A1(_0978_),
    .A2(_0968_),
    .ZN(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3706_ (.A1(_0987_),
    .A2(_0966_),
    .A3(_0988_),
    .ZN(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3707_ (.A1(_1419_),
    .A2(_0982_),
    .Z(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3708_ (.A1(_0983_),
    .A2(_0985_),
    .B(_0990_),
    .ZN(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _3709_ (.A1(_1464_),
    .A2(_0989_),
    .A3(_0992_),
    .ZN(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3710_ (.I(_0993_),
    .Z(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3711_ (.I(_0966_),
    .Z(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3712_ (.A1(_0978_),
    .A2(_0968_),
    .ZN(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3713_ (.A1(_0969_),
    .A2(_0995_),
    .ZN(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3714_ (.A1(_0994_),
    .A2(_0996_),
    .ZN(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3715_ (.A1(\dsynth.freeRunCntr[4] ),
    .A2(_0997_),
    .Z(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3716_ (.A1(\dsynth.freeRunCntr[3] ),
    .A2(_0989_),
    .ZN(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3717_ (.A1(_1417_),
    .A2(_0989_),
    .ZN(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3718_ (.A1(_0999_),
    .A2(_0992_),
    .B(_1000_),
    .ZN(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3719_ (.A1(_0998_),
    .A2(_1002_),
    .Z(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3720_ (.I(_1003_),
    .Z(_0027_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3721_ (.I(_0978_),
    .Z(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3722_ (.A1(_1004_),
    .A2(_0979_),
    .ZN(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3723_ (.A1(_0987_),
    .A2(_0967_),
    .A3(_1005_),
    .Z(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3724_ (.A1(_0905_),
    .A2(_0994_),
    .A3(_0996_),
    .ZN(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3725_ (.A1(_0998_),
    .A2(_1002_),
    .B(_1007_),
    .ZN(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3726_ (.A1(_0655_),
    .A2(_1006_),
    .A3(_1008_),
    .Z(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3727_ (.I(_1009_),
    .Z(_0028_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3728_ (.A1(_1004_),
    .A2(_0979_),
    .Z(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3729_ (.A1(_0987_),
    .A2(_1011_),
    .ZN(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3730_ (.A1(_0994_),
    .A2(_1012_),
    .ZN(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3731_ (.A1(\dsynth.freeRunCntr[6] ),
    .A2(_1013_),
    .Z(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3732_ (.A1(\dsynth.freeRunCntr[5] ),
    .A2(_1006_),
    .ZN(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3733_ (.A1(\dsynth.freeRunCntr[5] ),
    .A2(_1006_),
    .ZN(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3734_ (.A1(_1015_),
    .A2(_1008_),
    .B(_1016_),
    .ZN(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3735_ (.A1(_1014_),
    .A2(_1017_),
    .Z(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3736_ (.I(_1018_),
    .Z(_0029_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3737_ (.I(_0994_),
    .Z(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3738_ (.I(_0987_),
    .Z(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3739_ (.A1(_1004_),
    .A2(_0968_),
    .A3(_1021_),
    .ZN(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3740_ (.A1(_1019_),
    .A2(_1022_),
    .ZN(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3741_ (.A1(_0651_),
    .A2(_1019_),
    .A3(_1012_),
    .ZN(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3742_ (.A1(_1014_),
    .A2(_1017_),
    .B(_1024_),
    .ZN(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3743_ (.A1(_0647_),
    .A2(_1023_),
    .A3(_1025_),
    .Z(_1026_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3744_ (.I(_1026_),
    .Z(_0030_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3745_ (.I(_1019_),
    .Z(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3746_ (.A1(_1027_),
    .A2(_0970_),
    .B(_1313_),
    .ZN(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3747_ (.A1(\dsynth.freeRunCntr[8] ),
    .A2(_1019_),
    .A3(_0970_),
    .Z(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3748_ (.A1(_1028_),
    .A2(_1029_),
    .ZN(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3749_ (.A1(\dsynth.freeRunCntr[7] ),
    .A2(_1023_),
    .ZN(_1032_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3750_ (.A1(\dsynth.freeRunCntr[7] ),
    .A2(_1023_),
    .ZN(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3751_ (.A1(_1032_),
    .A2(_1025_),
    .B(_1033_),
    .ZN(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3752_ (.A1(_1031_),
    .A2(_1034_),
    .Z(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3753_ (.I(_1035_),
    .Z(_0031_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3754_ (.I(_1027_),
    .Z(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3755_ (.I(_1036_),
    .Z(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3756_ (.A1(_1004_),
    .A2(_0979_),
    .A3(_1021_),
    .ZN(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3757_ (.A1(_1037_),
    .A2(_1038_),
    .ZN(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3758_ (.A1(_1031_),
    .A2(_1034_),
    .B(_1029_),
    .ZN(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3759_ (.A1(_1290_),
    .A2(_1039_),
    .A3(_1041_),
    .Z(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3760_ (.I(_1042_),
    .Z(_0032_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _3761_ (.A1(_1021_),
    .A2(_0967_),
    .A3(_0980_),
    .Z(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3762_ (.A1(_0873_),
    .A2(_1043_),
    .Z(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3763_ (.A1(_1027_),
    .A2(_1038_),
    .B(\dsynth.freeRunCntr[9] ),
    .ZN(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3764_ (.A1(\dsynth.freeRunCntr[9] ),
    .A2(_1027_),
    .A3(_1038_),
    .ZN(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3765_ (.A1(_1045_),
    .A2(_1041_),
    .B(_1046_),
    .ZN(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3766_ (.A1(_1044_),
    .A2(_1047_),
    .Z(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3767_ (.I(_1048_),
    .Z(_0001_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3768_ (.I(_1021_),
    .Z(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3769_ (.A1(_1050_),
    .A2(_0988_),
    .ZN(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3770_ (.A1(_1037_),
    .A2(_1051_),
    .ZN(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3771_ (.A1(_0873_),
    .A2(_1043_),
    .ZN(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3772_ (.A1(_1044_),
    .A2(_1047_),
    .B(_1053_),
    .ZN(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3773_ (.A1(_1232_),
    .A2(_1052_),
    .A3(_1054_),
    .Z(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3774_ (.I(_1055_),
    .Z(_0002_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3775_ (.A1(_1050_),
    .A2(_1036_),
    .A3(_0995_),
    .ZN(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3776_ (.A1(_0697_),
    .A2(_1056_),
    .Z(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3777_ (.A1(_1036_),
    .A2(_1051_),
    .B(\dsynth.freeRunCntr[11] ),
    .ZN(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3778_ (.A1(\dsynth.freeRunCntr[11] ),
    .A2(_1037_),
    .A3(_1051_),
    .ZN(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3779_ (.A1(_1058_),
    .A2(_1054_),
    .B(_1060_),
    .ZN(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3780_ (.A1(_1057_),
    .A2(_1061_),
    .Z(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3781_ (.I(_1062_),
    .Z(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3782_ (.A1(_1050_),
    .A2(_1036_),
    .A3(_1005_),
    .ZN(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3783_ (.A1(_1136_),
    .A2(_1063_),
    .ZN(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3784_ (.A1(_1135_),
    .A2(_1063_),
    .Z(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3785_ (.A1(_1064_),
    .A2(_1065_),
    .ZN(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3786_ (.A1(_0697_),
    .A2(_1056_),
    .ZN(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3787_ (.A1(_1057_),
    .A2(_1061_),
    .B(_1067_),
    .ZN(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3788_ (.A1(_1066_),
    .A2(_1068_),
    .Z(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3789_ (.I(_1070_),
    .Z(_0004_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3790_ (.A1(_1050_),
    .A2(_1037_),
    .A3(_1011_),
    .ZN(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3791_ (.A1(_0849_),
    .A2(_1071_),
    .Z(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3792_ (.A1(_1066_),
    .A2(_1068_),
    .B(_1065_),
    .ZN(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3793_ (.A1(_1072_),
    .A2(_1073_),
    .Z(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3794_ (.I(_1074_),
    .Z(_0005_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3795_ (.A1(_0967_),
    .A2(_1022_),
    .Z(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3796_ (.A1(_0849_),
    .A2(_1071_),
    .ZN(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3797_ (.A1(_1072_),
    .A2(_1073_),
    .B(_1076_),
    .ZN(_1077_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3798_ (.A1(_1123_),
    .A2(_1075_),
    .A3(_1077_),
    .Z(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3799_ (.I(_1079_),
    .Z(_0006_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3800_ (.I(_1075_),
    .ZN(_1080_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3801_ (.A1(\dsynth.freeRunCntr[15] ),
    .A2(_1080_),
    .ZN(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3802_ (.A1(\dsynth.freeRunCntr[15] ),
    .A2(_1080_),
    .ZN(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3803_ (.A1(_1081_),
    .A2(_1077_),
    .B(_1082_),
    .ZN(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3804_ (.A1(_1131_),
    .A2(_1083_),
    .Z(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3805_ (.I(_1084_),
    .Z(_0007_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3806_ (.A1(\dsynth.freeRunCntr[16] ),
    .A2(_1083_),
    .Z(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3807_ (.A1(\dsynth.freeRunCntr[17] ),
    .A2(_1085_),
    .Z(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3808_ (.I(_1086_),
    .Z(_0008_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3809_ (.A1(\dsynth.freeRunCntr[17] ),
    .A2(_1085_),
    .ZN(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3810_ (.A1(_1145_),
    .A2(_1088_),
    .ZN(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3811_ (.I(_1089_),
    .Z(_0009_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3812_ (.I(_1144_),
    .ZN(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3813_ (.A1(_1145_),
    .A2(\dsynth.freeRunCntr[17] ),
    .A3(_1085_),
    .ZN(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3814_ (.A1(_1090_),
    .A2(_1091_),
    .Z(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3815_ (.I(_1092_),
    .Z(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3816_ (.I(_1157_),
    .Z(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3817_ (.A1(_1090_),
    .A2(_1091_),
    .ZN(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3818_ (.A1(_1093_),
    .A2(_1094_),
    .Z(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3819_ (.I(_1096_),
    .Z(_0012_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3820_ (.A1(_1093_),
    .A2(_1094_),
    .ZN(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3821_ (.A1(_0349_),
    .A2(_1097_),
    .ZN(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3822_ (.I(_1098_),
    .Z(_0013_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3823_ (.A1(_0349_),
    .A2(_1093_),
    .A3(_1094_),
    .ZN(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3824_ (.A1(\dsynth.csTable.address[4] ),
    .A2(_1099_),
    .ZN(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3825_ (.I(_1100_),
    .Z(_0014_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3826_ (.A1(_0349_),
    .A2(_1093_),
    .A3(\dsynth.csTable.address[4] ),
    .A4(_1094_),
    .Z(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3827_ (.A1(_0536_),
    .A2(_1101_),
    .Z(_1102_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3828_ (.I(_1102_),
    .Z(_0015_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3829_ (.A1(_0536_),
    .A2(_1101_),
    .ZN(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3830_ (.A1(_0085_),
    .A2(_1104_),
    .ZN(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3831_ (.I(_1105_),
    .Z(_0016_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3832_ (.A1(_1132_),
    .A2(_1104_),
    .ZN(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3833_ (.A1(_0112_),
    .A2(_1104_),
    .B(_1106_),
    .ZN(_0017_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3834_ (.A1(_0536_),
    .A2(_0085_),
    .A3(_1574_),
    .A4(_1101_),
    .Z(_1107_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3835_ (.A1(\dsynth.freeRunCntr[26] ),
    .A2(_1107_),
    .Z(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3836_ (.I(_1108_),
    .Z(_0018_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3837_ (.A1(\dsynth.freeRunCntr[26] ),
    .A2(_1107_),
    .Z(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3838_ (.A1(\dsynth.freeRunCntr[27] ),
    .A2(_1109_),
    .Z(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3839_ (.I(_1111_),
    .Z(_0019_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3840_ (.A1(\dsynth.freeRunCntr[27] ),
    .A2(_1109_),
    .Z(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3841_ (.A1(\dsynth.freeRunCntr[28] ),
    .A2(_1112_),
    .Z(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3842_ (.I(_1113_),
    .Z(_0020_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3843_ (.A1(\dsynth.freeRunCntr[28] ),
    .A2(_1112_),
    .B(_1477_),
    .ZN(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3844_ (.A1(_1477_),
    .A2(\dsynth.freeRunCntr[28] ),
    .A3(_1112_),
    .Z(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3845_ (.I(_1115_),
    .Z(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3846_ (.A1(_1114_),
    .A2(_1116_),
    .ZN(_0021_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3847_ (.A1(_1486_),
    .A2(_1116_),
    .Z(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3848_ (.I(_1117_),
    .Z(_0023_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3849_ (.A1(_1486_),
    .A2(_1116_),
    .B(_1476_),
    .ZN(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3850_ (.A1(_1485_),
    .A2(_1116_),
    .B(_1119_),
    .ZN(_0024_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3851_ (.A1(_1485_),
    .A2(_1115_),
    .ZN(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3852_ (.A1(_1473_),
    .A2(_1120_),
    .Z(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3853_ (.I(_1121_),
    .Z(_0025_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3854_ (.A1(\dsynth.freeRunCntr[0] ),
    .A2(_0972_),
    .Z(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3855_ (.I(_1122_),
    .Z(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3856_ (.I(net43),
    .ZN(_1919_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3857_ (.D(\tmux.clkapa ),
    .CLK(net43),
    .Q(\tmux.clkpaa ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3858_ (.D(\tmux.clkpaa ),
    .CLK(net44),
    .Q(\tmux.clkpab ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3859_ (.D(\tmux.clkbpb ),
    .CLK(net5),
    .Q(\tmux.clkpba ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3860_ (.D(\tmux.clkpba ),
    .CLK(net5),
    .Q(\tmux.clkpbb ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3861_ (.D(net6),
    .E(_1919_),
    .Q(\tgate.clkp ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3862_ (.D(_0000_),
    .RN(net53),
    .CLK(net41),
    .Q(\dsynth.freeRunCntr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3863_ (.D(_0011_),
    .RN(net54),
    .CLK(net41),
    .Q(\dsynth.freeRunCntr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3864_ (.D(_0022_),
    .RN(net55),
    .CLK(net40),
    .Q(\dsynth.freeRunCntr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3865_ (.D(_0026_),
    .RN(net55),
    .CLK(net42),
    .Q(\dsynth.freeRunCntr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3866_ (.D(_0027_),
    .RN(net55),
    .CLK(net40),
    .Q(\dsynth.freeRunCntr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3867_ (.D(_0028_),
    .RN(net55),
    .CLK(net40),
    .Q(\dsynth.freeRunCntr[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3868_ (.D(_0029_),
    .RN(net56),
    .CLK(net40),
    .Q(\dsynth.freeRunCntr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3869_ (.D(_0030_),
    .RN(net56),
    .CLK(net39),
    .Q(\dsynth.freeRunCntr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3870_ (.D(_0031_),
    .RN(net54),
    .CLK(net41),
    .Q(\dsynth.freeRunCntr[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3871_ (.D(_0032_),
    .RN(net53),
    .CLK(net37),
    .Q(\dsynth.freeRunCntr[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3872_ (.D(_0001_),
    .RN(net53),
    .CLK(net37),
    .Q(\dsynth.freeRunCntr[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3873_ (.D(_0002_),
    .RN(net53),
    .CLK(net37),
    .Q(\dsynth.freeRunCntr[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3874_ (.D(_0003_),
    .RN(net58),
    .CLK(net37),
    .Q(\dsynth.freeRunCntr[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3875_ (.D(_0004_),
    .RN(net58),
    .CLK(net38),
    .Q(\dsynth.freeRunCntr[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3876_ (.D(_0005_),
    .RN(net58),
    .CLK(net38),
    .Q(\dsynth.freeRunCntr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3877_ (.D(_0006_),
    .RN(net50),
    .CLK(net38),
    .Q(\dsynth.freeRunCntr[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3878_ (.D(_0007_),
    .RN(net50),
    .CLK(net33),
    .Q(\dsynth.freeRunCntr[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3879_ (.D(_0008_),
    .RN(net47),
    .CLK(net31),
    .Q(\dsynth.freeRunCntr[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3880_ (.D(_0009_),
    .RN(net47),
    .CLK(net31),
    .Q(\dsynth.csTable.address[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3881_ (.D(_0010_),
    .RN(net47),
    .CLK(net31),
    .Q(\dsynth.csTable.address[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3882_ (.D(_0012_),
    .RN(net47),
    .CLK(net31),
    .Q(\dsynth.csTable.address[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3883_ (.D(_0013_),
    .RN(net48),
    .CLK(net32),
    .Q(\dsynth.csTable.address[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3884_ (.D(_0014_),
    .RN(net48),
    .CLK(net32),
    .Q(\dsynth.csTable.address[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3885_ (.D(_0015_),
    .RN(net48),
    .CLK(net32),
    .Q(\dsynth.csTable.address[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3886_ (.D(_0016_),
    .RN(net52),
    .CLK(net36),
    .Q(\dsynth.csTable.address[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3887_ (.D(_0017_),
    .RN(net51),
    .CLK(net35),
    .Q(\dsynth.csTable.address[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3888_ (.D(_0018_),
    .RN(net49),
    .CLK(net33),
    .Q(\dsynth.freeRunCntr[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3889_ (.D(_0019_),
    .RN(net49),
    .CLK(net33),
    .Q(\dsynth.freeRunCntr[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3890_ (.D(_0020_),
    .RN(net49),
    .CLK(net33),
    .Q(\dsynth.freeRunCntr[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3891_ (.D(_0021_),
    .RN(net49),
    .CLK(net34),
    .Q(\dsynth.freeRunCntr[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3892_ (.D(_0023_),
    .RN(net51),
    .CLK(net35),
    .Q(\dsynth.freeRunCntr[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3893_ (.D(_0024_),
    .RN(net52),
    .CLK(net36),
    .Q(\dsynth.freeRunCntr[31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3894_ (.D(_0025_),
    .RN(net50),
    .CLK(net34),
    .Q(\dsynth.freeRunCntr[32] ));
 gf180mcu_fd_sc_mcu7t5v0__tieh user_proj_example_196 (.Z(net196));
 gf180mcu_fd_sc_mcu7t5v0__tieh user_proj_example_197 (.Z(net197));
 gf180mcu_fd_sc_mcu7t5v0__tieh user_proj_example_198 (.Z(net198));
 gf180mcu_fd_sc_mcu7t5v0__tieh user_proj_example_199 (.Z(net199));
 gf180mcu_fd_sc_mcu7t5v0__tieh user_proj_example_200 (.Z(net200));
 gf180mcu_fd_sc_mcu7t5v0__tieh user_proj_example_201 (.Z(net201));
 gf180mcu_fd_sc_mcu7t5v0__tieh user_proj_example_202 (.Z(net202));
 gf180mcu_fd_sc_mcu7t5v0__tieh user_proj_example_203 (.Z(net203));
 gf180mcu_fd_sc_mcu7t5v0__tieh user_proj_example_204 (.Z(net204));
 gf180mcu_fd_sc_mcu7t5v0__tieh user_proj_example_205 (.Z(net205));
 gf180mcu_fd_sc_mcu7t5v0__tieh user_proj_example_206 (.Z(net206));
 gf180mcu_fd_sc_mcu7t5v0__tieh user_proj_example_207 (.Z(net207));
 gf180mcu_fd_sc_mcu7t5v0__tieh user_proj_example_208 (.Z(net208));
 gf180mcu_fd_sc_mcu7t5v0__tieh user_proj_example_209 (.Z(net209));
 gf180mcu_fd_sc_mcu7t5v0__tieh user_proj_example_210 (.Z(net210));
 gf180mcu_fd_sc_mcu7t5v0__tieh user_proj_example_211 (.Z(net211));
 gf180mcu_fd_sc_mcu7t5v0__tieh user_proj_example_212 (.Z(net212));
 gf180mcu_fd_sc_mcu7t5v0__tieh user_proj_example_213 (.Z(net213));
 gf180mcu_fd_sc_mcu7t5v0__tieh user_proj_example_214 (.Z(net214));
 gf180mcu_fd_sc_mcu7t5v0__tieh user_proj_example_215 (.Z(net215));
 gf180mcu_fd_sc_mcu7t5v0__tieh user_proj_example_216 (.Z(net216));
 gf180mcu_fd_sc_mcu7t5v0__tieh user_proj_example_217 (.Z(net217));
 gf180mcu_fd_sc_mcu7t5v0__tieh user_proj_example_218 (.Z(net218));
 gf180mcu_fd_sc_mcu7t5v0__tieh user_proj_example_219 (.Z(net219));
 gf180mcu_fd_sc_mcu7t5v0__tieh user_proj_example_220 (.Z(net220));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3620__A2 (.I(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_61 (.ZN(net61));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_62 (.ZN(net62));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_63 (.ZN(net63));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_64 (.ZN(net64));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_65 (.ZN(net65));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_66 (.ZN(net66));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_67 (.ZN(net67));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_68 (.ZN(net68));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_69 (.ZN(net69));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_70 (.ZN(net70));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_71 (.ZN(net71));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_72 (.ZN(net72));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_73 (.ZN(net73));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_74 (.ZN(net74));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_75 (.ZN(net75));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_76 (.ZN(net76));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_77 (.ZN(net77));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_78 (.ZN(net78));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_79 (.ZN(net79));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_80 (.ZN(net80));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_81 (.ZN(net81));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_82 (.ZN(net82));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_83 (.ZN(net83));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_84 (.ZN(net84));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_85 (.ZN(net85));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_86 (.ZN(net86));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_87 (.ZN(net87));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_88 (.ZN(net88));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_89 (.ZN(net89));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_90 (.ZN(net90));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_91 (.ZN(net91));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_92 (.ZN(net92));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_93 (.ZN(net93));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_94 (.ZN(net94));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_95 (.ZN(net95));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_96 (.ZN(net96));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_97 (.ZN(net97));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_98 (.ZN(net98));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_99 (.ZN(net99));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_100 (.ZN(net100));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_101 (.ZN(net101));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_102 (.ZN(net102));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_103 (.ZN(net103));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_104 (.ZN(net104));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_105 (.ZN(net105));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_106 (.ZN(net106));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_107 (.ZN(net107));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_108 (.ZN(net108));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_109 (.ZN(net109));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_110 (.ZN(net110));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_111 (.ZN(net111));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_112 (.ZN(net112));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_113 (.ZN(net113));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_114 (.ZN(net114));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_115 (.ZN(net115));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_116 (.ZN(net116));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_117 (.ZN(net117));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_118 (.ZN(net118));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_119 (.ZN(net119));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_120 (.ZN(net120));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_121 (.ZN(net121));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_122 (.ZN(net122));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_123 (.ZN(net123));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_124 (.ZN(net124));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_125 (.ZN(net125));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_126 (.ZN(net126));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_127 (.ZN(net127));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_128 (.ZN(net128));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_129 (.ZN(net129));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_130 (.ZN(net130));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_131 (.ZN(net131));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_132 (.ZN(net132));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_133 (.ZN(net133));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_134 (.ZN(net134));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_135 (.ZN(net135));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_136 (.ZN(net136));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_137 (.ZN(net137));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_138 (.ZN(net138));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_139 (.ZN(net139));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_140 (.ZN(net140));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_141 (.ZN(net141));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_142 (.ZN(net142));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_143 (.ZN(net143));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_144 (.ZN(net144));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_145 (.ZN(net145));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_146 (.ZN(net146));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_147 (.ZN(net147));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_148 (.ZN(net148));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_149 (.ZN(net149));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_150 (.ZN(net150));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_151 (.ZN(net151));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_152 (.ZN(net152));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_153 (.ZN(net153));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_154 (.ZN(net154));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_155 (.ZN(net155));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_156 (.ZN(net156));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_157 (.ZN(net157));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_158 (.ZN(net158));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_159 (.ZN(net159));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_160 (.ZN(net160));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_161 (.ZN(net161));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_162 (.ZN(net162));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_163 (.ZN(net163));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_164 (.ZN(net164));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_165 (.ZN(net165));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_166 (.ZN(net166));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_167 (.ZN(net167));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_168 (.ZN(net168));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_169 (.ZN(net169));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_170 (.ZN(net170));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_171 (.ZN(net171));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_172 (.ZN(net172));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_173 (.ZN(net173));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_174 (.ZN(net174));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_175 (.ZN(net175));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_176 (.ZN(net176));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_177 (.ZN(net177));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_178 (.ZN(net178));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_179 (.ZN(net179));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_180 (.ZN(net180));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_181 (.ZN(net181));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_182 (.ZN(net182));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_183 (.ZN(net183));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_184 (.ZN(net184));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_185 (.ZN(net185));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_186 (.ZN(net186));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_187 (.ZN(net187));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_188 (.ZN(net188));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_189 (.ZN(net189));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_190 (.ZN(net190));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_191 (.ZN(net191));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_192 (.ZN(net192));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_193 (.ZN(net193));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_194 (.ZN(net194));
 gf180mcu_fd_sc_mcu7t5v0__tieh user_proj_example_195 (.Z(net195));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_289 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_290 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_291 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_292 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_293 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_294 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_295 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_296 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_297 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_298 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_299 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_300 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_301 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_302 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_303 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_304 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_305 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_306 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_307 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_308 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_309 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_310 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_311 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_312 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_313 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_314 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_315 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_316 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_317 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_318 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_319 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_320 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_321 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_322 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_323 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_324 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_325 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_326 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_327 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_328 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_329 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_330 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_331 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_332 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_333 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_334 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_335 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_336 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_337 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_338 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_339 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_340 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_341 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_342 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_343 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_344 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_345 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_346 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_347 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_348 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_349 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_350 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_351 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_352 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_353 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_354 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_355 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_356 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_357 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_358 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_359 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_360 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_361 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_362 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_363 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_364 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_365 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_366 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_367 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_368 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_369 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_370 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_371 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_372 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_373 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_374 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_375 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_376 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_377 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_378 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_379 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_380 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_381 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_382 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_383 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_384 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_385 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_386 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_387 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_388 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_389 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_390 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_391 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_392 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_393 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_394 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_395 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_396 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_397 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_398 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_399 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_400 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_401 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_402 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_403 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_404 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_405 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_406 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_407 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_408 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_409 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_410 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_411 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_412 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_413 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_414 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_415 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_416 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_417 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_418 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_419 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_420 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_421 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_422 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_423 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_424 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_425 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_426 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_427 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_428 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_429 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_430 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_431 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_432 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_433 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_434 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_435 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_436 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_437 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_438 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_439 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_440 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_441 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_442 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_443 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_444 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_445 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_446 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_447 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_448 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_449 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_450 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_451 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_452 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_453 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_454 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_455 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_456 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_457 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_458 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_459 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_460 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_461 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_462 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_463 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_464 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_465 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_466 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_467 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_468 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_469 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_470 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_471 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_472 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_473 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_474 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_475 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_476 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_477 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_478 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_479 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_480 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_481 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_482 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_483 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_484 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_485 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_486 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_487 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_488 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_489 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_490 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_491 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_492 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6595 ();
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1 (.I(io_in[11]),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input2 (.I(io_in[12]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input3 (.I(io_in[13]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input4 (.I(io_in[14]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input5 (.I(io_in[21]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input6 (.I(io_in[22]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input7 (.I(io_in[25]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input8 (.I(io_in[26]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input9 (.I(io_in[27]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input10 (.I(io_in[28]),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input11 (.I(io_in[35]),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input12 (.I(io_in[36]),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input13 (.I(io_in[37]),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input14 (.I(io_in[5]),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input15 (.I(io_in[6]),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output16 (.I(net16),
    .Z(io_out[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output17 (.I(net17),
    .Z(io_out[15]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output18 (.I(net18),
    .Z(io_out[16]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output19 (.I(net19),
    .Z(io_out[17]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output20 (.I(net20),
    .Z(io_out[18]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output21 (.I(net21),
    .Z(io_out[19]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output22 (.I(net22),
    .Z(io_out[20]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output23 (.I(net23),
    .Z(io_out[23]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output24 (.I(net24),
    .Z(io_out[24]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output25 (.I(net25),
    .Z(io_out[29]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output26 (.I(net26),
    .Z(io_out[30]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output27 (.I(net27),
    .Z(io_out[31]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output28 (.I(net28),
    .Z(io_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output29 (.I(net29),
    .Z(io_out[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output30 (.I(net30),
    .Z(io_out[9]));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout31 (.I(net32),
    .Z(net31));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout32 (.I(net36),
    .Z(net32));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout33 (.I(net35),
    .Z(net33));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout34 (.I(net35),
    .Z(net34));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout35 (.I(net36),
    .Z(net35));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout36 (.I(net39),
    .Z(net36));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout37 (.I(net38),
    .Z(net37));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout38 (.I(net39),
    .Z(net38));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout39 (.I(net46),
    .Z(net39));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout40 (.I(net41),
    .Z(net40));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout41 (.I(net42),
    .Z(net41));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout42 (.I(net45),
    .Z(net42));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout43 (.I(net44),
    .Z(net43));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout44 (.I(net45),
    .Z(net44));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout45 (.I(net46),
    .Z(net45));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout46 (.I(net13),
    .Z(net46));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout47 (.I(net48),
    .Z(net47));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout48 (.I(net52),
    .Z(net48));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout49 (.I(net51),
    .Z(net49));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout50 (.I(net51),
    .Z(net50));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout51 (.I(net52),
    .Z(net51));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout52 (.I(net59),
    .Z(net52));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout53 (.I(net57),
    .Z(net53));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout54 (.I(net57),
    .Z(net54));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout55 (.I(net56),
    .Z(net55));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout56 (.I(net57),
    .Z(net56));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout57 (.I(net58),
    .Z(net57));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout58 (.I(net59),
    .Z(net58));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout59 (.I(net12),
    .Z(net59));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_60 (.ZN(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2841__A2 (.I(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2831__A2 (.I(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2819__A2 (.I(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2832__A1 (.I(_0035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2823__A1 (.I(_0035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2822__A1 (.I(_0035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3616__A2 (.I(_0045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2946__A2 (.I(_0045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2831__B1 (.I(_0045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3640__B1 (.I(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2834__A1 (.I(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3243__A1 (.I(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3044__S (.I(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3042__B2 (.I(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2842__A2 (.I(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3066__B (.I(_0055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2976__A1 (.I(_0055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2912__I0 (.I(_0055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2841__B (.I(_0055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2848__A1 (.I(_0060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2847__A1 (.I(_0060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2848__A2 (.I(_0061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2847__A2 (.I(_0061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3204__A1 (.I(_0090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3202__I0 (.I(_0090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3139__A1 (.I(_0090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2873__A1 (.I(_0090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2906__A1 (.I(_0097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2881__A1 (.I(_0097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3100__A3 (.I(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3096__I (.I(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3062__A2 (.I(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2880__A2 (.I(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2907__A1 (.I(_0100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2898__A3 (.I(_0100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2883__A2 (.I(_0100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2893__A1 (.I(_0104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2891__A2 (.I(_0104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2890__A2 (.I(_0106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2022__I (.I(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1925__I (.I(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2893__A2 (.I(_0110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2891__A3 (.I(_0110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3833__A1 (.I(_0112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2957__B (.I(_0112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2956__A1 (.I(_0112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2893__B (.I(_0112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3066__A2 (.I(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3058__I (.I(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2896__A2 (.I(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3503__A1 (.I(_0129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3012__A1 (.I(_0129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2297__A1 (.I(_0129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1927__A2 (.I(_0129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3035__I1 (.I(_0130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3028__I (.I(_0130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2910__I0 (.I(_0130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3619__A2 (.I(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3035__I0 (.I(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3029__I1 (.I(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2910__I1 (.I(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2355__A1 (.I(_0140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2037__A1 (.I(_0140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2985__A1 (.I(_0142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2923__A1 (.I(_0142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2923__B (.I(_0145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3452__A2 (.I(_0159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2936__A2 (.I(_0159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3326__A1 (.I(_0160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2998__A1 (.I(_0160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3044__I1 (.I(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2970__A2 (.I(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2947__A2 (.I(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2964__A1 (.I(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2962__A3 (.I(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3139__B2 (.I(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3073__A1 (.I(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3021__A1 (.I(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2961__A1 (.I(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3261__I (.I(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3048__B1 (.I(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2960__A2 (.I(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3038__A1 (.I(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3011__I (.I(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2960__B (.I(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2520__B2 (.I(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2502__A2 (.I(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2220__B (.I(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1933__I (.I(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2293__C (.I(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2247__I (.I(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2080__A1 (.I(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1952__A1 (.I(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2983__A1 (.I(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2981__A1 (.I(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2983__A2 (.I(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2981__A2 (.I(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3188__A2 (.I(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3165__A2 (.I(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2988__A2 (.I(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2984__A2 (.I(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2547__A2 (.I(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2284__A2 (.I(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2245__A2 (.I(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1936__I (.I(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2422__A2 (.I(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2119__I (.I(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2045__A1 (.I(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1941__A1 (.I(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3297__A1 (.I(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3015__A1 (.I(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3013__A1 (.I(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3284__A2 (.I(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3106__A2 (.I(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3049__A2 (.I(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3018__A2 (.I(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3215__A1 (.I(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3203__A1 (.I(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3075__S (.I(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3020__S (.I(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3435__A2 (.I(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3431__A2 (.I(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3224__A2 (.I(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3025__A2 (.I(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3242__A2 (.I(_0260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3211__B (.I(_0260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3031__A2 (.I(_0260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3029__S (.I(_0260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3218__A1 (.I(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3039__A1 (.I(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3037__A1 (.I(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3301__A1 (.I(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3289__A2 (.I(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3262__A1 (.I(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3035__S (.I(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3218__A2 (.I(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3039__A2 (.I(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3037__A2 (.I(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2284__B (.I(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2103__A2 (.I(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1990__A2 (.I(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1940__I (.I(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3302__A1 (.I(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3288__A2 (.I(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3098__A2 (.I(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3042__A2 (.I(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3057__B2 (.I(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3046__A1 (.I(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3059__A3 (.I(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3045__A2 (.I(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3238__A1 (.I(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3061__A1 (.I(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3059__A1 (.I(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3048__A1 (.I(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2225__A2 (.I(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2144__I (.I(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2063__A2 (.I(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1941__A2 (.I(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3056__A1 (.I(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3055__A1 (.I(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3050__A2 (.I(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3084__I (.I(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3077__A1 (.I(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3057__A2 (.I(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3091__A1 (.I(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3071__A1 (.I(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2068__I (.I(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1951__A1 (.I(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3647__A2 (.I(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3613__A2 (.I(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3612__A2 (.I(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3059__B1 (.I(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3108__A1 (.I(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3069__A1 (.I(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3306__A1 (.I(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3305__A1 (.I(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3233__A1 (.I(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3069__A2 (.I(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3091__A2 (.I(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3071__A2 (.I(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3159__A2 (.I(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3117__A2 (.I(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3090__A2 (.I(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3288__A1 (.I(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3242__A1 (.I(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3211__A2 (.I(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3097__A2 (.I(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3134__A1 (.I(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3114__A1 (.I(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3121__A1 (.I(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3112__A1 (.I(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3232__A2 (.I(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3201__I (.I(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3110__S (.I(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2201__I (.I(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2111__I (.I(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2070__I (.I(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1949__B (.I(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3134__B (.I(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2588__A4 (.I(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2423__A1 (.I(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1950__I (.I(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3501__A2 (.I(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3446__B1 (.I(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3354__B1 (.I(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3150__I (.I(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3548__A2 (.I(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3182__A2 (.I(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3156__I (.I(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3151__A2 (.I(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3341__A2 (.I(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3327__A2 (.I(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3178__A2 (.I(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3157__A2 (.I(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3164__B (.I(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3189__A2 (.I(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3165__A3 (.I(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3186__A1 (.I(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3185__A1 (.I(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3171__A1 (.I(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2587__A1 (.I(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2422__B (.I(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2219__I (.I(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1956__I (.I(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3296__A1 (.I(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3287__A1 (.I(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3233__A2 (.I(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3202__I1 (.I(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2500__A1 (.I(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2418__A2 (.I(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2231__A3 (.I(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1957__I (.I(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3239__I0 (.I(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3238__A2 (.I(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3235__I (.I(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3212__A1 (.I(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3216__A1 (.I(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3214__A1 (.I(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2808__B2 (.I(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2304__I (.I(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2146__B2 (.I(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1968__A1 (.I(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3274__A3 (.I(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3246__A1 (.I(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3632__A2 (.I(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3611__A2 (.I(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3289__A1 (.I(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3241__A1 (.I(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2422__A1 (.I(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2225__A1 (.I(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2063__A1 (.I(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1960__I (.I(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3250__A1 (.I(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3248__A1 (.I(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2655__A2 (.I(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2200__A2 (.I(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2054__A1 (.I(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1962__A2 (.I(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3617__A2 (.I(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3612__B1 (.I(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3264__A1 (.I(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3263__A1 (.I(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2806__A1 (.I(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2285__I (.I(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1968__A2 (.I(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3317__B1 (.I(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3316__B (.I(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3281__A3 (.I(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3303__A1 (.I(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3301__A2 (.I(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3289__B1 (.I(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3286__A2 (.I(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3307__A2 (.I(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3300__A2 (.I(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3285__A2 (.I(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2294__A1 (.I(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2051__A1 (.I(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2002__I (.I(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1966__I (.I(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2458__B (.I(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2157__I (.I(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2058__A1 (.I(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1967__I (.I(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3322__A3 (.I(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3322__A4 (.I(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3400__B2 (.I(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3323__A2 (.I(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3414__A1 (.I(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3347__A1 (.I(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3404__A2 (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3346__B3 (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3339__A2 (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3527__A3 (.I(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3474__A3 (.I(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3347__B (.I(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3384__A2 (.I(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3380__A3 (.I(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3350__A3 (.I(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2172__A1 (.I(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2149__A1 (.I(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2038__I (.I(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1971__I (.I(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3388__A2 (.I(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3379__A2 (.I(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3351__B2 (.I(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3504__A2 (.I(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3454__A2 (.I(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3427__B2 (.I(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3358__B2 (.I(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2214__A1 (.I(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2180__I0 (.I(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2143__I (.I(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1975__A1 (.I(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3466__A2 (.I(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3465__A2 (.I(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3365__A3 (.I(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3492__A2 (.I(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3488__A2 (.I(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3478__A3 (.I(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3375__A2 (.I(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2451__A2 (.I(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2047__A2 (.I(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1979__I (.I(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1974__I (.I(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3743__A1 (.I(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3638__A1 (.I(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3383__A1 (.I(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3741__A1 (.I(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3618__A1 (.I(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3387__A1 (.I(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3383__B2 (.I(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3395__A2 (.I(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3387__B1 (.I(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3726__A1 (.I(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3618__B2 (.I(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3395__A1 (.I(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3387__B2 (.I(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3596__A1 (.I(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2742__B2 (.I(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2740__A1 (.I(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2523__A1 (.I(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1987__A1 (.I(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3417__A1 (.I(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3406__A1 (.I(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2437__B (.I(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2169__I (.I(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2103__B (.I(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1977__I (.I(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3647__A1 (.I(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3613__A1 (.I(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3612__A1 (.I(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3413__I (.I(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3606__A2 (.I(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3419__A2 (.I(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3416__A2 (.I(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3605__A2 (.I(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3418__A2 (.I(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2436__A1 (.I(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2054__B (.I(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2045__B (.I(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1978__I (.I(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3596__A2 (.I(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3639__B2 (.I(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3630__A1 (.I(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3599__B (.I(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3534__A1 (.I(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3458__A1 (.I(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3457__A1 (.I(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3432__A1 (.I(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2450__A1 (.I(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2204__A2 (.I(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2093__I (.I(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1987__A2 (.I(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3646__A2 (.I(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3626__A2 (.I(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3625__B1 (.I(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3429__A1 (.I(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3458__A2 (.I(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3457__A2 (.I(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3432__A2 (.I(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3459__A2 (.I(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3432__A3 (.I(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3639__B1 (.I(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3630__A2 (.I(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3436__A2 (.I(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3434__A2 (.I(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3451__A2 (.I(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3442__A2 (.I(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3447__A1 (.I(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3445__A1 (.I(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2094__I (.I(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2074__I (.I(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1981__I (.I(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3508__A1 (.I(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3456__A1 (.I(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3502__A3 (.I(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3455__A2 (.I(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2172__A2 (.I(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2149__A2 (.I(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2060__A2 (.I(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1982__I (.I(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3528__B (.I(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3481__A2 (.I(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3476__A2 (.I(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3590__A1 (.I(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3536__A1 (.I(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3491__A1 (.I(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3529__A3 (.I(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3482__A3 (.I(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3590__A2 (.I(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3536__A2 (.I(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3491__A2 (.I(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2950__A2 (.I(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2323__A2 (.I(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2254__A2 (.I(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1987__A3 (.I(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2523__B (.I(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2418__C (.I(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2078__I (.I(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1986__I (.I(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2654__C (.I(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2419__A1 (.I(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2253__I (.I(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1987__B (.I(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3581__A1 (.I(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3557__A1 (.I(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3531__A1 (.I(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2545__A1 (.I(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2172__B (.I(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2060__A1 (.I(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1990__B (.I(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3565__A1 (.I(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3549__A1 (.I(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2587__A2 (.I(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2469__A2 (.I(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2228__A1 (.I(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1998__A2 (.I(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3563__A1 (.I(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3560__A1 (.I(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2284__A1 (.I(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2117__I (.I(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2109__S (.I(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1994__A1 (.I(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3568__B (.I(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3597__A2 (.I(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3595__A2 (.I(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3639__A1 (.I(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3585__A1 (.I(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3771__A1 (.I(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3762__A1 (.I(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3585__B3 (.I(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3603__B (.I(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3610__B1 (.I(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3724__A1 (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3615__A1 (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3655__A1 (.I(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3630__B (.I(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2589__A1 (.I(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2001__B1 (.I(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3630__C (.I(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2500__B (.I(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2181__B (.I(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2058__A2 (.I(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2000__I (.I(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3655__A2 (.I(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2197__A1 (.I(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2159__A1 (.I(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2158__A1 (.I(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2001__B2 (.I(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3668__A1 (.I(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3666__B (.I(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3663__A1 (.I(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3659__A1 (.I(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3669__A1 (.I(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3662__A1 (.I(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3661__A1 (.I(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2622__A1 (.I(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2425__S (.I(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2258__I (.I(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2003__I (.I(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2228__C (.I(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2114__B (.I(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2080__C (.I(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2004__B2 (.I(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3747__A3 (.I(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3746__A2 (.I(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3688__A2 (.I(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2035__A2 (.I(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2005__A2 (.I(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3717__A2 (.I(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3716__A2 (.I(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3709__A2 (.I(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3446__A1 (.I(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3431__B2 (.I(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2720__A1 (.I(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2019__A2 (.I(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3737__I (.I(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3730__A1 (.I(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3724__A2 (.I(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3714__A1 (.I(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3724__A3 (.I(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3714__A2 (.I(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3733__A2 (.I(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3732__A2 (.I(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3726__A2 (.I(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2184__A1 (.I(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2086__I (.I(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2035__A1 (.I(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2009__I (.I(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3795__A2 (.I(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3740__A2 (.I(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2341__A1 (.I(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2326__A1 (.I(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2030__I (.I(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2017__A1 (.I(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3786__A2 (.I(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3776__A2 (.I(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2298__B (.I(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2178__B (.I(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2110__I (.I(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2014__I (.I(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3784__A2 (.I(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3783__A2 (.I(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2203__C (.I(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2153__C (.I(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2139__B (.I(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2015__A1 (.I(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3796__A2 (.I(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3791__A2 (.I(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3800__I (.I(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3798__A2 (.I(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3803__A2 (.I(_1077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3798__A3 (.I(_1077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3813__A3 (.I(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3809__A2 (.I(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3807__A2 (.I(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2763__A1 (.I(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2675__A1 (.I(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2600__A2 (.I(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2017__A2 (.I(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3624__A1 (.I(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3571__B (.I(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2028__B2 (.I(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2019__B2 (.I(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3626__A1 (.I(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3625__B2 (.I(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3567__A2 (.I(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2021__I (.I(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3798__A1 (.I(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3646__A1 (.I(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2031__B2 (.I(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2028__A1 (.I(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2271__A1 (.I(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2260__A1 (.I(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2234__A1 (.I(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2024__A1 (.I(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2025__A2 (.I(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3453__A1 (.I(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3435__A1 (.I(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2407__A1 (.I(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2027__I (.I(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3804__A1 (.I(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3646__B2 (.I(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3623__A1 (.I(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2031__A1 (.I(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3832__A1 (.I(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3548__A1 (.I(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3431__A1 (.I(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2031__A2 (.I(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3783__A1 (.I(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3569__A1 (.I(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3561__B (.I(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2036__A1 (.I(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2867__A1 (.I(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2764__A1 (.I(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2578__A1 (.I(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2036__A2 (.I(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2356__C (.I(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2355__B1 (.I(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2336__C (.I(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2244__A1 (.I(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2229__A1 (.I(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2041__A1 (.I(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2522__A1 (.I(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2306__A1 (.I(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2052__A1 (.I(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2249__I (.I(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2138__A2 (.I(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2045__A2 (.I(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2738__A1 (.I(_1148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2618__A1 (.I(_1148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2322__B (.I(_1148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2052__A2 (.I(_1148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2548__A1 (.I(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2544__A1 (.I(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2048__I (.I(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2621__A2 (.I(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2619__I0 (.I(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2438__A2 (.I(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2052__B1 (.I(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2544__A2 (.I(_1152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2288__B2 (.I(_1152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2052__B2 (.I(_1152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2652__A2 (.I(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2546__B2 (.I(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2052__C (.I(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2653__B2 (.I(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2458__A1 (.I(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2067__A1 (.I(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2148__A2 (.I(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2057__I (.I(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2505__A1 (.I(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2418__B1 (.I(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2079__B1 (.I(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2067__A2 (.I(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2623__A1 (.I(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2469__A3 (.I(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2206__B2 (.I(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2067__B (.I(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2519__B (.I(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2423__B2 (.I(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2159__A3 (.I(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2066__A2 (.I(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2196__B (.I(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2180__I1 (.I(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2073__I (.I(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2063__B (.I(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2504__A1 (.I(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2199__I (.I(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2066__B (.I(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2518__B (.I(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2266__B (.I(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2151__A2 (.I(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2065__I (.I(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2256__B (.I(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2191__A1 (.I(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2079__B2 (.I(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2066__C (.I(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2887__A1 (.I(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2742__A1 (.I(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2101__A2 (.I(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2072__A1 (.I(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2459__B (.I(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2416__A1 (.I(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2196__A1 (.I(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2071__A1 (.I(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2654__A1 (.I(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2458__A2 (.I(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2198__B2 (.I(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2072__A2 (.I(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2885__A1 (.I(_1174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2080__A2 (.I(_1174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2255__A1 (.I(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2221__I (.I(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2142__A2 (.I(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2076__A1 (.I(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2449__A1 (.I(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2180__S (.I(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2170__A2 (.I(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2075__I (.I(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2615__A2 (.I(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2231__A4 (.I(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2220__A3 (.I(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2076__A2 (.I(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2307__C (.I(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2178__C (.I(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2176__A1 (.I(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2079__A2 (.I(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2739__B (.I(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2481__A1 (.I(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2227__B (.I(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2079__C (.I(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2082__A2 (.I(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2805__A1 (.I(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2802__A1 (.I(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2579__A1 (.I(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2084__I (.I(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3446__B2 (.I(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3354__A1 (.I(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2129__A2 (.I(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2085__A2 (.I(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2439__B2 (.I(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2151__B (.I(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2104__I (.I(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2091__A2 (.I(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2656__C (.I(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2505__B2 (.I(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2092__I (.I(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2890__C2 (.I(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2461__A1 (.I(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2306__A2 (.I(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2124__A1 (.I(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2330__A2 (.I(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2192__I (.I(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2190__A3 (.I(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2096__A2 (.I(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2433__A1 (.I(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2298__A2 (.I(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2097__I (.I(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2334__A2 (.I(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2324__A2 (.I(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2106__B1 (.I(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2101__A3 (.I(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2518__A2 (.I(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2503__A2 (.I(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2204__A3 (.I(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2099__I (.I(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2889__A2 (.I(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2289__A2 (.I(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2270__C (.I(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2101__B2 (.I(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2739__A1 (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2319__A2 (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2159__A2 (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2106__A1 (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2433__A2 (.I(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2338__A2 (.I(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2153__B2 (.I(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2106__B2 (.I(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2740__C (.I(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2622__A2 (.I(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2616__B (.I(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2105__I (.I(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2810__A1 (.I(_1207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2809__A1 (.I(_1207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2274__A1 (.I(_1207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2106__C (.I(_1207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2655__B (.I(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2619__S (.I(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2420__A2 (.I(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2109__I1 (.I(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2806__B (.I(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2417__B1 (.I(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2203__B1 (.I(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2114__A1 (.I(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2268__I (.I(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2194__B (.I(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2120__B (.I(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2113__A1 (.I(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2524__A1 (.I(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2420__B (.I(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2200__B (.I(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2112__I (.I(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2230__A1 (.I(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2153__A1 (.I(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2120__A3 (.I(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2113__A2 (.I(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2501__C (.I(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2460__B (.I(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2182__B (.I(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2116__I (.I(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2309__I (.I(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2286__A1 (.I(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2206__A1 (.I(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2123__A1 (.I(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2617__A1 (.I(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2200__A1 (.I(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2151__A1 (.I(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2118__I (.I(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2953__A1 (.I(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2808__A1 (.I(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2256__A1 (.I(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2120__A1 (.I(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2273__C (.I(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2168__I (.I(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2122__I (.I(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2739__A2 (.I(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2338__A1 (.I(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2153__B1 (.I(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2123__A3 (.I(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2125__A2 (.I(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2404__A1 (.I(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2126__I (.I(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2938__A2 (.I(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2406__A1 (.I(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2394__A1 (.I(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2127__I (.I(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3354__B2 (.I(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2717__A1 (.I(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2167__A2 (.I(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2129__B1 (.I(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3640__B2 (.I(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3579__I (.I(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2130__I (.I(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2129__B2 (.I(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3773__A1 (.I(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3600__A1 (.I(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3578__B2 (.I(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2167__A1 (.I(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3641__A1 (.I(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3640__A1 (.I(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2187__A1 (.I(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2165__A1 (.I(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2524__B (.I(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2520__C (.I(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2502__A1 (.I(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2133__I (.I(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2482__A1 (.I(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2189__I (.I(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2183__A1 (.I(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2134__I (.I(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2888__B (.I(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2812__A1 (.I(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2494__A1 (.I(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2161__A1 (.I(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2273__A2 (.I(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2231__A2 (.I(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2220__A1 (.I(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2136__I (.I(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2336__B (.I(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2331__A1 (.I(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2225__B (.I(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2138__A1 (.I(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2452__A1 (.I(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2139__A2 (.I(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2952__A1 (.I(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2147__A1 (.I(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2524__A2 (.I(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2291__A2 (.I(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2148__A1 (.I(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2141__I (.I(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2621__A1 (.I(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2290__A2 (.I(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2153__A2 (.I(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2146__A1 (.I(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2810__A3 (.I(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2652__A1 (.I(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2146__A2 (.I(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2655__A1 (.I(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2265__A1 (.I(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2231__A1 (.I(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2145__A1 (.I(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2256__A2 (.I(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2255__A2 (.I(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2191__A2 (.I(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2145__A2 (.I(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2950__A3 (.I(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2333__B2 (.I(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2254__A3 (.I(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2146__B1 (.I(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2954__B1 (.I(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2307__A1 (.I(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2176__B1 (.I(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2152__A1 (.I(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2811__B1 (.I(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2619__I1 (.I(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2548__B1 (.I(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2150__I (.I(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2458__A3 (.I(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2308__A1 (.I(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2152__B (.I(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2622__A4 (.I(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2504__A2 (.I(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2171__A2 (.I(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2156__I (.I(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2740__A2 (.I(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2338__B1 (.I(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2270__A2 (.I(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2158__A2 (.I(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2324__B2 (.I(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2160__A2 (.I(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2161__B (.I(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2602__A1 (.I(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2163__I (.I(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3125__I0 (.I(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2937__A1 (.I(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2672__C2 (.I(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2164__I (.I(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2717__B2 (.I(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2570__A1 (.I(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2187__A2 (.I(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2165__A2 (.I(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2740__B2 (.I(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2521__A2 (.I(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2500__A3 (.I(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2171__A1 (.I(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2520__A2 (.I(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2423__C (.I(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2270__B (.I(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2171__B (.I(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2548__B2 (.I(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2438__A1 (.I(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2434__A3 (.I(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2176__A2 (.I(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2617__A3 (.I(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2523__A3 (.I(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2266__A2 (.I(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2175__A2 (.I(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2951__A2 (.I(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2293__A2 (.I(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2176__B2 (.I(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2621__B1 (.I(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2308__A2 (.I(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2181__A2 (.I(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2890__B2 (.I(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2182__A2 (.I(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2674__C2 (.I(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2661__A1 (.I(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2379__A1 (.I(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2185__I (.I(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2570__B2 (.I(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2356__A2 (.I(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2352__A2 (.I(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2187__B1 (.I(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3641__B2 (.I(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3593__A1 (.I(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3592__A1 (.I(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2187__B2 (.I(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3759__A1 (.I(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3642__A1 (.I(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2356__A1 (.I(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2352__A1 (.I(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2953__B (.I(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2288__A1 (.I(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2275__B (.I(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2207__A1 (.I(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2546__A2 (.I(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2275__A1 (.I(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2198__A1 (.I(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2456__A2 (.I(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2449__A2 (.I(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2240__A2 (.I(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2193__B (.I(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2436__A2 (.I(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2421__A2 (.I(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2233__A2 (.I(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2194__A2 (.I(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2950__B (.I(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2498__A1 (.I(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2251__A2 (.I(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2197__A2 (.I(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2889__B1 (.I(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2305__A2 (.I(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2270__A1 (.I(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2203__A1 (.I(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2651__A2 (.I(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2323__A3 (.I(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2203__A2 (.I(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2737__A2 (.I(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2208__A2 (.I(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3075__I0 (.I(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3010__A1 (.I(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2672__A1 (.I(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2210__I (.I(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2610__A1 (.I(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2358__A2 (.I(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2352__B1 (.I(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2239__A2 (.I(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3746__B (.I(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3635__B2 (.I(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2239__A1 (.I(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2212__I (.I(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2742__A2 (.I(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2423__A2 (.I(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2218__A2 (.I(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2588__A2 (.I(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2436__B (.I(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2433__C (.I(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2216__I (.I(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2653__C (.I(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2460__A1 (.I(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2424__A1 (.I(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2217__I (.I(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2811__C (.I(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2620__B2 (.I(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2319__A1 (.I(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2218__B (.I(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2743__B (.I(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2224__B1 (.I(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2886__A1 (.I(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2319__A3 (.I(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2290__A1 (.I(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2223__A1 (.I(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2433__B1 (.I(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2223__B (.I(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2224__B2 (.I(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2418__B2 (.I(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2293__B1 (.I(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2228__A2 (.I(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2651__A1 (.I(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2319__A4 (.I(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2241__A1 (.I(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2227__A3 (.I(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2889__A1 (.I(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2500__A2 (.I(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2289__A1 (.I(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2230__A2 (.I(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2494__A3 (.I(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2481__A2 (.I(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2470__B (.I(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2233__B (.I(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2885__B (.I(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2548__C (.I(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2233__C (.I(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2815__A1 (.I(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2799__A1 (.I(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2236__I (.I(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3106__A1 (.I(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3072__A1 (.I(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2674__A1 (.I(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2237__I (.I(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2672__B2 (.I(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2360__A2 (.I(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2350__A2 (.I(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2239__B1 (.I(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2740__B1 (.I(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2519__A2 (.I(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2248__A1 (.I(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2523__A2 (.I(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2298__A1 (.I(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2273__B (.I(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2243__A2 (.I(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2653__A1 (.I(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2322__A1 (.I(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2246__A1 (.I(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2811__A2 (.I(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2522__A2 (.I(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2246__A2 (.I(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2616__A1 (.I(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2542__A1 (.I(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2318__A1 (.I(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2246__B2 (.I(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2653__A2 (.I(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2420__A1 (.I(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2301__I (.I(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2250__A2 (.I(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2295__A3 (.I(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2259__A1 (.I(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2810__A2 (.I(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2469__A1 (.I(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2290__B (.I(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2254__A1 (.I(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2305__B (.I(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2264__A2 (.I(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2257__A2 (.I(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2333__A1 (.I(_1359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2259__B1 (.I(_1359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2809__B (.I(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2302__I (.I(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2295__A1 (.I(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2259__C (.I(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2895__A1 (.I(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2869__A1 (.I(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2262__I (.I(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3018__A1 (.I(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2765__A1 (.I(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2674__B2 (.I(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2263__I (.I(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3020__I0 (.I(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2360__B1 (.I(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2350__C1 (.I(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2281__A2 (.I(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2954__A2 (.I(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2293__B2 (.I(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2267__A1 (.I(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2654__B (.I(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2334__A3 (.I(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2267__A2 (.I(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2953__C (.I(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2332__I (.I(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2307__B (.I(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2269__B (.I(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2497__A1 (.I(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2418__A1 (.I(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2291__A1 (.I(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2273__A1 (.I(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2656__B (.I(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2274__A3 (.I(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2277__A2 (.I(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3341__A1 (.I(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2940__A1 (.I(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2347__B1 (.I(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2281__B1 (.I(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3619__A1 (.I(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3386__I (.I(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2347__B2 (.I(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2281__B2 (.I(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3616__A1 (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3421__A1 (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3411__A1 (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2316__A1 (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2433__B2 (.I(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2298__A3 (.I(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2288__A2 (.I(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2953__A2 (.I(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2889__B2 (.I(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2807__A1 (.I(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2288__C (.I(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2806__C (.I(_1393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2457__A2 (.I(_1393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2292__I (.I(_1393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2951__A1 (.I(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2807__A2 (.I(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2321__A1 (.I(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2293__A1 (.I(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2744__A1 (.I(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2522__A3 (.I(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2453__B (.I(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2295__B2 (.I(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2871__A2 (.I(_1398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2297__A2 (.I(_1398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3327__A1 (.I(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3126__A1 (.I(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2347__A2 (.I(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2316__A2 (.I(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2501__A1 (.I(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2311__A1 (.I(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2588__A3 (.I(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2300__I (.I(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2808__A2 (.I(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2622__A3 (.I(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2457__A1 (.I(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2303__A1 (.I(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2954__A1 (.I(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2886__A2 (.I(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2322__A2 (.I(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2303__A2 (.I(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2340__B2 (.I(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2335__A1 (.I(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2323__A1 (.I(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2303__B (.I(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2312__A2 (.I(_1413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3088__A1 (.I(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3067__A1 (.I(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2313__I (.I(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3267__I (.I(_1415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3232__A1 (.I(_1415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2941__A1 (.I(_1415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2314__I (.I(_1415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3182__A1 (.I(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2365__A2 (.I(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2346__A2 (.I(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2316__B1 (.I(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3717__A1 (.I(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2361__I (.I(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2346__A1 (.I(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2316__B2 (.I(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3707__A1 (.I(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3412__I (.I(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2344__A1 (.I(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2329__A1 (.I(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2326__A2 (.I(_1427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3166__A1 (.I(_1428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3123__A1 (.I(_1428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3049__A1 (.I(_1428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2327__I (.I(_1428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3286__A1 (.I(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3284__A1 (.I(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3025__A1 (.I(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2328__I (.I(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3178__A1 (.I(_1430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3157__A1 (.I(_1430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2344__A2 (.I(_1430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2329__A2 (.I(_1430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2499__A2 (.I(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2333__A2 (.I(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2331__A2 (.I(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2439__A1 (.I(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2333__B1 (.I(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2460__A2 (.I(_1438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2337__A2 (.I(_1438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3012__A2 (.I(_1442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2341__A2 (.I(_1442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3087__A1 (.I(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2342__I (.I(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3224__A1 (.I(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3151__A1 (.I(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2364__A2 (.I(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2344__B1 (.I(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3700__A1 (.I(_1445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3612__B2 (.I(_1445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2363__I (.I(_1445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2344__B2 (.I(_1445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2355__B2 (.I(_1456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3632__A1 (.I(_1463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3611__A1 (.I(_1463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3411__B2 (.I(_1463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2362__I (.I(_1463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3709__A1 (.I(_1464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3607__A1 (.I(_1464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3420__A1 (.I(_1464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2365__A1 (.I(_1464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3617__A1 (.I(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3605__A1 (.I(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3418__A1 (.I(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2364__A1 (.I(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2367__A3 (.I(_1468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2368__A2 (.I(_1469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2369__I (.I(_1470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3852__A1 (.I(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2541__A1 (.I(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2413__A3 (.I(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2378__A1 (.I(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3844__A1 (.I(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3843__B (.I(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2399__A1 (.I(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2377__A2 (.I(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2765__A2 (.I(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2565__I (.I(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2379__A2 (.I(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2428__A2 (.I(_1483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2383__I (.I(_1483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3851__A1 (.I(_1485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3850__A1 (.I(_1485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2444__A2 (.I(_1485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2387__A2 (.I(_1485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3849__A1 (.I(_1486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3847__A1 (.I(_1486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2568__A1 (.I(_1486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2386__A1 (.I(_1486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2762__A2 (.I(_1488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2388__A2 (.I(_1488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2799__A2 (.I(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2389__I (.I(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2748__A2 (.I(_1491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2604__A2 (.I(_1491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2578__A2 (.I(_1491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2391__I (.I(_1491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3109__A2 (.I(_1492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2959__A2 (.I(_1492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2763__A2 (.I(_1492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2392__I (.I(_1492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3205__A2 (.I(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3015__A2 (.I(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3013__A2 (.I(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2393__A2 (.I(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2397__I (.I(_1494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2394__B (.I(_1494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2562__A2 (.I(_1495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2395__A2 (.I(_1495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3435__C (.I(_1498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2675__A2 (.I(_1498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2609__A1 (.I(_1498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2409__A1 (.I(_1498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2661__A2 (.I(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2514__A2 (.I(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2403__I (.I(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2400__I (.I(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3358__C (.I(_1503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2668__A1 (.I(_1503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2608__B2 (.I(_1503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2408__A1 (.I(_1503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3074__A2 (.I(_1504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2895__A2 (.I(_1504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2406__A2 (.I(_1504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2404__A2 (.I(_1504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2882__A1 (.I(_1506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2867__A2 (.I(_1506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2817__A1 (.I(_1506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2408__A2 (.I(_1506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3088__B (.I(_1507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2407__A2 (.I(_1507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2411__A2 (.I(_1510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2410__A2 (.I(_1510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2960__A1 (.I(_1514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2896__A1 (.I(_1514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2816__A1 (.I(_1514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2414__I (.I(_1514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3547__A2 (.I(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2720__B2 (.I(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2579__B1 (.I(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2466__A1 (.I(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2892__I (.I(_1516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2483__A1 (.I(_1516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2462__B (.I(_1516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2426__A1 (.I(_1516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2887__A2 (.I(_1523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2742__A3 (.I(_1523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2423__B1 (.I(_1523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2425__I1 (.I(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3061__A2 (.I(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2834__A2 (.I(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2752__A1 (.I(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2427__I (.I(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3635__A2 (.I(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3059__A2 (.I(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3030__A2 (.I(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2466__A2 (.I(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2774__A1 (.I(_1530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2529__I (.I(_1530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2430__I (.I(_1530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2831__B2 (.I(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2583__A2 (.I(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2466__B1 (.I(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2435__A2 (.I(_1534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2656__A1 (.I(_1538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2621__B2 (.I(_1538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2542__A2 (.I(_1538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2438__B2 (.I(_1538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2441__A2 (.I(_1540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2440__A3 (.I(_1540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2974__I1 (.I(_1543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2686__I0 (.I(_1543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2443__I (.I(_1543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3637__A2 (.I(_1544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3635__B1 (.I(_1544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2665__A2 (.I(_1544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2466__B2 (.I(_1544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2819__A1 (.I(_1547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2752__A2 (.I(_1547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2665__A1 (.I(_1547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2447__I (.I(_1547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3429__A2 (.I(_1549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3361__A2 (.I(_1549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3048__B2 (.I(_1549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2466__C1 (.I(_1549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2808__B1 (.I(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2450__A2 (.I(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2546__B1 (.I(_1552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2452__A2 (.I(_1552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2955__A1 (.I(_1553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2453__A2 (.I(_1553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2497__A2 (.I(_1555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2459__A2 (.I(_1555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2456__A1 (.I(_1555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2455__A2 (.I(_1555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2742__B1 (.I(_1556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2457__B (.I(_1556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2464__A3 (.I(_1562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2462__A2 (.I(_1562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2582__I (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2480__A1 (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2466__C2 (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2745__A1 (.I(_1569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2624__B (.I(_1569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2495__A1 (.I(_1569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2471__A1 (.I(_1569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2474__A2 (.I(_1571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2471__A3 (.I(_1571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2658__A1 (.I(_1573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2507__B (.I(_1573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2506__A1 (.I(_1573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2473__I (.I(_1573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3834__A3 (.I(_1574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2879__A1 (.I(_1574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2746__B (.I(_1574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2474__B (.I(_1574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3454__A1 (.I(_1576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3427__C2 (.I(_1576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2636__A1 (.I(_1576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2492__A1 (.I(_1576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2685__B (.I(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2630__A1 (.I(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2477__I (.I(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3047__I (.I(_1579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2834__B (.I(_1579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2484__A1 (.I(_1579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2479__I (.I(_1579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3030__A1 (.I(_1580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2841__A1 (.I(_1580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2537__A1 (.I(_1580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2480__A2 (.I(_1580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2911__B2 (.I(_1581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2492__A2 (.I(_1581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2533__A2 (.I(_1583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2483__A2 (.I(_1583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3428__I (.I(_1584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2509__I1 (.I(_1584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2484__A2 (.I(_1584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3625__A2 (.I(_1586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3624__A2 (.I(_1586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3361__A1 (.I(_1586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2491__I0 (.I(_1586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2973__A1 (.I(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2908__B (.I(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2838__B (.I(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2487__B (.I(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2776__A1 (.I(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2751__A1 (.I(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2493__I (.I(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2490__B (.I(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2536__A2 (.I(_1595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2495__A2 (.I(_1595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3627__A2 (.I(_1596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3504__B2 (.I(_1596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3427__A1 (.I(_1596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2496__A2 (.I(_1596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2505__B1 (.I(_1605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2777__A1 (.I(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2776__B (.I(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2534__I (.I(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2509__S (.I(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2868__A1 (.I(_1615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2821__A1 (.I(_1615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2563__I (.I(_1615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2531__A1 (.I(_1615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2748__B1 (.I(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2662__A1 (.I(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2516__I (.I(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3060__A2 (.I(_1618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2975__A1 (.I(_1618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2687__A1 (.I(_1618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2530__A2 (.I(_1618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2884__A1 (.I(_1619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2806__A2 (.I(_1619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2520__A1 (.I(_1619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2527__A2 (.I(_1626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2526__A3 (.I(_1626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2628__B1 (.I(_1629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2576__I (.I(_1629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2530__B1 (.I(_1629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2970__A1 (.I(_1630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2880__A1 (.I(_1630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2753__A1 (.I(_1630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2530__B2 (.I(_1630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2564__A2 (.I(_1631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2531__A2 (.I(_1631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2659__B (.I(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2625__A1 (.I(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2612__A1 (.I(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2533__A1 (.I(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3504__A1 (.I(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3454__B2 (.I(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2751__A2 (.I(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2538__A1 (.I(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3097__B (.I(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2913__A1 (.I(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2842__B2 (.I(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2538__A2 (.I(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2891__A1 (.I(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2814__A1 (.I(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2590__A1 (.I(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2536__A1 (.I(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2572__A1 (.I(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2557__A1 (.I(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3639__A2 (.I(_1640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3358__B1 (.I(_1640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2722__A1 (.I(_1640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2556__A1 (.I(_1640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3097__A1 (.I(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2878__A1 (.I(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2584__I (.I(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2556__A2 (.I(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2955__B2 (.I(_1644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2589__A2 (.I(_1644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2544__B (.I(_1644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2951__B2 (.I(_1648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2548__A2 (.I(_1648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2946__B (.I(_1653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2778__A1 (.I(_1653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2581__A2 (.I(_1653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2553__A2 (.I(_1653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3433__I (.I(_1655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3360__A2 (.I(_1655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2585__A2 (.I(_1655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2555__A2 (.I(_1655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2572__A2 (.I(_1657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2557__A2 (.I(_1657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3125__S (.I(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2937__A2 (.I(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2749__A1 (.I(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2564__A1 (.I(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2712__A1 (.I(_1665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2711__A1 (.I(_1665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2571__A2 (.I(_1665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3087__A2 (.I(_1666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2941__A2 (.I(_1666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2674__A2 (.I(_1666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2566__I (.I(_1666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3166__A2 (.I(_1667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3123__A2 (.I(_1667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2672__A2 (.I(_1667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2567__I (.I(_1667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3453__A2 (.I(_1668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3431__C2 (.I(_1668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2716__I (.I(_1668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2570__A2 (.I(_1668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2935__A2 (.I(_1669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2569__A2 (.I(_1669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2674__B1 (.I(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2672__B1 (.I(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2599__I (.I(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2570__B1 (.I(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3126__A2 (.I(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3088__A2 (.I(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2674__C1 (.I(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2575__I (.I(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3023__I (.I(_1676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2720__A2 (.I(_1676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2672__C1 (.I(_1676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2579__A2 (.I(_1676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3642__A2 (.I(_1678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3641__B1 (.I(_1678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3048__A2 (.I(_1678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2579__B2 (.I(_1678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3646__B1 (.I(_1681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3623__A2 (.I(_1681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3547__A1 (.I(_1681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2581__A1 (.I(_1681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2718__A1 (.I(_1682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2594__A1 (.I(_1682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3641__A2 (.I(_1683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3640__A2 (.I(_1683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2720__B1 (.I(_1683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2583__A1 (.I(_1683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3100__A1 (.I(_1687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3062__B (.I(_1687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3060__A1 (.I(_1687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2591__A1 (.I(_1687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2637__A2 (.I(_1692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2592__A2 (.I(_1692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3431__B1 (.I(_1700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3149__I (.I(_1700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2717__B1 (.I(_1700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2610__A2 (.I(_1700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3452__A1 (.I(_1702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3358__A1 (.I(_1702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2667__I1 (.I(_1702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2608__A1 (.I(_1702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2667__S (.I(_1703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2606__I (.I(_1703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2603__I (.I(_1703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3125__I1 (.I(_1704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3107__B2 (.I(_1704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2897__A1 (.I(_1704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2608__A2 (.I(_1704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2868__A2 (.I(_1706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2805__A2 (.I(_1706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2720__C (.I(_1706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2607__A1 (.I(_1706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3076__A1 (.I(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2962__A1 (.I(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2948__A1 (.I(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2607__A2 (.I(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3638__A2 (.I(_1714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3100__A2 (.I(_1714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3062__A1 (.I(_1714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2628__A1 (.I(_1714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3098__A1 (.I(_1715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2947__A1 (.I(_1715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2664__I (.I(_1715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2628__A2 (.I(_1715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2620__B1 (.I(_1720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2625__A2 (.I(_1721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2624__A1 (.I(_1721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3618__A2 (.I(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3033__A2 (.I(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2666__A2 (.I(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2628__C1 (.I(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3627__B1 (.I(_1730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3624__B1 (.I(_1730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2682__I1 (.I(_1730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2630__A2 (.I(_1730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2878__B (.I(_1732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2687__B1 (.I(_1732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2682__I0 (.I(_1732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2634__A1 (.I(_1732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2910__S (.I(_1733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2682__S (.I(_1733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2633__I (.I(_1733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3102__A1 (.I(_1734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2975__B2 (.I(_1734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2911__A1 (.I(_1734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2634__A2 (.I(_1734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3043__A1 (.I(_1736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3034__A1 (.I(_1736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3032__I (.I(_1736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2636__A2 (.I(_1736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2831__C (.I(_1737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2637__B2 (.I(_1737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2659__A2 (.I(_1758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2658__A3 (.I(_1758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2750__I (.I(_1761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2662__A2 (.I(_1761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3141__A1 (.I(_1762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3111__A1 (.I(_1762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2949__I (.I(_1762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2662__B (.I(_1762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3437__A1 (.I(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2756__I (.I(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2722__A2 (.I(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2666__A1 (.I(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2690__A2 (.I(_1766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2666__A3 (.I(_1766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2820__A1 (.I(_1782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2724__B (.I(_1782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2688__A1 (.I(_1782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2683__A1 (.I(_1782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2836__B (.I(_1785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2835__A1 (.I(_1785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2687__A2 (.I(_1785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3015__A3 (.I(_1786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3014__A1 (.I(_1786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2974__I0 (.I(_1786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2686__I1 (.I(_1786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2700__A1 (.I(_1798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2699__A1 (.I(_1798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2700__A2 (.I(_1799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2699__A2 (.I(_1799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3479__A1 (.I(_1807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3351__A1 (.I(_1807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2735__A1 (.I(_1807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3502__A2 (.I(_1817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3446__A2 (.I(_1817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3354__A2 (.I(_1817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2717__A2 (.I(_1817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3478__A1 (.I(_1834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3353__A1 (.I(_1834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2734__A1 (.I(_1834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3205__A1 (.I(_1838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3107__A1 (.I(_1838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2763__B2 (.I(_1838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2748__A1 (.I(_1838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2741__A2 (.I(_1840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2744__A2 (.I(_1843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2746__A2 (.I(_1845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2745__A3 (.I(_1845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3615__A2 (.I(_1848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3210__A2 (.I(_1848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2820__B (.I(_1848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2748__B2 (.I(_1848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3361__B (.I(_1852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2752__B (.I(_1852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3436__A1 (.I(_1857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3426__I (.I(_1857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3360__A1 (.I(_1857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2758__A1 (.I(_1857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3618__B1 (.I(_1858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3031__A1 (.I(_1858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2911__A2 (.I(_1858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2758__A2 (.I(_1858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2769__A1 (.I(_1860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2761__A1 (.I(_1860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3358__A2 (.I(_1863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2763__B1 (.I(_1863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2768__A1 (.I(_1864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2766__A1 (.I(_1864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2800__A1 (.I(_1865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2768__A2 (.I(_1865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2766__A2 (.I(_1865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2781__A2 (.I(_1880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2780__A2 (.I(_1880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2850__A1 (.I(_1883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2785__A1 (.I(_1883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2784__A1 (.I(_1883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2850__A2 (.I(_1884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2785__A2 (.I(_1884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2784__A2 (.I(_1884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2789__A2 (.I(_1888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2788__A2 (.I(_1888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3067__A2 (.I(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3017__I (.I(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2938__B (.I(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2798__B (.I(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3503__A2 (.I(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2901__A2 (.I(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2873__A2 (.I(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2804__A2 (.I(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2857__A1 (.I(_1906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2827__A1 (.I(_1906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3209__I (.I(_1915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3061__A3 (.I(_1915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2816__A2 (.I(_1915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3019__I (.I(_1916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2816__B (.I(_1916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2898__A2 (.I(_1917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2882__A2 (.I(_1917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2817__A2 (.I(_1917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2095__A2 (.I(\dsynth.csTable.address[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2055__I (.I(\dsynth.csTable.address[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1972__A2 (.I(\dsynth.csTable.address[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1934__A2 (.I(\dsynth.csTable.address[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1953__A2 (.I(\dsynth.csTable.address[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1946__I (.I(\dsynth.csTable.address[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1969__A1 (.I(\dsynth.csTable.address[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1942__I (.I(\dsynth.csTable.address[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1928__I (.I(\dsynth.csTable.address[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1921__I (.I(\dsynth.csTable.address[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3578__A1 (.I(\dsynth.freeRunCntr[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3424__I (.I(\dsynth.freeRunCntr[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2129__A1 (.I(\dsynth.freeRunCntr[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2085__A1 (.I(\dsynth.freeRunCntr[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3627__B2 (.I(\dsynth.freeRunCntr[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3624__B2 (.I(\dsynth.freeRunCntr[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2033__I (.I(\dsynth.freeRunCntr[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2019__A1 (.I(\dsynth.freeRunCntr[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3625__A1 (.I(\dsynth.freeRunCntr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3562__I (.I(\dsynth.freeRunCntr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2018__I (.I(\dsynth.freeRunCntr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3715__A1 (.I(\dsynth.freeRunCntr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3614__I (.I(\dsynth.freeRunCntr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2347__A1 (.I(\dsynth.freeRunCntr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2283__I (.I(\dsynth.freeRunCntr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3731__A1 (.I(\dsynth.freeRunCntr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3382__I (.I(\dsynth.freeRunCntr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2349__I (.I(\dsynth.freeRunCntr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2281__A1 (.I(\dsynth.freeRunCntr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3750__A1 (.I(\dsynth.freeRunCntr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3749__A1 (.I(\dsynth.freeRunCntr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3635__A1 (.I(\dsynth.freeRunCntr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2238__I (.I(\dsynth.freeRunCntr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(io_in[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(io_in[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(io_in[21]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(io_in[22]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(io_in[25]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(io_in[26]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(io_in[27]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(io_in[28]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input11_I (.I(io_in[35]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input12_I (.I(io_in[36]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input13_I (.I(io_in[37]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input14_I (.I(io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input15_I (.I(io_in[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3675__A3 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3669__A2 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3667__B (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3665__B (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3672__C (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3670__B (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3664__I (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3672__A1 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3670__A1 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3667__A1 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3665__A1 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3860__CLK (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3859__CLK (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3676__B1 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3861__D (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3680__A2 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3678__I (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3690__I (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3685__I (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3695__I (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3691__A1 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3687__A1 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3691__A3 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3686__I (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3675__A1 (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3672__B (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3660__I (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3657__I (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout59_I (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout46_I (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3663__A2 (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3662__A2 (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3658__I (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3663__A3 (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3662__A3 (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3661__A3 (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3659__A3 (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output16_I (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output17_I (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output18_I (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output19_I (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output20_I (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output21_I (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output22_I (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output25_I (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output26_I (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output28_I (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output30_I (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3882__CLK (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3881__CLK (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3880__CLK (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3879__CLK (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3885__CLK (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3883__CLK (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3884__CLK (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout31_I (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3890__CLK (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3878__CLK (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3889__CLK (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3888__CLK (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3892__CLK (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3887__CLK (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout33_I (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout34_I (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3893__CLK (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout35_I (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3886__CLK (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout32_I (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3874__CLK (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3873__CLK (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3872__CLK (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3871__CLK (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout37_I (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3877__CLK (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3876__CLK (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3875__CLK (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3869__CLK (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout38_I (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout36_I (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3864__CLK (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3868__CLK (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3867__CLK (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3866__CLK (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout40_I (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3870__CLK (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3863__CLK (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3862__CLK (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3676__A1 (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3857__CLK (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3856__I (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3681__A1 (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3858__CLK (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout43_I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout44_I (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout42_I (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout45_I (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout39_I (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3882__RN (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3881__RN (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3880__RN (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3879__RN (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3885__RN (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3883__RN (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3884__RN (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout47_I (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3891__RN (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3890__RN (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3889__RN (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3888__RN (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3894__RN (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3878__RN (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3877__RN (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3892__RN (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3887__RN (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout49_I (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout50_I (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3893__RN (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout51_I (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3886__RN (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout48_I (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3862__RN (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3873__RN (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3872__RN (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3871__RN (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3867__RN (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3866__RN (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3865__RN (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3864__RN (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3868__RN (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout55_I (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3869__RN (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout56_I (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout53_I (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout54_I (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout57_I (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3876__RN (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3875__RN (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3874__RN (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout58_I (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout52_I (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_145_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_145_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_145_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_145_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_146_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_146_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_147_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_147_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_147_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_147_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_148_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_149_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_149_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_149_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_149_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_149_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_150_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_150_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_151_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_151_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_151_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_152_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_153_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_153_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_153_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_153_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_153_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_153_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_154_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_154_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_154_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_154_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_154_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_154_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_154_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_154_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_154_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_155_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_155_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_155_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_156_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_156_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_156_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_157_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_157_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_158_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_158_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_158_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_159_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_159_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_159_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_159_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_159_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_159_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_160_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_160_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_161_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_161_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_162_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_162_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_163_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_163_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_163_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_164_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_165_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_165_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_165_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_165_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_165_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_165_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_165_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_165_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_165_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_165_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_165_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_166_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_166_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_167_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_167_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_167_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_168_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_168_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_168_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_169_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_170_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_170_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_170_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_171_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_171_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_171_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_171_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_171_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_171_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_171_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_172_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_172_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_172_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_172_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_173_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_173_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_173_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_173_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_173_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_173_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_173_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_173_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_173_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_173_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_174_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_174_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_174_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_174_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_174_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_174_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_174_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_175_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_175_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_175_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_175_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_176_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_177_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_177_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_177_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_177_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_177_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_177_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_177_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_177_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_178_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_178_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_179_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_179_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_179_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_179_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_179_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_180_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_180_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_180_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_181_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_181_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_181_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_181_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_181_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_181_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_181_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_181_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_181_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_182_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_182_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_182_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_182_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_182_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_183_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_183_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_183_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_183_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_184_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_184_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_184_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_184_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_184_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_185_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_185_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_186_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_186_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_187_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_187_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_188_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_188_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_189_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_189_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_190_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_190_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_191_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_191_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_192_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_192_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_192_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_193_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_193_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_193_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_193_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_193_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_194_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_194_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_195_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_195_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_196_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_196_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_197_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_197_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_198_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_198_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_199_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_199_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_200_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_200_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_201_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_202_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_202_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_203_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_203_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_204_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_204_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_205_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_205_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_206_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_206_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_207_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_207_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_208_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_208_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_209_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_209_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_210_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_210_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_210_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_211_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_211_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_211_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_211_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_211_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_212_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_212_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_213_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_213_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_214_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_214_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_215_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_215_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_216_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_216_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_217_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_217_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_218_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_218_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_218_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_218_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_218_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_219_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_219_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_220_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_220_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_221_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_221_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_222_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_222_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_223_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_223_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_224_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_224_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_225_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_225_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_226_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_226_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_227_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_227_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_228_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_228_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_228_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_229_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_229_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_229_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_229_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_230_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_231_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_231_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_231_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_232_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_232_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_233_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_234_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_234_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_234_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_235_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_236_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_236_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_236_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_236_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_237_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_237_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_237_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_238_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_238_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_239_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_239_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_239_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_239_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_240_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_240_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_241_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_241_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_241_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_241_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_242_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_242_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_242_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_243_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_243_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_243_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_243_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_243_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_243_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_244_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_244_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_244_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_244_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_244_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_244_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_244_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_245_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_245_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_245_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_245_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_245_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1758 ();
 assign io_oeb[0] = net195;
 assign io_oeb[10] = net63;
 assign io_oeb[11] = net202;
 assign io_oeb[12] = net203;
 assign io_oeb[13] = net204;
 assign io_oeb[14] = net205;
 assign io_oeb[15] = net64;
 assign io_oeb[16] = net65;
 assign io_oeb[17] = net66;
 assign io_oeb[18] = net67;
 assign io_oeb[19] = net68;
 assign io_oeb[1] = net196;
 assign io_oeb[20] = net69;
 assign io_oeb[21] = net206;
 assign io_oeb[22] = net207;
 assign io_oeb[23] = net70;
 assign io_oeb[24] = net71;
 assign io_oeb[25] = net208;
 assign io_oeb[26] = net209;
 assign io_oeb[27] = net210;
 assign io_oeb[28] = net211;
 assign io_oeb[29] = net72;
 assign io_oeb[2] = net197;
 assign io_oeb[30] = net73;
 assign io_oeb[31] = net74;
 assign io_oeb[32] = net212;
 assign io_oeb[33] = net213;
 assign io_oeb[34] = net214;
 assign io_oeb[35] = net215;
 assign io_oeb[36] = net216;
 assign io_oeb[37] = net217;
 assign io_oeb[3] = net198;
 assign io_oeb[4] = net199;
 assign io_oeb[5] = net200;
 assign io_oeb[6] = net201;
 assign io_oeb[7] = net60;
 assign io_oeb[8] = net61;
 assign io_oeb[9] = net62;
 assign io_out[0] = net75;
 assign io_out[11] = net82;
 assign io_out[12] = net83;
 assign io_out[13] = net84;
 assign io_out[14] = net85;
 assign io_out[1] = net76;
 assign io_out[21] = net86;
 assign io_out[22] = net87;
 assign io_out[25] = net88;
 assign io_out[26] = net89;
 assign io_out[27] = net90;
 assign io_out[28] = net91;
 assign io_out[2] = net77;
 assign io_out[32] = net218;
 assign io_out[33] = net219;
 assign io_out[34] = net220;
 assign io_out[35] = net92;
 assign io_out[36] = net93;
 assign io_out[37] = net94;
 assign io_out[3] = net78;
 assign io_out[4] = net79;
 assign io_out[5] = net80;
 assign io_out[6] = net81;
 assign irq[0] = net95;
 assign irq[1] = net96;
 assign irq[2] = net97;
 assign la_data_out[0] = net98;
 assign la_data_out[10] = net108;
 assign la_data_out[11] = net109;
 assign la_data_out[12] = net110;
 assign la_data_out[13] = net111;
 assign la_data_out[14] = net112;
 assign la_data_out[15] = net113;
 assign la_data_out[16] = net114;
 assign la_data_out[17] = net115;
 assign la_data_out[18] = net116;
 assign la_data_out[19] = net117;
 assign la_data_out[1] = net99;
 assign la_data_out[20] = net118;
 assign la_data_out[21] = net119;
 assign la_data_out[22] = net120;
 assign la_data_out[23] = net121;
 assign la_data_out[24] = net122;
 assign la_data_out[25] = net123;
 assign la_data_out[26] = net124;
 assign la_data_out[27] = net125;
 assign la_data_out[28] = net126;
 assign la_data_out[29] = net127;
 assign la_data_out[2] = net100;
 assign la_data_out[30] = net128;
 assign la_data_out[31] = net129;
 assign la_data_out[32] = net130;
 assign la_data_out[33] = net131;
 assign la_data_out[34] = net132;
 assign la_data_out[35] = net133;
 assign la_data_out[36] = net134;
 assign la_data_out[37] = net135;
 assign la_data_out[38] = net136;
 assign la_data_out[39] = net137;
 assign la_data_out[3] = net101;
 assign la_data_out[40] = net138;
 assign la_data_out[41] = net139;
 assign la_data_out[42] = net140;
 assign la_data_out[43] = net141;
 assign la_data_out[44] = net142;
 assign la_data_out[45] = net143;
 assign la_data_out[46] = net144;
 assign la_data_out[47] = net145;
 assign la_data_out[48] = net146;
 assign la_data_out[49] = net147;
 assign la_data_out[4] = net102;
 assign la_data_out[50] = net148;
 assign la_data_out[51] = net149;
 assign la_data_out[52] = net150;
 assign la_data_out[53] = net151;
 assign la_data_out[54] = net152;
 assign la_data_out[55] = net153;
 assign la_data_out[56] = net154;
 assign la_data_out[57] = net155;
 assign la_data_out[58] = net156;
 assign la_data_out[59] = net157;
 assign la_data_out[5] = net103;
 assign la_data_out[60] = net158;
 assign la_data_out[61] = net159;
 assign la_data_out[62] = net160;
 assign la_data_out[63] = net161;
 assign la_data_out[6] = net104;
 assign la_data_out[7] = net105;
 assign la_data_out[8] = net106;
 assign la_data_out[9] = net107;
 assign wbs_ack_o = net162;
 assign wbs_dat_o[0] = net163;
 assign wbs_dat_o[10] = net173;
 assign wbs_dat_o[11] = net174;
 assign wbs_dat_o[12] = net175;
 assign wbs_dat_o[13] = net176;
 assign wbs_dat_o[14] = net177;
 assign wbs_dat_o[15] = net178;
 assign wbs_dat_o[16] = net179;
 assign wbs_dat_o[17] = net180;
 assign wbs_dat_o[18] = net181;
 assign wbs_dat_o[19] = net182;
 assign wbs_dat_o[1] = net164;
 assign wbs_dat_o[20] = net183;
 assign wbs_dat_o[21] = net184;
 assign wbs_dat_o[22] = net185;
 assign wbs_dat_o[23] = net186;
 assign wbs_dat_o[24] = net187;
 assign wbs_dat_o[25] = net188;
 assign wbs_dat_o[26] = net189;
 assign wbs_dat_o[27] = net190;
 assign wbs_dat_o[28] = net191;
 assign wbs_dat_o[29] = net192;
 assign wbs_dat_o[2] = net165;
 assign wbs_dat_o[30] = net193;
 assign wbs_dat_o[31] = net194;
 assign wbs_dat_o[3] = net166;
 assign wbs_dat_o[4] = net167;
 assign wbs_dat_o[5] = net168;
 assign wbs_dat_o[6] = net169;
 assign wbs_dat_o[7] = net170;
 assign wbs_dat_o[8] = net171;
 assign wbs_dat_o[9] = net172;
endmodule

