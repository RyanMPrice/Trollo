magic
tech gf180mcuC
magscale 1 5
timestamp 1670260625
<< metal1 >>
rect 672 6285 7360 6302
rect 672 6259 2259 6285
rect 2285 6259 2311 6285
rect 2337 6259 2363 6285
rect 2389 6259 3911 6285
rect 3937 6259 3963 6285
rect 3989 6259 4015 6285
rect 4041 6259 5563 6285
rect 5589 6259 5615 6285
rect 5641 6259 5667 6285
rect 5693 6259 7215 6285
rect 7241 6259 7267 6285
rect 7293 6259 7319 6285
rect 7345 6259 7360 6285
rect 672 6242 7360 6259
rect 4321 6063 4327 6089
rect 4353 6063 4359 6089
rect 4097 6007 4103 6033
rect 4129 6007 4135 6033
rect 672 5893 7280 5910
rect 672 5867 1433 5893
rect 1459 5867 1485 5893
rect 1511 5867 1537 5893
rect 1563 5867 3085 5893
rect 3111 5867 3137 5893
rect 3163 5867 3189 5893
rect 3215 5867 4737 5893
rect 4763 5867 4789 5893
rect 4815 5867 4841 5893
rect 4867 5867 6389 5893
rect 6415 5867 6441 5893
rect 6467 5867 6493 5893
rect 6519 5867 7280 5893
rect 672 5850 7280 5867
rect 672 5501 7360 5518
rect 672 5475 2259 5501
rect 2285 5475 2311 5501
rect 2337 5475 2363 5501
rect 2389 5475 3911 5501
rect 3937 5475 3963 5501
rect 3989 5475 4015 5501
rect 4041 5475 5563 5501
rect 5589 5475 5615 5501
rect 5641 5475 5667 5501
rect 5693 5475 7215 5501
rect 7241 5475 7267 5501
rect 7293 5475 7319 5501
rect 7345 5475 7360 5501
rect 672 5458 7360 5475
rect 672 5109 7280 5126
rect 672 5083 1433 5109
rect 1459 5083 1485 5109
rect 1511 5083 1537 5109
rect 1563 5083 3085 5109
rect 3111 5083 3137 5109
rect 3163 5083 3189 5109
rect 3215 5083 4737 5109
rect 4763 5083 4789 5109
rect 4815 5083 4841 5109
rect 4867 5083 6389 5109
rect 6415 5083 6441 5109
rect 6467 5083 6493 5109
rect 6519 5083 7280 5109
rect 672 5066 7280 5083
rect 672 4717 7360 4734
rect 672 4691 2259 4717
rect 2285 4691 2311 4717
rect 2337 4691 2363 4717
rect 2389 4691 3911 4717
rect 3937 4691 3963 4717
rect 3989 4691 4015 4717
rect 4041 4691 5563 4717
rect 5589 4691 5615 4717
rect 5641 4691 5667 4717
rect 5693 4691 7215 4717
rect 7241 4691 7267 4717
rect 7293 4691 7319 4717
rect 7345 4691 7360 4717
rect 672 4674 7360 4691
rect 4271 4633 4297 4639
rect 4271 4601 4297 4607
rect 3319 4521 3345 4527
rect 3145 4495 3151 4521
rect 3177 4495 3183 4521
rect 3319 4489 3345 4495
rect 3655 4521 3681 4527
rect 3655 4489 3681 4495
rect 3711 4521 3737 4527
rect 3711 4489 3737 4495
rect 3823 4521 3849 4527
rect 3823 4489 3849 4495
rect 3879 4521 3905 4527
rect 3879 4489 3905 4495
rect 3263 4465 3289 4471
rect 3263 4433 3289 4439
rect 3767 4465 3793 4471
rect 3767 4433 3793 4439
rect 4215 4465 4241 4471
rect 4215 4433 4241 4439
rect 672 4325 7280 4342
rect 672 4299 1433 4325
rect 1459 4299 1485 4325
rect 1511 4299 1537 4325
rect 1563 4299 3085 4325
rect 3111 4299 3137 4325
rect 3163 4299 3189 4325
rect 3215 4299 4737 4325
rect 4763 4299 4789 4325
rect 4815 4299 4841 4325
rect 4867 4299 6389 4325
rect 6415 4299 6441 4325
rect 6467 4299 6493 4325
rect 6519 4299 7280 4325
rect 672 4282 7280 4299
rect 1633 4159 1639 4185
rect 1665 4159 1671 4185
rect 3257 4159 3263 4185
rect 3289 4159 3295 4185
rect 2927 4129 2953 4135
rect 4713 4103 4719 4129
rect 4745 4103 4751 4129
rect 2927 4097 2953 4103
rect 961 4047 967 4073
rect 993 4047 999 4073
rect 4321 4047 4327 4073
rect 4353 4047 4359 4073
rect 2983 4017 3009 4023
rect 2983 3985 3009 3991
rect 672 3933 7360 3950
rect 672 3907 2259 3933
rect 2285 3907 2311 3933
rect 2337 3907 2363 3933
rect 2389 3907 3911 3933
rect 3937 3907 3963 3933
rect 3989 3907 4015 3933
rect 4041 3907 5563 3933
rect 5589 3907 5615 3933
rect 5641 3907 5667 3933
rect 5693 3907 7215 3933
rect 7241 3907 7267 3933
rect 7293 3907 7319 3933
rect 7345 3907 7360 3933
rect 672 3890 7360 3907
rect 911 3849 937 3855
rect 911 3817 937 3823
rect 4943 3849 4969 3855
rect 4943 3817 4969 3823
rect 4999 3849 5025 3855
rect 4999 3817 5025 3823
rect 3033 3711 3039 3737
rect 3065 3711 3071 3737
rect 4887 3681 4913 3687
rect 3369 3655 3375 3681
rect 3401 3655 3407 3681
rect 4433 3655 4439 3681
rect 4465 3655 4471 3681
rect 4887 3649 4913 3655
rect 672 3541 7280 3558
rect 672 3515 1433 3541
rect 1459 3515 1485 3541
rect 1511 3515 1537 3541
rect 1563 3515 3085 3541
rect 3111 3515 3137 3541
rect 3163 3515 3189 3541
rect 3215 3515 4737 3541
rect 4763 3515 4789 3541
rect 4815 3515 4841 3541
rect 4867 3515 6389 3541
rect 6415 3515 6441 3541
rect 6467 3515 6493 3541
rect 6519 3515 7280 3541
rect 672 3498 7280 3515
rect 3593 3375 3599 3401
rect 3625 3375 3631 3401
rect 4657 3319 4663 3345
rect 4689 3319 4695 3345
rect 5049 3319 5055 3345
rect 5081 3319 5087 3345
rect 672 3149 7360 3166
rect 672 3123 2259 3149
rect 2285 3123 2311 3149
rect 2337 3123 2363 3149
rect 2389 3123 3911 3149
rect 3937 3123 3963 3149
rect 3989 3123 4015 3149
rect 4041 3123 5563 3149
rect 5589 3123 5615 3149
rect 5641 3123 5667 3149
rect 5693 3123 7215 3149
rect 7241 3123 7267 3149
rect 7293 3123 7319 3149
rect 7345 3123 7360 3149
rect 672 3106 7360 3123
rect 3145 2983 3151 3009
rect 3177 2983 3183 3009
rect 2809 2927 2815 2953
rect 2841 2927 2847 2953
rect 4209 2871 4215 2897
rect 4241 2871 4247 2897
rect 672 2757 7280 2774
rect 672 2731 1433 2757
rect 1459 2731 1485 2757
rect 1511 2731 1537 2757
rect 1563 2731 3085 2757
rect 3111 2731 3137 2757
rect 3163 2731 3189 2757
rect 3215 2731 4737 2757
rect 4763 2731 4789 2757
rect 4815 2731 4841 2757
rect 4867 2731 6389 2757
rect 6415 2731 6441 2757
rect 6467 2731 6493 2757
rect 6519 2731 7280 2757
rect 672 2714 7280 2731
rect 672 2365 7360 2382
rect 672 2339 2259 2365
rect 2285 2339 2311 2365
rect 2337 2339 2363 2365
rect 2389 2339 3911 2365
rect 3937 2339 3963 2365
rect 3989 2339 4015 2365
rect 4041 2339 5563 2365
rect 5589 2339 5615 2365
rect 5641 2339 5667 2365
rect 5693 2339 7215 2365
rect 7241 2339 7267 2365
rect 7293 2339 7319 2365
rect 7345 2339 7360 2365
rect 672 2322 7360 2339
rect 672 1973 7280 1990
rect 672 1947 1433 1973
rect 1459 1947 1485 1973
rect 1511 1947 1537 1973
rect 1563 1947 3085 1973
rect 3111 1947 3137 1973
rect 3163 1947 3189 1973
rect 3215 1947 4737 1973
rect 4763 1947 4789 1973
rect 4815 1947 4841 1973
rect 4867 1947 6389 1973
rect 6415 1947 6441 1973
rect 6467 1947 6493 1973
rect 6519 1947 7280 1973
rect 672 1930 7280 1947
rect 2473 1807 2479 1833
rect 2505 1807 2511 1833
rect 5441 1807 5447 1833
rect 5473 1807 5479 1833
rect 2815 1721 2841 1727
rect 6399 1721 6425 1727
rect 1969 1695 1975 1721
rect 2001 1695 2007 1721
rect 5945 1695 5951 1721
rect 5977 1695 5983 1721
rect 2815 1689 2841 1695
rect 6399 1689 6425 1695
rect 672 1581 7360 1598
rect 672 1555 2259 1581
rect 2285 1555 2311 1581
rect 2337 1555 2363 1581
rect 2389 1555 3911 1581
rect 3937 1555 3963 1581
rect 3989 1555 4015 1581
rect 4041 1555 5563 1581
rect 5589 1555 5615 1581
rect 5641 1555 5667 1581
rect 5693 1555 7215 1581
rect 7241 1555 7267 1581
rect 7293 1555 7319 1581
rect 7345 1555 7360 1581
rect 672 1538 7360 1555
<< via1 >>
rect 2259 6259 2285 6285
rect 2311 6259 2337 6285
rect 2363 6259 2389 6285
rect 3911 6259 3937 6285
rect 3963 6259 3989 6285
rect 4015 6259 4041 6285
rect 5563 6259 5589 6285
rect 5615 6259 5641 6285
rect 5667 6259 5693 6285
rect 7215 6259 7241 6285
rect 7267 6259 7293 6285
rect 7319 6259 7345 6285
rect 4327 6063 4353 6089
rect 4103 6007 4129 6033
rect 1433 5867 1459 5893
rect 1485 5867 1511 5893
rect 1537 5867 1563 5893
rect 3085 5867 3111 5893
rect 3137 5867 3163 5893
rect 3189 5867 3215 5893
rect 4737 5867 4763 5893
rect 4789 5867 4815 5893
rect 4841 5867 4867 5893
rect 6389 5867 6415 5893
rect 6441 5867 6467 5893
rect 6493 5867 6519 5893
rect 2259 5475 2285 5501
rect 2311 5475 2337 5501
rect 2363 5475 2389 5501
rect 3911 5475 3937 5501
rect 3963 5475 3989 5501
rect 4015 5475 4041 5501
rect 5563 5475 5589 5501
rect 5615 5475 5641 5501
rect 5667 5475 5693 5501
rect 7215 5475 7241 5501
rect 7267 5475 7293 5501
rect 7319 5475 7345 5501
rect 1433 5083 1459 5109
rect 1485 5083 1511 5109
rect 1537 5083 1563 5109
rect 3085 5083 3111 5109
rect 3137 5083 3163 5109
rect 3189 5083 3215 5109
rect 4737 5083 4763 5109
rect 4789 5083 4815 5109
rect 4841 5083 4867 5109
rect 6389 5083 6415 5109
rect 6441 5083 6467 5109
rect 6493 5083 6519 5109
rect 2259 4691 2285 4717
rect 2311 4691 2337 4717
rect 2363 4691 2389 4717
rect 3911 4691 3937 4717
rect 3963 4691 3989 4717
rect 4015 4691 4041 4717
rect 5563 4691 5589 4717
rect 5615 4691 5641 4717
rect 5667 4691 5693 4717
rect 7215 4691 7241 4717
rect 7267 4691 7293 4717
rect 7319 4691 7345 4717
rect 4271 4607 4297 4633
rect 3151 4495 3177 4521
rect 3319 4495 3345 4521
rect 3655 4495 3681 4521
rect 3711 4495 3737 4521
rect 3823 4495 3849 4521
rect 3879 4495 3905 4521
rect 3263 4439 3289 4465
rect 3767 4439 3793 4465
rect 4215 4439 4241 4465
rect 1433 4299 1459 4325
rect 1485 4299 1511 4325
rect 1537 4299 1563 4325
rect 3085 4299 3111 4325
rect 3137 4299 3163 4325
rect 3189 4299 3215 4325
rect 4737 4299 4763 4325
rect 4789 4299 4815 4325
rect 4841 4299 4867 4325
rect 6389 4299 6415 4325
rect 6441 4299 6467 4325
rect 6493 4299 6519 4325
rect 1639 4159 1665 4185
rect 3263 4159 3289 4185
rect 2927 4103 2953 4129
rect 4719 4103 4745 4129
rect 967 4047 993 4073
rect 4327 4047 4353 4073
rect 2983 3991 3009 4017
rect 2259 3907 2285 3933
rect 2311 3907 2337 3933
rect 2363 3907 2389 3933
rect 3911 3907 3937 3933
rect 3963 3907 3989 3933
rect 4015 3907 4041 3933
rect 5563 3907 5589 3933
rect 5615 3907 5641 3933
rect 5667 3907 5693 3933
rect 7215 3907 7241 3933
rect 7267 3907 7293 3933
rect 7319 3907 7345 3933
rect 911 3823 937 3849
rect 4943 3823 4969 3849
rect 4999 3823 5025 3849
rect 3039 3711 3065 3737
rect 3375 3655 3401 3681
rect 4439 3655 4465 3681
rect 4887 3655 4913 3681
rect 1433 3515 1459 3541
rect 1485 3515 1511 3541
rect 1537 3515 1563 3541
rect 3085 3515 3111 3541
rect 3137 3515 3163 3541
rect 3189 3515 3215 3541
rect 4737 3515 4763 3541
rect 4789 3515 4815 3541
rect 4841 3515 4867 3541
rect 6389 3515 6415 3541
rect 6441 3515 6467 3541
rect 6493 3515 6519 3541
rect 3599 3375 3625 3401
rect 4663 3319 4689 3345
rect 5055 3319 5081 3345
rect 2259 3123 2285 3149
rect 2311 3123 2337 3149
rect 2363 3123 2389 3149
rect 3911 3123 3937 3149
rect 3963 3123 3989 3149
rect 4015 3123 4041 3149
rect 5563 3123 5589 3149
rect 5615 3123 5641 3149
rect 5667 3123 5693 3149
rect 7215 3123 7241 3149
rect 7267 3123 7293 3149
rect 7319 3123 7345 3149
rect 3151 2983 3177 3009
rect 2815 2927 2841 2953
rect 4215 2871 4241 2897
rect 1433 2731 1459 2757
rect 1485 2731 1511 2757
rect 1537 2731 1563 2757
rect 3085 2731 3111 2757
rect 3137 2731 3163 2757
rect 3189 2731 3215 2757
rect 4737 2731 4763 2757
rect 4789 2731 4815 2757
rect 4841 2731 4867 2757
rect 6389 2731 6415 2757
rect 6441 2731 6467 2757
rect 6493 2731 6519 2757
rect 2259 2339 2285 2365
rect 2311 2339 2337 2365
rect 2363 2339 2389 2365
rect 3911 2339 3937 2365
rect 3963 2339 3989 2365
rect 4015 2339 4041 2365
rect 5563 2339 5589 2365
rect 5615 2339 5641 2365
rect 5667 2339 5693 2365
rect 7215 2339 7241 2365
rect 7267 2339 7293 2365
rect 7319 2339 7345 2365
rect 1433 1947 1459 1973
rect 1485 1947 1511 1973
rect 1537 1947 1563 1973
rect 3085 1947 3111 1973
rect 3137 1947 3163 1973
rect 3189 1947 3215 1973
rect 4737 1947 4763 1973
rect 4789 1947 4815 1973
rect 4841 1947 4867 1973
rect 6389 1947 6415 1973
rect 6441 1947 6467 1973
rect 6493 1947 6519 1973
rect 2479 1807 2505 1833
rect 5447 1807 5473 1833
rect 1975 1695 2001 1721
rect 2815 1695 2841 1721
rect 5951 1695 5977 1721
rect 6399 1695 6425 1721
rect 2259 1555 2285 1581
rect 2311 1555 2337 1581
rect 2363 1555 2389 1581
rect 3911 1555 3937 1581
rect 3963 1555 3989 1581
rect 4015 1555 4041 1581
rect 5563 1555 5589 1581
rect 5615 1555 5641 1581
rect 5667 1555 5693 1581
rect 7215 1555 7241 1581
rect 7267 1555 7293 1581
rect 7319 1555 7345 1581
<< metal2 >>
rect 3976 7600 4032 8000
rect 3990 6874 4018 7600
rect 3990 6846 4130 6874
rect 2258 6286 2390 6291
rect 2286 6258 2310 6286
rect 2338 6258 2362 6286
rect 2258 6253 2390 6258
rect 3910 6286 4042 6291
rect 3938 6258 3962 6286
rect 3990 6258 4014 6286
rect 3910 6253 4042 6258
rect 4102 6033 4130 6846
rect 5562 6286 5694 6291
rect 5590 6258 5614 6286
rect 5642 6258 5666 6286
rect 5562 6253 5694 6258
rect 7214 6286 7346 6291
rect 7242 6258 7266 6286
rect 7294 6258 7318 6286
rect 7214 6253 7346 6258
rect 4102 6007 4103 6033
rect 4129 6007 4130 6033
rect 4102 6001 4130 6007
rect 4326 6089 4354 6095
rect 4326 6063 4327 6089
rect 4353 6063 4354 6089
rect 1432 5894 1564 5899
rect 1460 5866 1484 5894
rect 1512 5866 1536 5894
rect 1432 5861 1564 5866
rect 3084 5894 3216 5899
rect 4326 5894 4354 6063
rect 3112 5866 3136 5894
rect 3164 5866 3188 5894
rect 3084 5861 3216 5866
rect 4270 5866 4354 5894
rect 4736 5894 4868 5899
rect 4764 5866 4788 5894
rect 4816 5866 4840 5894
rect 2258 5502 2390 5507
rect 2286 5474 2310 5502
rect 2338 5474 2362 5502
rect 2258 5469 2390 5474
rect 3910 5502 4042 5507
rect 3938 5474 3962 5502
rect 3990 5474 4014 5502
rect 3910 5469 4042 5474
rect 1432 5110 1564 5115
rect 1460 5082 1484 5110
rect 1512 5082 1536 5110
rect 1432 5077 1564 5082
rect 3084 5110 3216 5115
rect 3112 5082 3136 5110
rect 3164 5082 3188 5110
rect 3084 5077 3216 5082
rect 2258 4718 2390 4723
rect 2286 4690 2310 4718
rect 2338 4690 2362 4718
rect 2258 4685 2390 4690
rect 3910 4718 4042 4723
rect 3938 4690 3962 4718
rect 3990 4690 4014 4718
rect 3910 4685 4042 4690
rect 4270 4633 4298 5866
rect 4736 5861 4868 5866
rect 6388 5894 6520 5899
rect 6416 5866 6440 5894
rect 6468 5866 6492 5894
rect 6388 5861 6520 5866
rect 5562 5502 5694 5507
rect 5590 5474 5614 5502
rect 5642 5474 5666 5502
rect 5562 5469 5694 5474
rect 7214 5502 7346 5507
rect 7242 5474 7266 5502
rect 7294 5474 7318 5502
rect 7214 5469 7346 5474
rect 4736 5110 4868 5115
rect 4764 5082 4788 5110
rect 4816 5082 4840 5110
rect 4736 5077 4868 5082
rect 6388 5110 6520 5115
rect 6416 5082 6440 5110
rect 6468 5082 6492 5110
rect 6388 5077 6520 5082
rect 5562 4718 5694 4723
rect 5590 4690 5614 4718
rect 5642 4690 5666 4718
rect 5562 4685 5694 4690
rect 7214 4718 7346 4723
rect 7242 4690 7266 4718
rect 7294 4690 7318 4718
rect 7214 4685 7346 4690
rect 4270 4607 4271 4633
rect 4297 4607 4298 4633
rect 4270 4601 4298 4607
rect 3150 4522 3178 4527
rect 2982 4521 3178 4522
rect 2982 4495 3151 4521
rect 3177 4495 3178 4521
rect 2982 4494 3178 4495
rect 1432 4326 1564 4331
rect 1460 4298 1484 4326
rect 1512 4298 1536 4326
rect 1432 4293 1564 4298
rect 1638 4186 1666 4191
rect 1638 4185 1722 4186
rect 1638 4159 1639 4185
rect 1665 4159 1722 4185
rect 1638 4158 1722 4159
rect 1638 4153 1666 4158
rect 1694 4130 1722 4158
rect 1694 4097 1722 4102
rect 2926 4130 2954 4135
rect 2982 4130 3010 4494
rect 3150 4489 3178 4494
rect 3318 4522 3346 4527
rect 3318 4475 3346 4494
rect 3598 4522 3626 4527
rect 3262 4465 3290 4471
rect 3262 4439 3263 4465
rect 3289 4439 3290 4465
rect 3084 4326 3216 4331
rect 3112 4298 3136 4326
rect 3164 4298 3188 4326
rect 3084 4293 3216 4298
rect 3262 4298 3290 4439
rect 3262 4270 3346 4298
rect 2954 4102 3010 4130
rect 3038 4242 3066 4247
rect 2926 4083 2954 4102
rect 966 4073 994 4079
rect 966 4047 967 4073
rect 993 4047 994 4073
rect 966 4018 994 4047
rect 910 3850 938 3855
rect 966 3850 994 3990
rect 2982 4017 3010 4023
rect 2982 3991 2983 4017
rect 3009 3991 3010 4017
rect 2258 3934 2390 3939
rect 2286 3906 2310 3934
rect 2338 3906 2362 3934
rect 2258 3901 2390 3906
rect 910 3849 994 3850
rect 910 3823 911 3849
rect 937 3823 994 3849
rect 910 3822 994 3823
rect 2982 3850 3010 3991
rect 910 3817 938 3822
rect 2982 3817 3010 3822
rect 3038 3738 3066 4214
rect 2814 3737 3066 3738
rect 2814 3711 3039 3737
rect 3065 3711 3066 3737
rect 2814 3710 3066 3711
rect 1432 3542 1564 3547
rect 1460 3514 1484 3542
rect 1512 3514 1536 3542
rect 1432 3509 1564 3514
rect 2258 3150 2390 3155
rect 2286 3122 2310 3150
rect 2338 3122 2362 3150
rect 2258 3117 2390 3122
rect 2814 2954 2842 3710
rect 3038 3705 3066 3710
rect 3262 4185 3290 4191
rect 3262 4159 3263 4185
rect 3289 4159 3290 4185
rect 3262 3626 3290 4159
rect 3262 3593 3290 3598
rect 3084 3542 3216 3547
rect 3112 3514 3136 3542
rect 3164 3514 3188 3542
rect 3084 3509 3216 3514
rect 3318 3402 3346 4270
rect 3150 3374 3346 3402
rect 3374 3681 3402 3687
rect 3374 3655 3375 3681
rect 3401 3655 3402 3681
rect 3150 3009 3178 3374
rect 3150 2983 3151 3009
rect 3177 2983 3178 3009
rect 3150 2977 3178 2983
rect 2534 2953 2842 2954
rect 2534 2927 2815 2953
rect 2841 2927 2842 2953
rect 2534 2926 2842 2927
rect 1432 2758 1564 2763
rect 1460 2730 1484 2758
rect 1512 2730 1536 2758
rect 1432 2725 1564 2730
rect 2258 2366 2390 2371
rect 2286 2338 2310 2366
rect 2338 2338 2362 2366
rect 2258 2333 2390 2338
rect 1432 1974 1564 1979
rect 1460 1946 1484 1974
rect 1512 1946 1536 1974
rect 1432 1941 1564 1946
rect 2478 1834 2506 1839
rect 2534 1834 2562 2926
rect 2814 2921 2842 2926
rect 3374 2898 3402 3655
rect 3598 3401 3626 4494
rect 3654 4521 3682 4527
rect 3654 4495 3655 4521
rect 3681 4495 3682 4521
rect 3654 4242 3682 4495
rect 3654 4209 3682 4214
rect 3710 4521 3738 4527
rect 3710 4495 3711 4521
rect 3737 4495 3738 4521
rect 3710 3682 3738 4495
rect 3822 4521 3850 4527
rect 3822 4495 3823 4521
rect 3849 4495 3850 4521
rect 3766 4466 3794 4471
rect 3766 4419 3794 4438
rect 3822 4242 3850 4495
rect 3878 4522 3906 4527
rect 3878 4475 3906 4494
rect 4214 4466 4242 4471
rect 4214 4419 4242 4438
rect 4736 4326 4868 4331
rect 4764 4298 4788 4326
rect 4816 4298 4840 4326
rect 4736 4293 4868 4298
rect 6388 4326 6520 4331
rect 6416 4298 6440 4326
rect 6468 4298 6492 4326
rect 6388 4293 6520 4298
rect 3822 4209 3850 4214
rect 4718 4130 4746 4135
rect 4718 4083 4746 4102
rect 5054 4130 5082 4135
rect 4326 4074 4354 4079
rect 4326 4073 4634 4074
rect 4326 4047 4327 4073
rect 4353 4047 4634 4073
rect 4326 4046 4634 4047
rect 4326 4041 4354 4046
rect 3910 3934 4042 3939
rect 3938 3906 3962 3934
rect 3990 3906 4014 3934
rect 3910 3901 4042 3906
rect 4606 3906 4634 4046
rect 4606 3878 4970 3906
rect 4942 3849 4970 3878
rect 4942 3823 4943 3849
rect 4969 3823 4970 3849
rect 4942 3817 4970 3823
rect 4998 3850 5026 3855
rect 4998 3803 5026 3822
rect 3710 3649 3738 3654
rect 4438 3682 4466 3687
rect 4438 3635 4466 3654
rect 4886 3682 4914 3687
rect 4886 3635 4914 3654
rect 3598 3375 3599 3401
rect 3625 3375 3626 3401
rect 3598 3369 3626 3375
rect 4662 3626 4690 3631
rect 4662 3345 4690 3598
rect 4736 3542 4868 3547
rect 4764 3514 4788 3542
rect 4816 3514 4840 3542
rect 4736 3509 4868 3514
rect 4662 3319 4663 3345
rect 4689 3319 4690 3345
rect 4662 3313 4690 3319
rect 5054 3402 5082 4102
rect 5562 3934 5694 3939
rect 5590 3906 5614 3934
rect 5642 3906 5666 3934
rect 5562 3901 5694 3906
rect 7214 3934 7346 3939
rect 7242 3906 7266 3934
rect 7294 3906 7318 3934
rect 7214 3901 7346 3906
rect 6388 3542 6520 3547
rect 6416 3514 6440 3542
rect 6468 3514 6492 3542
rect 6388 3509 6520 3514
rect 5054 3345 5082 3374
rect 5054 3319 5055 3345
rect 5081 3319 5082 3345
rect 5054 3313 5082 3319
rect 5446 3402 5474 3407
rect 3910 3150 4042 3155
rect 3938 3122 3962 3150
rect 3990 3122 4014 3150
rect 3910 3117 4042 3122
rect 3374 2865 3402 2870
rect 4214 2898 4242 2903
rect 4214 2851 4242 2870
rect 3084 2758 3216 2763
rect 3112 2730 3136 2758
rect 3164 2730 3188 2758
rect 3084 2725 3216 2730
rect 4736 2758 4868 2763
rect 4764 2730 4788 2758
rect 4816 2730 4840 2758
rect 4736 2725 4868 2730
rect 3910 2366 4042 2371
rect 3938 2338 3962 2366
rect 3990 2338 4014 2366
rect 3910 2333 4042 2338
rect 3084 1974 3216 1979
rect 3112 1946 3136 1974
rect 3164 1946 3188 1974
rect 3084 1941 3216 1946
rect 4736 1974 4868 1979
rect 4764 1946 4788 1974
rect 4816 1946 4840 1974
rect 4736 1941 4868 1946
rect 2478 1833 2562 1834
rect 2478 1807 2479 1833
rect 2505 1807 2562 1833
rect 2478 1806 2562 1807
rect 5446 1833 5474 3374
rect 5562 3150 5694 3155
rect 5590 3122 5614 3150
rect 5642 3122 5666 3150
rect 5562 3117 5694 3122
rect 7214 3150 7346 3155
rect 7242 3122 7266 3150
rect 7294 3122 7318 3150
rect 7214 3117 7346 3122
rect 6388 2758 6520 2763
rect 6416 2730 6440 2758
rect 6468 2730 6492 2758
rect 6388 2725 6520 2730
rect 5562 2366 5694 2371
rect 5590 2338 5614 2366
rect 5642 2338 5666 2366
rect 5562 2333 5694 2338
rect 7214 2366 7346 2371
rect 7242 2338 7266 2366
rect 7294 2338 7318 2366
rect 7214 2333 7346 2338
rect 6388 1974 6520 1979
rect 6416 1946 6440 1974
rect 6468 1946 6492 1974
rect 6388 1941 6520 1946
rect 5446 1807 5447 1833
rect 5473 1807 5474 1833
rect 2478 1801 2506 1806
rect 5446 1801 5474 1807
rect 1974 1722 2002 1727
rect 1974 400 2002 1694
rect 2814 1722 2842 1727
rect 2814 1675 2842 1694
rect 5950 1722 5978 1727
rect 2258 1582 2390 1587
rect 2286 1554 2310 1582
rect 2338 1554 2362 1582
rect 2258 1549 2390 1554
rect 3910 1582 4042 1587
rect 3938 1554 3962 1582
rect 3990 1554 4014 1582
rect 3910 1549 4042 1554
rect 5562 1582 5694 1587
rect 5590 1554 5614 1582
rect 5642 1554 5666 1582
rect 5562 1549 5694 1554
rect 5950 400 5978 1694
rect 6398 1722 6426 1727
rect 6398 1675 6426 1694
rect 7214 1582 7346 1587
rect 7242 1554 7266 1582
rect 7294 1554 7318 1582
rect 7214 1549 7346 1554
rect 1960 0 2016 400
rect 5936 0 5992 400
<< via2 >>
rect 2258 6285 2286 6286
rect 2258 6259 2259 6285
rect 2259 6259 2285 6285
rect 2285 6259 2286 6285
rect 2258 6258 2286 6259
rect 2310 6285 2338 6286
rect 2310 6259 2311 6285
rect 2311 6259 2337 6285
rect 2337 6259 2338 6285
rect 2310 6258 2338 6259
rect 2362 6285 2390 6286
rect 2362 6259 2363 6285
rect 2363 6259 2389 6285
rect 2389 6259 2390 6285
rect 2362 6258 2390 6259
rect 3910 6285 3938 6286
rect 3910 6259 3911 6285
rect 3911 6259 3937 6285
rect 3937 6259 3938 6285
rect 3910 6258 3938 6259
rect 3962 6285 3990 6286
rect 3962 6259 3963 6285
rect 3963 6259 3989 6285
rect 3989 6259 3990 6285
rect 3962 6258 3990 6259
rect 4014 6285 4042 6286
rect 4014 6259 4015 6285
rect 4015 6259 4041 6285
rect 4041 6259 4042 6285
rect 4014 6258 4042 6259
rect 5562 6285 5590 6286
rect 5562 6259 5563 6285
rect 5563 6259 5589 6285
rect 5589 6259 5590 6285
rect 5562 6258 5590 6259
rect 5614 6285 5642 6286
rect 5614 6259 5615 6285
rect 5615 6259 5641 6285
rect 5641 6259 5642 6285
rect 5614 6258 5642 6259
rect 5666 6285 5694 6286
rect 5666 6259 5667 6285
rect 5667 6259 5693 6285
rect 5693 6259 5694 6285
rect 5666 6258 5694 6259
rect 7214 6285 7242 6286
rect 7214 6259 7215 6285
rect 7215 6259 7241 6285
rect 7241 6259 7242 6285
rect 7214 6258 7242 6259
rect 7266 6285 7294 6286
rect 7266 6259 7267 6285
rect 7267 6259 7293 6285
rect 7293 6259 7294 6285
rect 7266 6258 7294 6259
rect 7318 6285 7346 6286
rect 7318 6259 7319 6285
rect 7319 6259 7345 6285
rect 7345 6259 7346 6285
rect 7318 6258 7346 6259
rect 1432 5893 1460 5894
rect 1432 5867 1433 5893
rect 1433 5867 1459 5893
rect 1459 5867 1460 5893
rect 1432 5866 1460 5867
rect 1484 5893 1512 5894
rect 1484 5867 1485 5893
rect 1485 5867 1511 5893
rect 1511 5867 1512 5893
rect 1484 5866 1512 5867
rect 1536 5893 1564 5894
rect 1536 5867 1537 5893
rect 1537 5867 1563 5893
rect 1563 5867 1564 5893
rect 1536 5866 1564 5867
rect 3084 5893 3112 5894
rect 3084 5867 3085 5893
rect 3085 5867 3111 5893
rect 3111 5867 3112 5893
rect 3084 5866 3112 5867
rect 3136 5893 3164 5894
rect 3136 5867 3137 5893
rect 3137 5867 3163 5893
rect 3163 5867 3164 5893
rect 3136 5866 3164 5867
rect 3188 5893 3216 5894
rect 3188 5867 3189 5893
rect 3189 5867 3215 5893
rect 3215 5867 3216 5893
rect 3188 5866 3216 5867
rect 4736 5893 4764 5894
rect 4736 5867 4737 5893
rect 4737 5867 4763 5893
rect 4763 5867 4764 5893
rect 4736 5866 4764 5867
rect 4788 5893 4816 5894
rect 4788 5867 4789 5893
rect 4789 5867 4815 5893
rect 4815 5867 4816 5893
rect 4788 5866 4816 5867
rect 4840 5893 4868 5894
rect 4840 5867 4841 5893
rect 4841 5867 4867 5893
rect 4867 5867 4868 5893
rect 4840 5866 4868 5867
rect 2258 5501 2286 5502
rect 2258 5475 2259 5501
rect 2259 5475 2285 5501
rect 2285 5475 2286 5501
rect 2258 5474 2286 5475
rect 2310 5501 2338 5502
rect 2310 5475 2311 5501
rect 2311 5475 2337 5501
rect 2337 5475 2338 5501
rect 2310 5474 2338 5475
rect 2362 5501 2390 5502
rect 2362 5475 2363 5501
rect 2363 5475 2389 5501
rect 2389 5475 2390 5501
rect 2362 5474 2390 5475
rect 3910 5501 3938 5502
rect 3910 5475 3911 5501
rect 3911 5475 3937 5501
rect 3937 5475 3938 5501
rect 3910 5474 3938 5475
rect 3962 5501 3990 5502
rect 3962 5475 3963 5501
rect 3963 5475 3989 5501
rect 3989 5475 3990 5501
rect 3962 5474 3990 5475
rect 4014 5501 4042 5502
rect 4014 5475 4015 5501
rect 4015 5475 4041 5501
rect 4041 5475 4042 5501
rect 4014 5474 4042 5475
rect 1432 5109 1460 5110
rect 1432 5083 1433 5109
rect 1433 5083 1459 5109
rect 1459 5083 1460 5109
rect 1432 5082 1460 5083
rect 1484 5109 1512 5110
rect 1484 5083 1485 5109
rect 1485 5083 1511 5109
rect 1511 5083 1512 5109
rect 1484 5082 1512 5083
rect 1536 5109 1564 5110
rect 1536 5083 1537 5109
rect 1537 5083 1563 5109
rect 1563 5083 1564 5109
rect 1536 5082 1564 5083
rect 3084 5109 3112 5110
rect 3084 5083 3085 5109
rect 3085 5083 3111 5109
rect 3111 5083 3112 5109
rect 3084 5082 3112 5083
rect 3136 5109 3164 5110
rect 3136 5083 3137 5109
rect 3137 5083 3163 5109
rect 3163 5083 3164 5109
rect 3136 5082 3164 5083
rect 3188 5109 3216 5110
rect 3188 5083 3189 5109
rect 3189 5083 3215 5109
rect 3215 5083 3216 5109
rect 3188 5082 3216 5083
rect 2258 4717 2286 4718
rect 2258 4691 2259 4717
rect 2259 4691 2285 4717
rect 2285 4691 2286 4717
rect 2258 4690 2286 4691
rect 2310 4717 2338 4718
rect 2310 4691 2311 4717
rect 2311 4691 2337 4717
rect 2337 4691 2338 4717
rect 2310 4690 2338 4691
rect 2362 4717 2390 4718
rect 2362 4691 2363 4717
rect 2363 4691 2389 4717
rect 2389 4691 2390 4717
rect 2362 4690 2390 4691
rect 3910 4717 3938 4718
rect 3910 4691 3911 4717
rect 3911 4691 3937 4717
rect 3937 4691 3938 4717
rect 3910 4690 3938 4691
rect 3962 4717 3990 4718
rect 3962 4691 3963 4717
rect 3963 4691 3989 4717
rect 3989 4691 3990 4717
rect 3962 4690 3990 4691
rect 4014 4717 4042 4718
rect 4014 4691 4015 4717
rect 4015 4691 4041 4717
rect 4041 4691 4042 4717
rect 4014 4690 4042 4691
rect 6388 5893 6416 5894
rect 6388 5867 6389 5893
rect 6389 5867 6415 5893
rect 6415 5867 6416 5893
rect 6388 5866 6416 5867
rect 6440 5893 6468 5894
rect 6440 5867 6441 5893
rect 6441 5867 6467 5893
rect 6467 5867 6468 5893
rect 6440 5866 6468 5867
rect 6492 5893 6520 5894
rect 6492 5867 6493 5893
rect 6493 5867 6519 5893
rect 6519 5867 6520 5893
rect 6492 5866 6520 5867
rect 5562 5501 5590 5502
rect 5562 5475 5563 5501
rect 5563 5475 5589 5501
rect 5589 5475 5590 5501
rect 5562 5474 5590 5475
rect 5614 5501 5642 5502
rect 5614 5475 5615 5501
rect 5615 5475 5641 5501
rect 5641 5475 5642 5501
rect 5614 5474 5642 5475
rect 5666 5501 5694 5502
rect 5666 5475 5667 5501
rect 5667 5475 5693 5501
rect 5693 5475 5694 5501
rect 5666 5474 5694 5475
rect 7214 5501 7242 5502
rect 7214 5475 7215 5501
rect 7215 5475 7241 5501
rect 7241 5475 7242 5501
rect 7214 5474 7242 5475
rect 7266 5501 7294 5502
rect 7266 5475 7267 5501
rect 7267 5475 7293 5501
rect 7293 5475 7294 5501
rect 7266 5474 7294 5475
rect 7318 5501 7346 5502
rect 7318 5475 7319 5501
rect 7319 5475 7345 5501
rect 7345 5475 7346 5501
rect 7318 5474 7346 5475
rect 4736 5109 4764 5110
rect 4736 5083 4737 5109
rect 4737 5083 4763 5109
rect 4763 5083 4764 5109
rect 4736 5082 4764 5083
rect 4788 5109 4816 5110
rect 4788 5083 4789 5109
rect 4789 5083 4815 5109
rect 4815 5083 4816 5109
rect 4788 5082 4816 5083
rect 4840 5109 4868 5110
rect 4840 5083 4841 5109
rect 4841 5083 4867 5109
rect 4867 5083 4868 5109
rect 4840 5082 4868 5083
rect 6388 5109 6416 5110
rect 6388 5083 6389 5109
rect 6389 5083 6415 5109
rect 6415 5083 6416 5109
rect 6388 5082 6416 5083
rect 6440 5109 6468 5110
rect 6440 5083 6441 5109
rect 6441 5083 6467 5109
rect 6467 5083 6468 5109
rect 6440 5082 6468 5083
rect 6492 5109 6520 5110
rect 6492 5083 6493 5109
rect 6493 5083 6519 5109
rect 6519 5083 6520 5109
rect 6492 5082 6520 5083
rect 5562 4717 5590 4718
rect 5562 4691 5563 4717
rect 5563 4691 5589 4717
rect 5589 4691 5590 4717
rect 5562 4690 5590 4691
rect 5614 4717 5642 4718
rect 5614 4691 5615 4717
rect 5615 4691 5641 4717
rect 5641 4691 5642 4717
rect 5614 4690 5642 4691
rect 5666 4717 5694 4718
rect 5666 4691 5667 4717
rect 5667 4691 5693 4717
rect 5693 4691 5694 4717
rect 5666 4690 5694 4691
rect 7214 4717 7242 4718
rect 7214 4691 7215 4717
rect 7215 4691 7241 4717
rect 7241 4691 7242 4717
rect 7214 4690 7242 4691
rect 7266 4717 7294 4718
rect 7266 4691 7267 4717
rect 7267 4691 7293 4717
rect 7293 4691 7294 4717
rect 7266 4690 7294 4691
rect 7318 4717 7346 4718
rect 7318 4691 7319 4717
rect 7319 4691 7345 4717
rect 7345 4691 7346 4717
rect 7318 4690 7346 4691
rect 1432 4325 1460 4326
rect 1432 4299 1433 4325
rect 1433 4299 1459 4325
rect 1459 4299 1460 4325
rect 1432 4298 1460 4299
rect 1484 4325 1512 4326
rect 1484 4299 1485 4325
rect 1485 4299 1511 4325
rect 1511 4299 1512 4325
rect 1484 4298 1512 4299
rect 1536 4325 1564 4326
rect 1536 4299 1537 4325
rect 1537 4299 1563 4325
rect 1563 4299 1564 4325
rect 1536 4298 1564 4299
rect 1694 4102 1722 4130
rect 3318 4521 3346 4522
rect 3318 4495 3319 4521
rect 3319 4495 3345 4521
rect 3345 4495 3346 4521
rect 3318 4494 3346 4495
rect 3598 4494 3626 4522
rect 3084 4325 3112 4326
rect 3084 4299 3085 4325
rect 3085 4299 3111 4325
rect 3111 4299 3112 4325
rect 3084 4298 3112 4299
rect 3136 4325 3164 4326
rect 3136 4299 3137 4325
rect 3137 4299 3163 4325
rect 3163 4299 3164 4325
rect 3136 4298 3164 4299
rect 3188 4325 3216 4326
rect 3188 4299 3189 4325
rect 3189 4299 3215 4325
rect 3215 4299 3216 4325
rect 3188 4298 3216 4299
rect 2926 4129 2954 4130
rect 2926 4103 2927 4129
rect 2927 4103 2953 4129
rect 2953 4103 2954 4129
rect 2926 4102 2954 4103
rect 3038 4214 3066 4242
rect 966 3990 994 4018
rect 2258 3933 2286 3934
rect 2258 3907 2259 3933
rect 2259 3907 2285 3933
rect 2285 3907 2286 3933
rect 2258 3906 2286 3907
rect 2310 3933 2338 3934
rect 2310 3907 2311 3933
rect 2311 3907 2337 3933
rect 2337 3907 2338 3933
rect 2310 3906 2338 3907
rect 2362 3933 2390 3934
rect 2362 3907 2363 3933
rect 2363 3907 2389 3933
rect 2389 3907 2390 3933
rect 2362 3906 2390 3907
rect 2982 3822 3010 3850
rect 1432 3541 1460 3542
rect 1432 3515 1433 3541
rect 1433 3515 1459 3541
rect 1459 3515 1460 3541
rect 1432 3514 1460 3515
rect 1484 3541 1512 3542
rect 1484 3515 1485 3541
rect 1485 3515 1511 3541
rect 1511 3515 1512 3541
rect 1484 3514 1512 3515
rect 1536 3541 1564 3542
rect 1536 3515 1537 3541
rect 1537 3515 1563 3541
rect 1563 3515 1564 3541
rect 1536 3514 1564 3515
rect 2258 3149 2286 3150
rect 2258 3123 2259 3149
rect 2259 3123 2285 3149
rect 2285 3123 2286 3149
rect 2258 3122 2286 3123
rect 2310 3149 2338 3150
rect 2310 3123 2311 3149
rect 2311 3123 2337 3149
rect 2337 3123 2338 3149
rect 2310 3122 2338 3123
rect 2362 3149 2390 3150
rect 2362 3123 2363 3149
rect 2363 3123 2389 3149
rect 2389 3123 2390 3149
rect 2362 3122 2390 3123
rect 3262 3598 3290 3626
rect 3084 3541 3112 3542
rect 3084 3515 3085 3541
rect 3085 3515 3111 3541
rect 3111 3515 3112 3541
rect 3084 3514 3112 3515
rect 3136 3541 3164 3542
rect 3136 3515 3137 3541
rect 3137 3515 3163 3541
rect 3163 3515 3164 3541
rect 3136 3514 3164 3515
rect 3188 3541 3216 3542
rect 3188 3515 3189 3541
rect 3189 3515 3215 3541
rect 3215 3515 3216 3541
rect 3188 3514 3216 3515
rect 1432 2757 1460 2758
rect 1432 2731 1433 2757
rect 1433 2731 1459 2757
rect 1459 2731 1460 2757
rect 1432 2730 1460 2731
rect 1484 2757 1512 2758
rect 1484 2731 1485 2757
rect 1485 2731 1511 2757
rect 1511 2731 1512 2757
rect 1484 2730 1512 2731
rect 1536 2757 1564 2758
rect 1536 2731 1537 2757
rect 1537 2731 1563 2757
rect 1563 2731 1564 2757
rect 1536 2730 1564 2731
rect 2258 2365 2286 2366
rect 2258 2339 2259 2365
rect 2259 2339 2285 2365
rect 2285 2339 2286 2365
rect 2258 2338 2286 2339
rect 2310 2365 2338 2366
rect 2310 2339 2311 2365
rect 2311 2339 2337 2365
rect 2337 2339 2338 2365
rect 2310 2338 2338 2339
rect 2362 2365 2390 2366
rect 2362 2339 2363 2365
rect 2363 2339 2389 2365
rect 2389 2339 2390 2365
rect 2362 2338 2390 2339
rect 1432 1973 1460 1974
rect 1432 1947 1433 1973
rect 1433 1947 1459 1973
rect 1459 1947 1460 1973
rect 1432 1946 1460 1947
rect 1484 1973 1512 1974
rect 1484 1947 1485 1973
rect 1485 1947 1511 1973
rect 1511 1947 1512 1973
rect 1484 1946 1512 1947
rect 1536 1973 1564 1974
rect 1536 1947 1537 1973
rect 1537 1947 1563 1973
rect 1563 1947 1564 1973
rect 1536 1946 1564 1947
rect 3654 4214 3682 4242
rect 3766 4465 3794 4466
rect 3766 4439 3767 4465
rect 3767 4439 3793 4465
rect 3793 4439 3794 4465
rect 3766 4438 3794 4439
rect 3878 4521 3906 4522
rect 3878 4495 3879 4521
rect 3879 4495 3905 4521
rect 3905 4495 3906 4521
rect 3878 4494 3906 4495
rect 4214 4465 4242 4466
rect 4214 4439 4215 4465
rect 4215 4439 4241 4465
rect 4241 4439 4242 4465
rect 4214 4438 4242 4439
rect 4736 4325 4764 4326
rect 4736 4299 4737 4325
rect 4737 4299 4763 4325
rect 4763 4299 4764 4325
rect 4736 4298 4764 4299
rect 4788 4325 4816 4326
rect 4788 4299 4789 4325
rect 4789 4299 4815 4325
rect 4815 4299 4816 4325
rect 4788 4298 4816 4299
rect 4840 4325 4868 4326
rect 4840 4299 4841 4325
rect 4841 4299 4867 4325
rect 4867 4299 4868 4325
rect 4840 4298 4868 4299
rect 6388 4325 6416 4326
rect 6388 4299 6389 4325
rect 6389 4299 6415 4325
rect 6415 4299 6416 4325
rect 6388 4298 6416 4299
rect 6440 4325 6468 4326
rect 6440 4299 6441 4325
rect 6441 4299 6467 4325
rect 6467 4299 6468 4325
rect 6440 4298 6468 4299
rect 6492 4325 6520 4326
rect 6492 4299 6493 4325
rect 6493 4299 6519 4325
rect 6519 4299 6520 4325
rect 6492 4298 6520 4299
rect 3822 4214 3850 4242
rect 4718 4129 4746 4130
rect 4718 4103 4719 4129
rect 4719 4103 4745 4129
rect 4745 4103 4746 4129
rect 4718 4102 4746 4103
rect 5054 4102 5082 4130
rect 3910 3933 3938 3934
rect 3910 3907 3911 3933
rect 3911 3907 3937 3933
rect 3937 3907 3938 3933
rect 3910 3906 3938 3907
rect 3962 3933 3990 3934
rect 3962 3907 3963 3933
rect 3963 3907 3989 3933
rect 3989 3907 3990 3933
rect 3962 3906 3990 3907
rect 4014 3933 4042 3934
rect 4014 3907 4015 3933
rect 4015 3907 4041 3933
rect 4041 3907 4042 3933
rect 4014 3906 4042 3907
rect 4998 3849 5026 3850
rect 4998 3823 4999 3849
rect 4999 3823 5025 3849
rect 5025 3823 5026 3849
rect 4998 3822 5026 3823
rect 3710 3654 3738 3682
rect 4438 3681 4466 3682
rect 4438 3655 4439 3681
rect 4439 3655 4465 3681
rect 4465 3655 4466 3681
rect 4438 3654 4466 3655
rect 4886 3681 4914 3682
rect 4886 3655 4887 3681
rect 4887 3655 4913 3681
rect 4913 3655 4914 3681
rect 4886 3654 4914 3655
rect 4662 3598 4690 3626
rect 4736 3541 4764 3542
rect 4736 3515 4737 3541
rect 4737 3515 4763 3541
rect 4763 3515 4764 3541
rect 4736 3514 4764 3515
rect 4788 3541 4816 3542
rect 4788 3515 4789 3541
rect 4789 3515 4815 3541
rect 4815 3515 4816 3541
rect 4788 3514 4816 3515
rect 4840 3541 4868 3542
rect 4840 3515 4841 3541
rect 4841 3515 4867 3541
rect 4867 3515 4868 3541
rect 4840 3514 4868 3515
rect 5562 3933 5590 3934
rect 5562 3907 5563 3933
rect 5563 3907 5589 3933
rect 5589 3907 5590 3933
rect 5562 3906 5590 3907
rect 5614 3933 5642 3934
rect 5614 3907 5615 3933
rect 5615 3907 5641 3933
rect 5641 3907 5642 3933
rect 5614 3906 5642 3907
rect 5666 3933 5694 3934
rect 5666 3907 5667 3933
rect 5667 3907 5693 3933
rect 5693 3907 5694 3933
rect 5666 3906 5694 3907
rect 7214 3933 7242 3934
rect 7214 3907 7215 3933
rect 7215 3907 7241 3933
rect 7241 3907 7242 3933
rect 7214 3906 7242 3907
rect 7266 3933 7294 3934
rect 7266 3907 7267 3933
rect 7267 3907 7293 3933
rect 7293 3907 7294 3933
rect 7266 3906 7294 3907
rect 7318 3933 7346 3934
rect 7318 3907 7319 3933
rect 7319 3907 7345 3933
rect 7345 3907 7346 3933
rect 7318 3906 7346 3907
rect 6388 3541 6416 3542
rect 6388 3515 6389 3541
rect 6389 3515 6415 3541
rect 6415 3515 6416 3541
rect 6388 3514 6416 3515
rect 6440 3541 6468 3542
rect 6440 3515 6441 3541
rect 6441 3515 6467 3541
rect 6467 3515 6468 3541
rect 6440 3514 6468 3515
rect 6492 3541 6520 3542
rect 6492 3515 6493 3541
rect 6493 3515 6519 3541
rect 6519 3515 6520 3541
rect 6492 3514 6520 3515
rect 5054 3374 5082 3402
rect 5446 3374 5474 3402
rect 3910 3149 3938 3150
rect 3910 3123 3911 3149
rect 3911 3123 3937 3149
rect 3937 3123 3938 3149
rect 3910 3122 3938 3123
rect 3962 3149 3990 3150
rect 3962 3123 3963 3149
rect 3963 3123 3989 3149
rect 3989 3123 3990 3149
rect 3962 3122 3990 3123
rect 4014 3149 4042 3150
rect 4014 3123 4015 3149
rect 4015 3123 4041 3149
rect 4041 3123 4042 3149
rect 4014 3122 4042 3123
rect 3374 2870 3402 2898
rect 4214 2897 4242 2898
rect 4214 2871 4215 2897
rect 4215 2871 4241 2897
rect 4241 2871 4242 2897
rect 4214 2870 4242 2871
rect 3084 2757 3112 2758
rect 3084 2731 3085 2757
rect 3085 2731 3111 2757
rect 3111 2731 3112 2757
rect 3084 2730 3112 2731
rect 3136 2757 3164 2758
rect 3136 2731 3137 2757
rect 3137 2731 3163 2757
rect 3163 2731 3164 2757
rect 3136 2730 3164 2731
rect 3188 2757 3216 2758
rect 3188 2731 3189 2757
rect 3189 2731 3215 2757
rect 3215 2731 3216 2757
rect 3188 2730 3216 2731
rect 4736 2757 4764 2758
rect 4736 2731 4737 2757
rect 4737 2731 4763 2757
rect 4763 2731 4764 2757
rect 4736 2730 4764 2731
rect 4788 2757 4816 2758
rect 4788 2731 4789 2757
rect 4789 2731 4815 2757
rect 4815 2731 4816 2757
rect 4788 2730 4816 2731
rect 4840 2757 4868 2758
rect 4840 2731 4841 2757
rect 4841 2731 4867 2757
rect 4867 2731 4868 2757
rect 4840 2730 4868 2731
rect 3910 2365 3938 2366
rect 3910 2339 3911 2365
rect 3911 2339 3937 2365
rect 3937 2339 3938 2365
rect 3910 2338 3938 2339
rect 3962 2365 3990 2366
rect 3962 2339 3963 2365
rect 3963 2339 3989 2365
rect 3989 2339 3990 2365
rect 3962 2338 3990 2339
rect 4014 2365 4042 2366
rect 4014 2339 4015 2365
rect 4015 2339 4041 2365
rect 4041 2339 4042 2365
rect 4014 2338 4042 2339
rect 3084 1973 3112 1974
rect 3084 1947 3085 1973
rect 3085 1947 3111 1973
rect 3111 1947 3112 1973
rect 3084 1946 3112 1947
rect 3136 1973 3164 1974
rect 3136 1947 3137 1973
rect 3137 1947 3163 1973
rect 3163 1947 3164 1973
rect 3136 1946 3164 1947
rect 3188 1973 3216 1974
rect 3188 1947 3189 1973
rect 3189 1947 3215 1973
rect 3215 1947 3216 1973
rect 3188 1946 3216 1947
rect 4736 1973 4764 1974
rect 4736 1947 4737 1973
rect 4737 1947 4763 1973
rect 4763 1947 4764 1973
rect 4736 1946 4764 1947
rect 4788 1973 4816 1974
rect 4788 1947 4789 1973
rect 4789 1947 4815 1973
rect 4815 1947 4816 1973
rect 4788 1946 4816 1947
rect 4840 1973 4868 1974
rect 4840 1947 4841 1973
rect 4841 1947 4867 1973
rect 4867 1947 4868 1973
rect 4840 1946 4868 1947
rect 5562 3149 5590 3150
rect 5562 3123 5563 3149
rect 5563 3123 5589 3149
rect 5589 3123 5590 3149
rect 5562 3122 5590 3123
rect 5614 3149 5642 3150
rect 5614 3123 5615 3149
rect 5615 3123 5641 3149
rect 5641 3123 5642 3149
rect 5614 3122 5642 3123
rect 5666 3149 5694 3150
rect 5666 3123 5667 3149
rect 5667 3123 5693 3149
rect 5693 3123 5694 3149
rect 5666 3122 5694 3123
rect 7214 3149 7242 3150
rect 7214 3123 7215 3149
rect 7215 3123 7241 3149
rect 7241 3123 7242 3149
rect 7214 3122 7242 3123
rect 7266 3149 7294 3150
rect 7266 3123 7267 3149
rect 7267 3123 7293 3149
rect 7293 3123 7294 3149
rect 7266 3122 7294 3123
rect 7318 3149 7346 3150
rect 7318 3123 7319 3149
rect 7319 3123 7345 3149
rect 7345 3123 7346 3149
rect 7318 3122 7346 3123
rect 6388 2757 6416 2758
rect 6388 2731 6389 2757
rect 6389 2731 6415 2757
rect 6415 2731 6416 2757
rect 6388 2730 6416 2731
rect 6440 2757 6468 2758
rect 6440 2731 6441 2757
rect 6441 2731 6467 2757
rect 6467 2731 6468 2757
rect 6440 2730 6468 2731
rect 6492 2757 6520 2758
rect 6492 2731 6493 2757
rect 6493 2731 6519 2757
rect 6519 2731 6520 2757
rect 6492 2730 6520 2731
rect 5562 2365 5590 2366
rect 5562 2339 5563 2365
rect 5563 2339 5589 2365
rect 5589 2339 5590 2365
rect 5562 2338 5590 2339
rect 5614 2365 5642 2366
rect 5614 2339 5615 2365
rect 5615 2339 5641 2365
rect 5641 2339 5642 2365
rect 5614 2338 5642 2339
rect 5666 2365 5694 2366
rect 5666 2339 5667 2365
rect 5667 2339 5693 2365
rect 5693 2339 5694 2365
rect 5666 2338 5694 2339
rect 7214 2365 7242 2366
rect 7214 2339 7215 2365
rect 7215 2339 7241 2365
rect 7241 2339 7242 2365
rect 7214 2338 7242 2339
rect 7266 2365 7294 2366
rect 7266 2339 7267 2365
rect 7267 2339 7293 2365
rect 7293 2339 7294 2365
rect 7266 2338 7294 2339
rect 7318 2365 7346 2366
rect 7318 2339 7319 2365
rect 7319 2339 7345 2365
rect 7345 2339 7346 2365
rect 7318 2338 7346 2339
rect 6388 1973 6416 1974
rect 6388 1947 6389 1973
rect 6389 1947 6415 1973
rect 6415 1947 6416 1973
rect 6388 1946 6416 1947
rect 6440 1973 6468 1974
rect 6440 1947 6441 1973
rect 6441 1947 6467 1973
rect 6467 1947 6468 1973
rect 6440 1946 6468 1947
rect 6492 1973 6520 1974
rect 6492 1947 6493 1973
rect 6493 1947 6519 1973
rect 6519 1947 6520 1973
rect 6492 1946 6520 1947
rect 1974 1721 2002 1722
rect 1974 1695 1975 1721
rect 1975 1695 2001 1721
rect 2001 1695 2002 1721
rect 1974 1694 2002 1695
rect 2814 1721 2842 1722
rect 2814 1695 2815 1721
rect 2815 1695 2841 1721
rect 2841 1695 2842 1721
rect 2814 1694 2842 1695
rect 5950 1721 5978 1722
rect 5950 1695 5951 1721
rect 5951 1695 5977 1721
rect 5977 1695 5978 1721
rect 5950 1694 5978 1695
rect 2258 1581 2286 1582
rect 2258 1555 2259 1581
rect 2259 1555 2285 1581
rect 2285 1555 2286 1581
rect 2258 1554 2286 1555
rect 2310 1581 2338 1582
rect 2310 1555 2311 1581
rect 2311 1555 2337 1581
rect 2337 1555 2338 1581
rect 2310 1554 2338 1555
rect 2362 1581 2390 1582
rect 2362 1555 2363 1581
rect 2363 1555 2389 1581
rect 2389 1555 2390 1581
rect 2362 1554 2390 1555
rect 3910 1581 3938 1582
rect 3910 1555 3911 1581
rect 3911 1555 3937 1581
rect 3937 1555 3938 1581
rect 3910 1554 3938 1555
rect 3962 1581 3990 1582
rect 3962 1555 3963 1581
rect 3963 1555 3989 1581
rect 3989 1555 3990 1581
rect 3962 1554 3990 1555
rect 4014 1581 4042 1582
rect 4014 1555 4015 1581
rect 4015 1555 4041 1581
rect 4041 1555 4042 1581
rect 4014 1554 4042 1555
rect 5562 1581 5590 1582
rect 5562 1555 5563 1581
rect 5563 1555 5589 1581
rect 5589 1555 5590 1581
rect 5562 1554 5590 1555
rect 5614 1581 5642 1582
rect 5614 1555 5615 1581
rect 5615 1555 5641 1581
rect 5641 1555 5642 1581
rect 5614 1554 5642 1555
rect 5666 1581 5694 1582
rect 5666 1555 5667 1581
rect 5667 1555 5693 1581
rect 5693 1555 5694 1581
rect 5666 1554 5694 1555
rect 6398 1721 6426 1722
rect 6398 1695 6399 1721
rect 6399 1695 6425 1721
rect 6425 1695 6426 1721
rect 6398 1694 6426 1695
rect 7214 1581 7242 1582
rect 7214 1555 7215 1581
rect 7215 1555 7241 1581
rect 7241 1555 7242 1581
rect 7214 1554 7242 1555
rect 7266 1581 7294 1582
rect 7266 1555 7267 1581
rect 7267 1555 7293 1581
rect 7293 1555 7294 1581
rect 7266 1554 7294 1555
rect 7318 1581 7346 1582
rect 7318 1555 7319 1581
rect 7319 1555 7345 1581
rect 7345 1555 7346 1581
rect 7318 1554 7346 1555
<< metal3 >>
rect 2253 6258 2258 6286
rect 2286 6258 2310 6286
rect 2338 6258 2362 6286
rect 2390 6258 2395 6286
rect 3905 6258 3910 6286
rect 3938 6258 3962 6286
rect 3990 6258 4014 6286
rect 4042 6258 4047 6286
rect 5557 6258 5562 6286
rect 5590 6258 5614 6286
rect 5642 6258 5666 6286
rect 5694 6258 5699 6286
rect 7209 6258 7214 6286
rect 7242 6258 7266 6286
rect 7294 6258 7318 6286
rect 7346 6258 7351 6286
rect 1427 5866 1432 5894
rect 1460 5866 1484 5894
rect 1512 5866 1536 5894
rect 1564 5866 1569 5894
rect 3079 5866 3084 5894
rect 3112 5866 3136 5894
rect 3164 5866 3188 5894
rect 3216 5866 3221 5894
rect 4731 5866 4736 5894
rect 4764 5866 4788 5894
rect 4816 5866 4840 5894
rect 4868 5866 4873 5894
rect 6383 5866 6388 5894
rect 6416 5866 6440 5894
rect 6468 5866 6492 5894
rect 6520 5866 6525 5894
rect 2253 5474 2258 5502
rect 2286 5474 2310 5502
rect 2338 5474 2362 5502
rect 2390 5474 2395 5502
rect 3905 5474 3910 5502
rect 3938 5474 3962 5502
rect 3990 5474 4014 5502
rect 4042 5474 4047 5502
rect 5557 5474 5562 5502
rect 5590 5474 5614 5502
rect 5642 5474 5666 5502
rect 5694 5474 5699 5502
rect 7209 5474 7214 5502
rect 7242 5474 7266 5502
rect 7294 5474 7318 5502
rect 7346 5474 7351 5502
rect 1427 5082 1432 5110
rect 1460 5082 1484 5110
rect 1512 5082 1536 5110
rect 1564 5082 1569 5110
rect 3079 5082 3084 5110
rect 3112 5082 3136 5110
rect 3164 5082 3188 5110
rect 3216 5082 3221 5110
rect 4731 5082 4736 5110
rect 4764 5082 4788 5110
rect 4816 5082 4840 5110
rect 4868 5082 4873 5110
rect 6383 5082 6388 5110
rect 6416 5082 6440 5110
rect 6468 5082 6492 5110
rect 6520 5082 6525 5110
rect 2253 4690 2258 4718
rect 2286 4690 2310 4718
rect 2338 4690 2362 4718
rect 2390 4690 2395 4718
rect 3905 4690 3910 4718
rect 3938 4690 3962 4718
rect 3990 4690 4014 4718
rect 4042 4690 4047 4718
rect 5557 4690 5562 4718
rect 5590 4690 5614 4718
rect 5642 4690 5666 4718
rect 5694 4690 5699 4718
rect 7209 4690 7214 4718
rect 7242 4690 7266 4718
rect 7294 4690 7318 4718
rect 7346 4690 7351 4718
rect 3313 4494 3318 4522
rect 3346 4494 3598 4522
rect 3626 4494 3878 4522
rect 3906 4494 3911 4522
rect 3761 4438 3766 4466
rect 3794 4438 4214 4466
rect 4242 4438 4247 4466
rect 1427 4298 1432 4326
rect 1460 4298 1484 4326
rect 1512 4298 1536 4326
rect 1564 4298 1569 4326
rect 3079 4298 3084 4326
rect 3112 4298 3136 4326
rect 3164 4298 3188 4326
rect 3216 4298 3221 4326
rect 4731 4298 4736 4326
rect 4764 4298 4788 4326
rect 4816 4298 4840 4326
rect 4868 4298 4873 4326
rect 6383 4298 6388 4326
rect 6416 4298 6440 4326
rect 6468 4298 6492 4326
rect 6520 4298 6525 4326
rect 3033 4214 3038 4242
rect 3066 4214 3654 4242
rect 3682 4214 3687 4242
rect 3817 4214 3822 4242
rect 3850 4214 4746 4242
rect 4718 4130 4746 4214
rect 1689 4102 1694 4130
rect 1722 4102 2926 4130
rect 2954 4102 2959 4130
rect 4713 4102 4718 4130
rect 4746 4102 5054 4130
rect 5082 4102 5087 4130
rect 0 4018 400 4032
rect 0 3990 966 4018
rect 994 3990 999 4018
rect 0 3976 400 3990
rect 2253 3906 2258 3934
rect 2286 3906 2310 3934
rect 2338 3906 2362 3934
rect 2390 3906 2395 3934
rect 3905 3906 3910 3934
rect 3938 3906 3962 3934
rect 3990 3906 4014 3934
rect 4042 3906 4047 3934
rect 5557 3906 5562 3934
rect 5590 3906 5614 3934
rect 5642 3906 5666 3934
rect 5694 3906 5699 3934
rect 7209 3906 7214 3934
rect 7242 3906 7266 3934
rect 7294 3906 7318 3934
rect 7346 3906 7351 3934
rect 2977 3822 2982 3850
rect 3010 3822 4998 3850
rect 5026 3822 5031 3850
rect 3705 3654 3710 3682
rect 3738 3654 4438 3682
rect 4466 3654 4886 3682
rect 4914 3654 4919 3682
rect 3257 3598 3262 3626
rect 3290 3598 4662 3626
rect 4690 3598 4695 3626
rect 1427 3514 1432 3542
rect 1460 3514 1484 3542
rect 1512 3514 1536 3542
rect 1564 3514 1569 3542
rect 3079 3514 3084 3542
rect 3112 3514 3136 3542
rect 3164 3514 3188 3542
rect 3216 3514 3221 3542
rect 4731 3514 4736 3542
rect 4764 3514 4788 3542
rect 4816 3514 4840 3542
rect 4868 3514 4873 3542
rect 6383 3514 6388 3542
rect 6416 3514 6440 3542
rect 6468 3514 6492 3542
rect 6520 3514 6525 3542
rect 5049 3374 5054 3402
rect 5082 3374 5446 3402
rect 5474 3374 5479 3402
rect 2253 3122 2258 3150
rect 2286 3122 2310 3150
rect 2338 3122 2362 3150
rect 2390 3122 2395 3150
rect 3905 3122 3910 3150
rect 3938 3122 3962 3150
rect 3990 3122 4014 3150
rect 4042 3122 4047 3150
rect 5557 3122 5562 3150
rect 5590 3122 5614 3150
rect 5642 3122 5666 3150
rect 5694 3122 5699 3150
rect 7209 3122 7214 3150
rect 7242 3122 7266 3150
rect 7294 3122 7318 3150
rect 7346 3122 7351 3150
rect 3369 2870 3374 2898
rect 3402 2870 4214 2898
rect 4242 2870 4247 2898
rect 1427 2730 1432 2758
rect 1460 2730 1484 2758
rect 1512 2730 1536 2758
rect 1564 2730 1569 2758
rect 3079 2730 3084 2758
rect 3112 2730 3136 2758
rect 3164 2730 3188 2758
rect 3216 2730 3221 2758
rect 4731 2730 4736 2758
rect 4764 2730 4788 2758
rect 4816 2730 4840 2758
rect 4868 2730 4873 2758
rect 6383 2730 6388 2758
rect 6416 2730 6440 2758
rect 6468 2730 6492 2758
rect 6520 2730 6525 2758
rect 2253 2338 2258 2366
rect 2286 2338 2310 2366
rect 2338 2338 2362 2366
rect 2390 2338 2395 2366
rect 3905 2338 3910 2366
rect 3938 2338 3962 2366
rect 3990 2338 4014 2366
rect 4042 2338 4047 2366
rect 5557 2338 5562 2366
rect 5590 2338 5614 2366
rect 5642 2338 5666 2366
rect 5694 2338 5699 2366
rect 7209 2338 7214 2366
rect 7242 2338 7266 2366
rect 7294 2338 7318 2366
rect 7346 2338 7351 2366
rect 1427 1946 1432 1974
rect 1460 1946 1484 1974
rect 1512 1946 1536 1974
rect 1564 1946 1569 1974
rect 3079 1946 3084 1974
rect 3112 1946 3136 1974
rect 3164 1946 3188 1974
rect 3216 1946 3221 1974
rect 4731 1946 4736 1974
rect 4764 1946 4788 1974
rect 4816 1946 4840 1974
rect 4868 1946 4873 1974
rect 6383 1946 6388 1974
rect 6416 1946 6440 1974
rect 6468 1946 6492 1974
rect 6520 1946 6525 1974
rect 1969 1694 1974 1722
rect 2002 1694 2814 1722
rect 2842 1694 2847 1722
rect 5945 1694 5950 1722
rect 5978 1694 6398 1722
rect 6426 1694 6431 1722
rect 2253 1554 2258 1582
rect 2286 1554 2310 1582
rect 2338 1554 2362 1582
rect 2390 1554 2395 1582
rect 3905 1554 3910 1582
rect 3938 1554 3962 1582
rect 3990 1554 4014 1582
rect 4042 1554 4047 1582
rect 5557 1554 5562 1582
rect 5590 1554 5614 1582
rect 5642 1554 5666 1582
rect 5694 1554 5699 1582
rect 7209 1554 7214 1582
rect 7242 1554 7266 1582
rect 7294 1554 7318 1582
rect 7346 1554 7351 1582
<< via3 >>
rect 2258 6258 2286 6286
rect 2310 6258 2338 6286
rect 2362 6258 2390 6286
rect 3910 6258 3938 6286
rect 3962 6258 3990 6286
rect 4014 6258 4042 6286
rect 5562 6258 5590 6286
rect 5614 6258 5642 6286
rect 5666 6258 5694 6286
rect 7214 6258 7242 6286
rect 7266 6258 7294 6286
rect 7318 6258 7346 6286
rect 1432 5866 1460 5894
rect 1484 5866 1512 5894
rect 1536 5866 1564 5894
rect 3084 5866 3112 5894
rect 3136 5866 3164 5894
rect 3188 5866 3216 5894
rect 4736 5866 4764 5894
rect 4788 5866 4816 5894
rect 4840 5866 4868 5894
rect 6388 5866 6416 5894
rect 6440 5866 6468 5894
rect 6492 5866 6520 5894
rect 2258 5474 2286 5502
rect 2310 5474 2338 5502
rect 2362 5474 2390 5502
rect 3910 5474 3938 5502
rect 3962 5474 3990 5502
rect 4014 5474 4042 5502
rect 5562 5474 5590 5502
rect 5614 5474 5642 5502
rect 5666 5474 5694 5502
rect 7214 5474 7242 5502
rect 7266 5474 7294 5502
rect 7318 5474 7346 5502
rect 1432 5082 1460 5110
rect 1484 5082 1512 5110
rect 1536 5082 1564 5110
rect 3084 5082 3112 5110
rect 3136 5082 3164 5110
rect 3188 5082 3216 5110
rect 4736 5082 4764 5110
rect 4788 5082 4816 5110
rect 4840 5082 4868 5110
rect 6388 5082 6416 5110
rect 6440 5082 6468 5110
rect 6492 5082 6520 5110
rect 2258 4690 2286 4718
rect 2310 4690 2338 4718
rect 2362 4690 2390 4718
rect 3910 4690 3938 4718
rect 3962 4690 3990 4718
rect 4014 4690 4042 4718
rect 5562 4690 5590 4718
rect 5614 4690 5642 4718
rect 5666 4690 5694 4718
rect 7214 4690 7242 4718
rect 7266 4690 7294 4718
rect 7318 4690 7346 4718
rect 1432 4298 1460 4326
rect 1484 4298 1512 4326
rect 1536 4298 1564 4326
rect 3084 4298 3112 4326
rect 3136 4298 3164 4326
rect 3188 4298 3216 4326
rect 4736 4298 4764 4326
rect 4788 4298 4816 4326
rect 4840 4298 4868 4326
rect 6388 4298 6416 4326
rect 6440 4298 6468 4326
rect 6492 4298 6520 4326
rect 2258 3906 2286 3934
rect 2310 3906 2338 3934
rect 2362 3906 2390 3934
rect 3910 3906 3938 3934
rect 3962 3906 3990 3934
rect 4014 3906 4042 3934
rect 5562 3906 5590 3934
rect 5614 3906 5642 3934
rect 5666 3906 5694 3934
rect 7214 3906 7242 3934
rect 7266 3906 7294 3934
rect 7318 3906 7346 3934
rect 1432 3514 1460 3542
rect 1484 3514 1512 3542
rect 1536 3514 1564 3542
rect 3084 3514 3112 3542
rect 3136 3514 3164 3542
rect 3188 3514 3216 3542
rect 4736 3514 4764 3542
rect 4788 3514 4816 3542
rect 4840 3514 4868 3542
rect 6388 3514 6416 3542
rect 6440 3514 6468 3542
rect 6492 3514 6520 3542
rect 2258 3122 2286 3150
rect 2310 3122 2338 3150
rect 2362 3122 2390 3150
rect 3910 3122 3938 3150
rect 3962 3122 3990 3150
rect 4014 3122 4042 3150
rect 5562 3122 5590 3150
rect 5614 3122 5642 3150
rect 5666 3122 5694 3150
rect 7214 3122 7242 3150
rect 7266 3122 7294 3150
rect 7318 3122 7346 3150
rect 1432 2730 1460 2758
rect 1484 2730 1512 2758
rect 1536 2730 1564 2758
rect 3084 2730 3112 2758
rect 3136 2730 3164 2758
rect 3188 2730 3216 2758
rect 4736 2730 4764 2758
rect 4788 2730 4816 2758
rect 4840 2730 4868 2758
rect 6388 2730 6416 2758
rect 6440 2730 6468 2758
rect 6492 2730 6520 2758
rect 2258 2338 2286 2366
rect 2310 2338 2338 2366
rect 2362 2338 2390 2366
rect 3910 2338 3938 2366
rect 3962 2338 3990 2366
rect 4014 2338 4042 2366
rect 5562 2338 5590 2366
rect 5614 2338 5642 2366
rect 5666 2338 5694 2366
rect 7214 2338 7242 2366
rect 7266 2338 7294 2366
rect 7318 2338 7346 2366
rect 1432 1946 1460 1974
rect 1484 1946 1512 1974
rect 1536 1946 1564 1974
rect 3084 1946 3112 1974
rect 3136 1946 3164 1974
rect 3188 1946 3216 1974
rect 4736 1946 4764 1974
rect 4788 1946 4816 1974
rect 4840 1946 4868 1974
rect 6388 1946 6416 1974
rect 6440 1946 6468 1974
rect 6492 1946 6520 1974
rect 2258 1554 2286 1582
rect 2310 1554 2338 1582
rect 2362 1554 2390 1582
rect 3910 1554 3938 1582
rect 3962 1554 3990 1582
rect 4014 1554 4042 1582
rect 5562 1554 5590 1582
rect 5614 1554 5642 1582
rect 5666 1554 5694 1582
rect 7214 1554 7242 1582
rect 7266 1554 7294 1582
rect 7318 1554 7346 1582
<< metal4 >>
rect 1418 5894 1578 6302
rect 1418 5866 1432 5894
rect 1460 5866 1484 5894
rect 1512 5866 1536 5894
rect 1564 5866 1578 5894
rect 1418 5110 1578 5866
rect 1418 5082 1432 5110
rect 1460 5082 1484 5110
rect 1512 5082 1536 5110
rect 1564 5082 1578 5110
rect 1418 4326 1578 5082
rect 1418 4298 1432 4326
rect 1460 4298 1484 4326
rect 1512 4298 1536 4326
rect 1564 4298 1578 4326
rect 1418 3542 1578 4298
rect 1418 3514 1432 3542
rect 1460 3514 1484 3542
rect 1512 3514 1536 3542
rect 1564 3514 1578 3542
rect 1418 2758 1578 3514
rect 1418 2730 1432 2758
rect 1460 2730 1484 2758
rect 1512 2730 1536 2758
rect 1564 2730 1578 2758
rect 1418 1974 1578 2730
rect 1418 1946 1432 1974
rect 1460 1946 1484 1974
rect 1512 1946 1536 1974
rect 1564 1946 1578 1974
rect 1418 1538 1578 1946
rect 2244 6286 2404 6302
rect 2244 6258 2258 6286
rect 2286 6258 2310 6286
rect 2338 6258 2362 6286
rect 2390 6258 2404 6286
rect 2244 5502 2404 6258
rect 2244 5474 2258 5502
rect 2286 5474 2310 5502
rect 2338 5474 2362 5502
rect 2390 5474 2404 5502
rect 2244 4718 2404 5474
rect 2244 4690 2258 4718
rect 2286 4690 2310 4718
rect 2338 4690 2362 4718
rect 2390 4690 2404 4718
rect 2244 3934 2404 4690
rect 2244 3906 2258 3934
rect 2286 3906 2310 3934
rect 2338 3906 2362 3934
rect 2390 3906 2404 3934
rect 2244 3150 2404 3906
rect 2244 3122 2258 3150
rect 2286 3122 2310 3150
rect 2338 3122 2362 3150
rect 2390 3122 2404 3150
rect 2244 2366 2404 3122
rect 2244 2338 2258 2366
rect 2286 2338 2310 2366
rect 2338 2338 2362 2366
rect 2390 2338 2404 2366
rect 2244 1582 2404 2338
rect 2244 1554 2258 1582
rect 2286 1554 2310 1582
rect 2338 1554 2362 1582
rect 2390 1554 2404 1582
rect 2244 1538 2404 1554
rect 3070 5894 3230 6302
rect 3070 5866 3084 5894
rect 3112 5866 3136 5894
rect 3164 5866 3188 5894
rect 3216 5866 3230 5894
rect 3070 5110 3230 5866
rect 3070 5082 3084 5110
rect 3112 5082 3136 5110
rect 3164 5082 3188 5110
rect 3216 5082 3230 5110
rect 3070 4326 3230 5082
rect 3070 4298 3084 4326
rect 3112 4298 3136 4326
rect 3164 4298 3188 4326
rect 3216 4298 3230 4326
rect 3070 3542 3230 4298
rect 3070 3514 3084 3542
rect 3112 3514 3136 3542
rect 3164 3514 3188 3542
rect 3216 3514 3230 3542
rect 3070 2758 3230 3514
rect 3070 2730 3084 2758
rect 3112 2730 3136 2758
rect 3164 2730 3188 2758
rect 3216 2730 3230 2758
rect 3070 1974 3230 2730
rect 3070 1946 3084 1974
rect 3112 1946 3136 1974
rect 3164 1946 3188 1974
rect 3216 1946 3230 1974
rect 3070 1538 3230 1946
rect 3896 6286 4056 6302
rect 3896 6258 3910 6286
rect 3938 6258 3962 6286
rect 3990 6258 4014 6286
rect 4042 6258 4056 6286
rect 3896 5502 4056 6258
rect 3896 5474 3910 5502
rect 3938 5474 3962 5502
rect 3990 5474 4014 5502
rect 4042 5474 4056 5502
rect 3896 4718 4056 5474
rect 3896 4690 3910 4718
rect 3938 4690 3962 4718
rect 3990 4690 4014 4718
rect 4042 4690 4056 4718
rect 3896 3934 4056 4690
rect 3896 3906 3910 3934
rect 3938 3906 3962 3934
rect 3990 3906 4014 3934
rect 4042 3906 4056 3934
rect 3896 3150 4056 3906
rect 3896 3122 3910 3150
rect 3938 3122 3962 3150
rect 3990 3122 4014 3150
rect 4042 3122 4056 3150
rect 3896 2366 4056 3122
rect 3896 2338 3910 2366
rect 3938 2338 3962 2366
rect 3990 2338 4014 2366
rect 4042 2338 4056 2366
rect 3896 1582 4056 2338
rect 3896 1554 3910 1582
rect 3938 1554 3962 1582
rect 3990 1554 4014 1582
rect 4042 1554 4056 1582
rect 3896 1538 4056 1554
rect 4722 5894 4882 6302
rect 4722 5866 4736 5894
rect 4764 5866 4788 5894
rect 4816 5866 4840 5894
rect 4868 5866 4882 5894
rect 4722 5110 4882 5866
rect 4722 5082 4736 5110
rect 4764 5082 4788 5110
rect 4816 5082 4840 5110
rect 4868 5082 4882 5110
rect 4722 4326 4882 5082
rect 4722 4298 4736 4326
rect 4764 4298 4788 4326
rect 4816 4298 4840 4326
rect 4868 4298 4882 4326
rect 4722 3542 4882 4298
rect 4722 3514 4736 3542
rect 4764 3514 4788 3542
rect 4816 3514 4840 3542
rect 4868 3514 4882 3542
rect 4722 2758 4882 3514
rect 4722 2730 4736 2758
rect 4764 2730 4788 2758
rect 4816 2730 4840 2758
rect 4868 2730 4882 2758
rect 4722 1974 4882 2730
rect 4722 1946 4736 1974
rect 4764 1946 4788 1974
rect 4816 1946 4840 1974
rect 4868 1946 4882 1974
rect 4722 1538 4882 1946
rect 5548 6286 5708 6302
rect 5548 6258 5562 6286
rect 5590 6258 5614 6286
rect 5642 6258 5666 6286
rect 5694 6258 5708 6286
rect 5548 5502 5708 6258
rect 5548 5474 5562 5502
rect 5590 5474 5614 5502
rect 5642 5474 5666 5502
rect 5694 5474 5708 5502
rect 5548 4718 5708 5474
rect 5548 4690 5562 4718
rect 5590 4690 5614 4718
rect 5642 4690 5666 4718
rect 5694 4690 5708 4718
rect 5548 3934 5708 4690
rect 5548 3906 5562 3934
rect 5590 3906 5614 3934
rect 5642 3906 5666 3934
rect 5694 3906 5708 3934
rect 5548 3150 5708 3906
rect 5548 3122 5562 3150
rect 5590 3122 5614 3150
rect 5642 3122 5666 3150
rect 5694 3122 5708 3150
rect 5548 2366 5708 3122
rect 5548 2338 5562 2366
rect 5590 2338 5614 2366
rect 5642 2338 5666 2366
rect 5694 2338 5708 2366
rect 5548 1582 5708 2338
rect 5548 1554 5562 1582
rect 5590 1554 5614 1582
rect 5642 1554 5666 1582
rect 5694 1554 5708 1582
rect 5548 1538 5708 1554
rect 6374 5894 6534 6302
rect 6374 5866 6388 5894
rect 6416 5866 6440 5894
rect 6468 5866 6492 5894
rect 6520 5866 6534 5894
rect 6374 5110 6534 5866
rect 6374 5082 6388 5110
rect 6416 5082 6440 5110
rect 6468 5082 6492 5110
rect 6520 5082 6534 5110
rect 6374 4326 6534 5082
rect 6374 4298 6388 4326
rect 6416 4298 6440 4326
rect 6468 4298 6492 4326
rect 6520 4298 6534 4326
rect 6374 3542 6534 4298
rect 6374 3514 6388 3542
rect 6416 3514 6440 3542
rect 6468 3514 6492 3542
rect 6520 3514 6534 3542
rect 6374 2758 6534 3514
rect 6374 2730 6388 2758
rect 6416 2730 6440 2758
rect 6468 2730 6492 2758
rect 6520 2730 6534 2758
rect 6374 1974 6534 2730
rect 6374 1946 6388 1974
rect 6416 1946 6440 1974
rect 6468 1946 6492 1974
rect 6520 1946 6534 1974
rect 6374 1538 6534 1946
rect 7200 6286 7360 6302
rect 7200 6258 7214 6286
rect 7242 6258 7266 6286
rect 7294 6258 7318 6286
rect 7346 6258 7360 6286
rect 7200 5502 7360 6258
rect 7200 5474 7214 5502
rect 7242 5474 7266 5502
rect 7294 5474 7318 5502
rect 7346 5474 7360 5502
rect 7200 4718 7360 5474
rect 7200 4690 7214 4718
rect 7242 4690 7266 4718
rect 7294 4690 7318 4718
rect 7346 4690 7360 4718
rect 7200 3934 7360 4690
rect 7200 3906 7214 3934
rect 7242 3906 7266 3934
rect 7294 3906 7318 3934
rect 7346 3906 7360 3934
rect 7200 3150 7360 3906
rect 7200 3122 7214 3150
rect 7242 3122 7266 3150
rect 7294 3122 7318 3150
rect 7346 3122 7360 3150
rect 7200 2366 7360 3122
rect 7200 2338 7214 2366
rect 7242 2338 7266 2366
rect 7294 2338 7318 2366
rect 7346 2338 7360 2366
rect 7200 1582 7360 2338
rect 7200 1554 7214 1582
rect 7242 1554 7266 1582
rect 7294 1554 7318 1582
rect 7346 1554 7360 1582
rect 7200 1538 7360 1554
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 2800 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1669390400
transform 1 0 6384 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1669390400
transform -1 0 952 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2 Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 784 0 1 1568
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34 Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 2576 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37
timestamp 1669390400
transform 1 0 2744 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40
timestamp 1669390400
transform 1 0 2912 0 1 1568
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56 Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 3808 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64 Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 4256 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68 Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 4480 0 1 1568
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_72
timestamp 1669390400
transform 1 0 4704 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80
timestamp 1669390400
transform 1 0 5152 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_100
timestamp 1669390400
transform 1 0 6272 0 1 1568
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_104
timestamp 1669390400
transform 1 0 6496 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_107
timestamp 1669390400
transform 1 0 6664 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_115
timestamp 1669390400
transform 1 0 7112 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_2 Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 784 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_66
timestamp 1669390400
transform 1 0 4368 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_70
timestamp 1669390400
transform 1 0 4592 0 -1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_73 Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 4760 0 -1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_105
timestamp 1669390400
transform 1 0 6552 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_113
timestamp 1669390400
transform 1 0 7000 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_115
timestamp 1669390400
transform 1 0 7112 0 -1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_2
timestamp 1669390400
transform 1 0 784 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_34
timestamp 1669390400
transform 1 0 2576 0 1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_37
timestamp 1669390400
transform 1 0 2744 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_101
timestamp 1669390400
transform 1 0 6328 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_105
timestamp 1669390400
transform 1 0 6552 0 1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_108
timestamp 1669390400
transform 1 0 6720 0 1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_2
timestamp 1669390400
transform 1 0 784 0 -1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_34
timestamp 1669390400
transform 1 0 2576 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_65
timestamp 1669390400
transform 1 0 4312 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_69
timestamp 1669390400
transform 1 0 4536 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_73
timestamp 1669390400
transform 1 0 4760 0 -1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_105
timestamp 1669390400
transform 1 0 6552 0 -1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_113
timestamp 1669390400
transform 1 0 7000 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_115
timestamp 1669390400
transform 1 0 7112 0 -1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_2
timestamp 1669390400
transform 1 0 784 0 1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_34
timestamp 1669390400
transform 1 0 2576 0 1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_37
timestamp 1669390400
transform 1 0 2744 0 1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_45
timestamp 1669390400
transform 1 0 3192 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_49
timestamp 1669390400
transform 1 0 3416 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_80
timestamp 1669390400
transform 1 0 5152 0 1 3136
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_96
timestamp 1669390400
transform 1 0 6048 0 1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_104
timestamp 1669390400
transform 1 0 6496 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_108
timestamp 1669390400
transform 1 0 6720 0 1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_2
timestamp 1669390400
transform 1 0 784 0 -1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_5
timestamp 1669390400
transform 1 0 952 0 -1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_37
timestamp 1669390400
transform 1 0 2744 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_39
timestamp 1669390400
transform 1 0 2856 0 -1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_69
timestamp 1669390400
transform 1 0 4536 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_73
timestamp 1669390400
transform 1 0 4760 0 -1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_80
timestamp 1669390400
transform 1 0 5152 0 -1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_112
timestamp 1669390400
transform 1 0 6944 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_2
timestamp 1669390400
transform 1 0 784 0 1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_19
timestamp 1669390400
transform 1 0 1736 0 1 3920
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_37
timestamp 1669390400
transform 1 0 2744 0 1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_43
timestamp 1669390400
transform 1 0 3080 0 1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_74
timestamp 1669390400
transform 1 0 4816 0 1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_108
timestamp 1669390400
transform 1 0 6720 0 1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_2
timestamp 1669390400
transform 1 0 784 0 -1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_34
timestamp 1669390400
transform 1 0 2576 0 -1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_42
timestamp 1669390400
transform 1 0 3024 0 -1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_49
timestamp 1669390400
transform 1 0 3416 0 -1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_60
timestamp 1669390400
transform 1 0 4032 0 -1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_66
timestamp 1669390400
transform 1 0 4368 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_70
timestamp 1669390400
transform 1 0 4592 0 -1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_73
timestamp 1669390400
transform 1 0 4760 0 -1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_105
timestamp 1669390400
transform 1 0 6552 0 -1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_113
timestamp 1669390400
transform 1 0 7000 0 -1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_115
timestamp 1669390400
transform 1 0 7112 0 -1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_2
timestamp 1669390400
transform 1 0 784 0 1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_34
timestamp 1669390400
transform 1 0 2576 0 1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_37
timestamp 1669390400
transform 1 0 2744 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_101
timestamp 1669390400
transform 1 0 6328 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_105
timestamp 1669390400
transform 1 0 6552 0 1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_108
timestamp 1669390400
transform 1 0 6720 0 1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_2
timestamp 1669390400
transform 1 0 784 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_66
timestamp 1669390400
transform 1 0 4368 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_70
timestamp 1669390400
transform 1 0 4592 0 -1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_9_73
timestamp 1669390400
transform 1 0 4760 0 -1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_105
timestamp 1669390400
transform 1 0 6552 0 -1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_113
timestamp 1669390400
transform 1 0 7000 0 -1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_115
timestamp 1669390400
transform 1 0 7112 0 -1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_2
timestamp 1669390400
transform 1 0 784 0 1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_34
timestamp 1669390400
transform 1 0 2576 0 1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_37
timestamp 1669390400
transform 1 0 2744 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_101
timestamp 1669390400
transform 1 0 6328 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_105
timestamp 1669390400
transform 1 0 6552 0 1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_108
timestamp 1669390400
transform 1 0 6720 0 1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_11_2
timestamp 1669390400
transform 1 0 784 0 -1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_34
timestamp 1669390400
transform 1 0 2576 0 -1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_37
timestamp 1669390400
transform 1 0 2744 0 -1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_53
timestamp 1669390400
transform 1 0 3640 0 -1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_69
timestamp 1669390400
transform 1 0 4536 0 -1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_11_72
timestamp 1669390400
transform 1 0 4704 0 -1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_104
timestamp 1669390400
transform 1 0 6496 0 -1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_107
timestamp 1669390400
transform 1 0 6664 0 -1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_115
timestamp 1669390400
transform 1 0 7112 0 -1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_0 Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 672 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_1
timestamp 1669390400
transform -1 0 7280 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_2
timestamp 1669390400
transform 1 0 672 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_3
timestamp 1669390400
transform -1 0 7280 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_4
timestamp 1669390400
transform 1 0 672 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_5
timestamp 1669390400
transform -1 0 7280 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_6
timestamp 1669390400
transform 1 0 672 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_7
timestamp 1669390400
transform -1 0 7280 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_8
timestamp 1669390400
transform 1 0 672 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_9
timestamp 1669390400
transform -1 0 7280 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_10
timestamp 1669390400
transform 1 0 672 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_11
timestamp 1669390400
transform -1 0 7280 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_12
timestamp 1669390400
transform 1 0 672 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_13
timestamp 1669390400
transform -1 0 7280 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_14
timestamp 1669390400
transform 1 0 672 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_15
timestamp 1669390400
transform -1 0 7280 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_16
timestamp 1669390400
transform 1 0 672 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_17
timestamp 1669390400
transform -1 0 7280 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_18
timestamp 1669390400
transform 1 0 672 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_19
timestamp 1669390400
transform -1 0 7280 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_20
timestamp 1669390400
transform 1 0 672 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_21
timestamp 1669390400
transform -1 0 7280 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_22
timestamp 1669390400
transform 1 0 672 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_23
timestamp 1669390400
transform -1 0 7280 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_24 Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 2632 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_25
timestamp 1669390400
transform 1 0 4592 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_26
timestamp 1669390400
transform 1 0 6552 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_27
timestamp 1669390400
transform 1 0 4648 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_28
timestamp 1669390400
transform 1 0 2632 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_29
timestamp 1669390400
transform 1 0 6608 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_30
timestamp 1669390400
transform 1 0 4648 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_31
timestamp 1669390400
transform 1 0 2632 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_32
timestamp 1669390400
transform 1 0 6608 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_33
timestamp 1669390400
transform 1 0 4648 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_34
timestamp 1669390400
transform 1 0 2632 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_35
timestamp 1669390400
transform 1 0 6608 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_36
timestamp 1669390400
transform 1 0 4648 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_37
timestamp 1669390400
transform 1 0 2632 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_38
timestamp 1669390400
transform 1 0 6608 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_39
timestamp 1669390400
transform 1 0 4648 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_40
timestamp 1669390400
transform 1 0 2632 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_41
timestamp 1669390400
transform 1 0 6608 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_42
timestamp 1669390400
transform 1 0 2632 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_43
timestamp 1669390400
transform 1 0 4592 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_44
timestamp 1669390400
transform 1 0 6552 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _02_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 2856 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _03_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 4816 0 -1 3920
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _04_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 4032 0 -1 4704
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _05_
timestamp 1669390400
transform 1 0 4144 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _06_
timestamp 1669390400
transform -1 0 3416 0 -1 4704
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _07_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 5152 0 1 3136
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _08_
timestamp 1669390400
transform -1 0 4816 0 1 3920
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _09_
timestamp 1669390400
transform 1 0 2912 0 -1 3920
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _10_
timestamp 1669390400
transform 1 0 2688 0 -1 3136
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input1 Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 1680 0 1 1568
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input2
timestamp 1669390400
transform -1 0 6272 0 1 1568
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input3
timestamp 1669390400
transform 1 0 840 0 1 3920
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output4 Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 4536 0 -1 6272
box -43 -43 827 435
<< labels >>
flabel metal2 s 1960 0 2016 400 0 FreeSans 224 90 0 0 clka
port 0 nsew signal input
flabel metal2 s 5936 0 5992 400 0 FreeSans 224 90 0 0 clkb
port 1 nsew signal input
flabel metal2 s 3976 7600 4032 8000 0 FreeSans 224 90 0 0 gclk
port 2 nsew signal tristate
flabel metal3 s 0 3976 400 4032 0 FreeSans 224 0 0 0 select
port 3 nsew signal input
flabel metal4 s 1418 1538 1578 6302 0 FreeSans 640 90 0 0 vdd
port 4 nsew power bidirectional
flabel metal4 s 3070 1538 3230 6302 0 FreeSans 640 90 0 0 vdd
port 4 nsew power bidirectional
flabel metal4 s 4722 1538 4882 6302 0 FreeSans 640 90 0 0 vdd
port 4 nsew power bidirectional
flabel metal4 s 6374 1538 6534 6302 0 FreeSans 640 90 0 0 vdd
port 4 nsew power bidirectional
flabel metal4 s 2244 1538 2404 6302 0 FreeSans 640 90 0 0 vss
port 5 nsew ground bidirectional
flabel metal4 s 3896 1538 4056 6302 0 FreeSans 640 90 0 0 vss
port 5 nsew ground bidirectional
flabel metal4 s 5548 1538 5708 6302 0 FreeSans 640 90 0 0 vss
port 5 nsew ground bidirectional
flabel metal4 s 7200 1538 7360 6302 0 FreeSans 640 90 0 0 vss
port 5 nsew ground bidirectional
rlabel metal1 3976 5880 3976 5880 0 vdd
rlabel via1 4016 6272 4016 6272 0 vss
rlabel metal3 4004 4452 4004 4452 0 _00_
rlabel metal3 4004 3836 4004 3836 0 _01_
rlabel metal2 1988 1043 1988 1043 0 clka
rlabel metal2 3164 3192 3164 3192 0 clkapa
rlabel metal2 5964 1043 5964 1043 0 clkb
rlabel metal2 4956 3864 4956 3864 0 clkbpb
rlabel metal3 3808 2884 3808 2884 0 clkpaa
rlabel metal3 4088 3668 4088 3668 0 clkpab
rlabel metal2 4676 3472 4676 3472 0 clkpba
rlabel via2 3612 4508 3612 4508 0 clkpbb
rlabel metal2 4116 6440 4116 6440 0 gclk
rlabel metal2 3052 3976 3052 3976 0 net1
rlabel metal2 5068 3360 5068 3360 0 net2
rlabel metal3 2324 4116 2324 4116 0 net3
rlabel metal2 4284 5250 4284 5250 0 net4
rlabel metal2 980 4032 980 4032 0 select
<< properties >>
string FIXED_BBOX 0 0 8000 8000
<< end >>
