magic
tech gf180mcuC
magscale 1 5
timestamp 1670260779
<< obsm1 >>
rect 672 1538 7360 6302
<< metal2 >>
rect 1008 7600 1064 8000
rect 2968 7600 3024 8000
rect 4928 7600 4984 8000
rect 6888 7600 6944 8000
rect 840 0 896 400
rect 2408 0 2464 400
rect 3976 0 4032 400
rect 5544 0 5600 400
rect 7112 0 7168 400
<< obsm2 >>
rect 854 7570 978 7600
rect 1094 7570 2938 7600
rect 3054 7570 4898 7600
rect 5014 7570 6858 7600
rect 6974 7570 7346 7600
rect 854 430 7346 7570
rect 926 350 2378 430
rect 2494 350 3946 430
rect 4062 350 5514 430
rect 5630 350 7082 430
rect 7198 350 7346 430
<< metal3 >>
rect 0 5936 400 5992
rect 0 1960 400 2016
<< obsm3 >>
rect 400 6022 7351 6286
rect 430 5906 7351 6022
rect 400 2046 7351 5906
rect 430 1930 7351 2046
rect 400 1554 7351 1930
<< metal4 >>
rect 1418 1538 1578 6302
rect 2244 1538 2404 6302
rect 3070 1538 3230 6302
rect 3896 1538 4056 6302
rect 4722 1538 4882 6302
rect 5548 1538 5708 6302
rect 6374 1538 6534 6302
rect 7200 1538 7360 6302
<< labels >>
rlabel metal2 s 2408 0 2464 400 6 INmb
port 1 nsew signal input
rlabel metal2 s 840 0 896 400 6 INpb
port 2 nsew signal input
rlabel metal2 s 5544 0 5600 400 6 OUTm
port 3 nsew signal input
rlabel metal2 s 3976 0 4032 400 6 OUTp
port 4 nsew signal input
rlabel metal3 s 0 5936 400 5992 6 cmnmos
port 5 nsew signal output
rlabel metal3 s 0 1960 400 2016 6 cmpmos
port 6 nsew signal output
rlabel metal2 s 7112 0 7168 400 6 oe
port 7 nsew signal input
rlabel metal2 s 6888 7600 6944 8000 6 omnmos
port 8 nsew signal output
rlabel metal2 s 4928 7600 4984 8000 6 ompmos
port 9 nsew signal output
rlabel metal2 s 2968 7600 3024 8000 6 opnmos
port 10 nsew signal output
rlabel metal2 s 1008 7600 1064 8000 6 oppmos
port 11 nsew signal output
rlabel metal4 s 1418 1538 1578 6302 6 vdd
port 12 nsew power bidirectional
rlabel metal4 s 3070 1538 3230 6302 6 vdd
port 12 nsew power bidirectional
rlabel metal4 s 4722 1538 4882 6302 6 vdd
port 12 nsew power bidirectional
rlabel metal4 s 6374 1538 6534 6302 6 vdd
port 12 nsew power bidirectional
rlabel metal4 s 2244 1538 2404 6302 6 vss
port 13 nsew ground bidirectional
rlabel metal4 s 3896 1538 4056 6302 6 vss
port 13 nsew ground bidirectional
rlabel metal4 s 5548 1538 5708 6302 6 vss
port 13 nsew ground bidirectional
rlabel metal4 s 7200 1538 7360 6302 6 vss
port 13 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 8000 8000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 157044
string GDS_FILE /mnt/c/Users/rmprice/Documents/Github/Trollo/openlane/user_DiffDigota/runs/22_12_05_10_18/results/signoff/DiffDigota.magic.gds
string GDS_START 71906
<< end >>

