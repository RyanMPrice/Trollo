// SPDX-FileCopyrightText: 2022 Ryan M Price
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

module clkgate(
  input       clk
, input       gate
, output wire gclk
);

  wire clki = ~clk;
  reg  clkp;

  assign gclk = clkp & clk;
  
  always @*
    if( clki )
      clkp <= gate;
    else
      clkp <= clkp;
  
  initial clkp = 0;
  
endmodule
