* NGSPICE file created from user_proj_example.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_4 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tieh abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tieh Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_2 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_1 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 D RN CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_2 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai33_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai33_4 A1 A2 A3 B1 B2 B3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai222_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai222_4 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyc_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyc_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_4 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyb_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyb_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_2 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_2 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_4 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai33_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai33_1 A1 A2 A3 B1 B2 B3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai222_1 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_4 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__latq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__latq_1 D E Q VDD VSS
.ends

.subckt user_proj_example io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30]
+ io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12]
+ io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ irq[0] irq[1] irq[2] la_data_in[0] la_data_in[10] la_data_in[11] la_data_in[12]
+ la_data_in[13] la_data_in[14] la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[18]
+ la_data_in[19] la_data_in[1] la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23]
+ la_data_in[24] la_data_in[25] la_data_in[26] la_data_in[27] la_data_in[28] la_data_in[29]
+ la_data_in[2] la_data_in[30] la_data_in[31] la_data_in[32] la_data_in[33] la_data_in[34]
+ la_data_in[35] la_data_in[36] la_data_in[37] la_data_in[38] la_data_in[39] la_data_in[3]
+ la_data_in[40] la_data_in[41] la_data_in[42] la_data_in[43] la_data_in[44] la_data_in[45]
+ la_data_in[46] la_data_in[47] la_data_in[48] la_data_in[49] la_data_in[4] la_data_in[50]
+ la_data_in[51] la_data_in[52] la_data_in[53] la_data_in[54] la_data_in[55] la_data_in[56]
+ la_data_in[57] la_data_in[58] la_data_in[59] la_data_in[5] la_data_in[60] la_data_in[61]
+ la_data_in[62] la_data_in[63] la_data_in[6] la_data_in[7] la_data_in[8] la_data_in[9]
+ la_data_out[0] la_data_out[10] la_data_out[11] la_data_out[12] la_data_out[13] la_data_out[14]
+ la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19]
+ la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24]
+ la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29]
+ la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34]
+ la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39]
+ la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44]
+ la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49]
+ la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54]
+ la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59]
+ la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[6]
+ la_data_out[7] la_data_out[8] la_data_out[9] la_oenb[0] la_oenb[10] la_oenb[11]
+ la_oenb[12] la_oenb[13] la_oenb[14] la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18]
+ la_oenb[19] la_oenb[1] la_oenb[20] la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24]
+ la_oenb[25] la_oenb[26] la_oenb[27] la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30]
+ la_oenb[31] la_oenb[32] la_oenb[33] la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37]
+ la_oenb[38] la_oenb[39] la_oenb[3] la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43]
+ la_oenb[44] la_oenb[45] la_oenb[46] la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4]
+ la_oenb[50] la_oenb[51] la_oenb[52] la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56]
+ la_oenb[57] la_oenb[58] la_oenb[59] la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62]
+ la_oenb[63] la_oenb[6] la_oenb[7] la_oenb[8] la_oenb[9] vdd vss wb_clk_i wb_rst_i
+ wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14]
+ wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1]
+ wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25]
+ wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30]
+ wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8]
+ wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13]
+ wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19]
+ wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24]
+ wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2]
+ wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6]
+ wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11]
+ wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17]
+ wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22]
+ wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28]
+ wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4]
+ wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1]
+ wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
XFILLER_140_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3155_ _0394_ _0400_ _0401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2494__A3 _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2106_ _1204_ _1195_ _1199_ _1205_ _1207_ _1208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XANTENNA_fanout56_I net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3086_ _0322_ _0315_ _0324_ _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_199_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2037_ _0140_ _1133_ _1110_ _1138_ _1139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_58_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_167_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2939_ _0084_ _0163_ _0164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_182_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2954__A1 _1403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2182__A2 _1283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_246_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2890__C2 _1194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_165_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3434__A2 _0707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_201_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1942__I dsynth.csTable.address\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_184_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_232_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1987__A2 _0701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3842_ _1113_ _0020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_242_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3773_ _1232_ _1052_ _1054_ _1055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_164_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2724_ _1685_ _1824_ _1782_ _1825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_157_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2655_ _1245_ _0514_ _1210_ _1756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_146_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2586_ _1594_ _1687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3361__A1 _1586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3207_ _0457_ _0458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_67_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_228_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3138_ _0380_ _0381_ _0383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_83_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3069_ _0303_ _0306_ _0307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__3416__A2 _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_145_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3019__I _1916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2458__A3 _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3655__A2 _0940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_246_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_202_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_127_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2440_ _1533_ _1536_ _1540_ _1541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_154_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2146__A2 _1244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2371_ _1471_ _1472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3646__A2 _0702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_224_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3886__RN net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_177_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3825_ _1100_ _0014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_203_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3756_ _1004_ _0979_ _1021_ _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_14_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2707_ _1662_ _1698_ _1808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_134_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3687_ net8 _0968_ _0969_ _0970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_118_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2638_ _1585_ _1592_ _1739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_82_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_216_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2569_ _1484_ _1669_ _1670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_99_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_181_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_210_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3637__A2 _1544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_216_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_229_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3877__RN net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_245_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_227_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_231_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xuser_proj_example_206 io_oeb[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_149_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xuser_proj_example_217 io_oeb[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_128_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_206_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3868__RN net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1940_ _0272_ _0283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_206_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3610_ _0886_ _0894_ _0901_ _0885_ net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_200_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3541_ _0793_ _0795_ _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_196_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3472_ _0747_ _0749_ _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_142_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2423_ _0382_ _1316_ _1523_ _1163_ _1272_ _1524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_233_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2354_ _1187_ _1231_ _1269_ _1455_ _1456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_229_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_215_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2285_ _0525_ _1387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3619__A2 _0131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_225_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_20_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_213_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2182__B _1217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3808_ _1086_ _0008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_165_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2358__A2 _1312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3739_ _1004_ _0968_ _1021_ _1022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_238_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2201__I _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_173_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3322__A4 _0584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2530__A2 _1618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_125_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2294__A1 _0558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3032__I _1736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_229_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_186_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_245_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_200_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2820__B _1848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_197_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2111__I _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2521__A2 _1270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1950__I _0382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2070_ _0371_ _1172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_93_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2037__A1 _0140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2972_ _0199_ _0200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_241_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2588__A2 _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_187_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1923_ dsynth.csTable.address\[7\] _0096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_163_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3524_ _0751_ _0807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_143_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3455_ _0729_ _0730_ _0731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_118_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2021__I _1118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2406_ _1228_ _1504_ _1507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_48_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3386_ _1382_ _0655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_170_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3561__B _1136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2337_ _1434_ _1438_ _1439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_26_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2268_ _1212_ _1370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3859__CLK net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2199_ _1165_ _1301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_240_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2028__A1 _1123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2028__B2 _1103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2579__A2 _1676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_205_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2200__A1 _1219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2751__A2 _1634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3700__A1 _1445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2503__A2 _1200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_195_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3059__A3 _0279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2267__A1 _1367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_205_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2019__A1 dsynth.freeRunCntr\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2019__B2 _1103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_242_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_236_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2742__A2 _1316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_193_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3240_ _0262_ _0494_ _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_234_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3171_ _0417_ _0418_ _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_239_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2122_ _1223_ _1224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_43_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_212_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2053_ _0899_ _1155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_222_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2955_ _1553_ _0179_ _0180_ _1644_ _0181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_148_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2886_ _1323_ _1403_ _0105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_30_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2981__A2 _0209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2460__B _1217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_198_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3507_ _0782_ _0787_ _0788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_143_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3438_ _0711_ _0703_ _0713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_83_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2497__A1 _1374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3369_ _0632_ _0634_ _0637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_211_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3446__B1 _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_246_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3749__A1 dsynth.freeRunCntr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_224_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_194_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_208_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput20 net20 io_out[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_134_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_235_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_204_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2740_ _0668_ _1258_ _1342_ _1270_ _1206_ _1841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XPHY_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_200_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2671_ _1764_ _1770_ _1771_ _1772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_157_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2176__B1 _1250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3223_ _0474_ _0475_ _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_80_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3676__B1 net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3154_ _0397_ _0399_ _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3691__A3 net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2105_ _1206_ _1207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3085_ _0323_ _0314_ _0324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_167_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2036_ _1136_ _1137_ _1130_ _1138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_fanout49_I net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_223_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2651__A1 _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_206_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2938_ _0981_ _1228_ _1898_ _0163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_241_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2954__A2 _1367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2869_ _1363_ _1490_ _0087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_148_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_232_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2890__B2 _1283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_107_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_218_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2259__C _1360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2881__A1 _0097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_209_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2275__B _1291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1987__A3 _0767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3841_ dsynth.freeRunCntr\[28\] _1112_ _1113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_189_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3189__A2 _0411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3772_ _1044_ _1047_ _1053_ _1054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_207_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2723_ _1691_ _1824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__2936__A2 _0159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2654_ _1173_ _1279_ _1368_ _0789_ _1755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_105_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2585_ _1685_ _1655_ _1686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3361__A2 _1549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_236_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3206_ _0456_ _0241_ _0242_ _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_151_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3137_ _0199_ _0205_ _0381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_82_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3068_ _0304_ _0306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2019_ dsynth.freeRunCntr\[13\] _0991_ _1095_ _1103_ _1110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__2624__A1 _1721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_242_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_164_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2079__C _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2091__A2 _1192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_226_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2370_ dsynth.freeRunCntr\[32\] _1471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_155_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_238_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_224_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3892__CLK net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_205_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2082__A2 _1183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3824_ dsynth.csTable.address\[4\] _1099_ _1100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_242_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3031__A1 _1858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3755_ _1036_ _1037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2706_ _1751_ _1806_ _1807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3686_ net9 _0969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2637_ _1677_ _1692_ _1735_ _1737_ _1738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_160_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2568_ _1486_ _1476_ _1669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_160_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2499_ _1281_ _1432_ _1600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_134_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3098__A1 _1715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2908__B _1587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_228_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_example_207 io_oeb[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_7_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xuser_proj_example_218 io_out[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_109_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_232_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_235_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3013__A1 _0244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3540_ _0793_ _0796_ _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__2367__A3 _1468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3471_ _0636_ _0748_ _0749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_100_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2422_ _0492_ _0239_ _0448_ _1523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2353_ _1289_ _1454_ _1455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_123_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2284_ _0844_ _0228_ _0272_ _1386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_245_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2827__A1 _1906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_231_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout31_I net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3807_ dsynth.freeRunCntr\[17\] _1085_ _1086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_14_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1999_ _0173_ _0931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3738_ _0987_ _1021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_147_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2763__B1 _1863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3669_ _0954_ net1 _0959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_106_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3307__A2 _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_192_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_6428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_138_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_125_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_229_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3491__A1 _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_217_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3243__A1 _0054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_166_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2599__I _1670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_166_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2809__A1 _1207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2971_ _0171_ _0198_ _0199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_206_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2588__A3 _1401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1922_ _0074_ _0085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_128_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3523_ _0751_ _0781_ _0805_ _0806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_155_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2302__I _1360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_235_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3454_ _1576_ _0623_ _0699_ _1634_ _0730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_157_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_217_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2405_ _1505_ _1506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3385_ _0079_ _0653_ _0654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_44_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2336_ _1142_ _1155_ _1239_ _1141_ _1438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__2458__B _0569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_217_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2267_ _1367_ _1368_ _1369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2198_ _1292_ _1296_ _1299_ _1173_ _1300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_93_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_241_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_228_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2193__B _1294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3776__A2 _1056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2200__A2 _0514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2212__I _1313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_235_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_4845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2267__A2 _1368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2672__C1 _1676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3216__A1 _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2019__A2 _0991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_223_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_184_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_199_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2122__I _1223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2742__A3 _1523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3170_ _0166_ _0167_ _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_6_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2121_ _1145_ _1157_ _1223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2052_ _1143_ _1148_ _1150_ _1152_ _1153_ _1154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_75_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2954_ _1403_ _1367_ _1250_ _1406_ _0180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_163_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2885_ _1174_ _0103_ _1334_ _0104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_175_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_219_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_176_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3506_ _0783_ _0786_ _0787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_85_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1941__A1 _0239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3437_ _1765_ _1824_ _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3368_ _0632_ _0634_ _0636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_246_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2497__A2 _1555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2319_ _1319_ _1204_ _1323_ _1328_ _1421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XTAP_3407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3299_ _0557_ _0559_ _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_3418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input11_I io_in[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3446__A1 _0991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3446__B2 _1186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_81_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_220_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2421__A2 _1295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_181_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput21 net21 io_out[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_218_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3437__A1 _1765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_232_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2117__I _0844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1956__I _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2670_ _1767_ _1769_ _1771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_157_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2176__A1 _1179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2176__B2 _1277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_236_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_193_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3222_ _0287_ _0288_ _0475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_98_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3676__A1 net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input3_I io_in[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_239_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3153_ _0398_ _0392_ _0399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2104_ _1192_ _1206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3084_ _0291_ _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2035_ _1010_ _0971_ _1137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_36_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2651__A2 _1302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2027__I _1128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_221_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2937_ _1265_ _1664_ _0161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3600__A1 _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2868_ _1615_ _1706_ _1903_ _0086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_108_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2799_ _1337_ _1489_ _1900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2167__A1 _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3667__A1 net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2890__A2 _0106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_241_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_198_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_220_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2158__A1 _0942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_237_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_174_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2400__I _1500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3840_ dsynth.freeRunCntr\[27\] _1109_ _1112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_220_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3771_ _0873_ _1043_ _1053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2722_ _1640_ _1765_ _1823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_218_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2653_ _1345_ _1351_ _1718_ _1156_ _1318_ _1754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__2149__A1 _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2584_ _1642_ _1685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_86_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_214_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3205_ _1838_ _1493_ _0456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2321__A1 _1394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3136_ _0340_ _0344_ _0379_ _0380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_216_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3067_ _1414_ _1898_ _0304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_97_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2018_ dsynth.freeRunCntr\[14\] _1103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_223_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_225_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_211_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_2_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2615__A2 _1177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2379__A1 _1286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2130__I _1230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3670__B net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2303__A1 _1402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_231_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_221_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3823_ _0349_ _1093_ _1094_ _1099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_222_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3754_ _1027_ _1036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3031__A2 _0260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_174_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2705_ _1779_ _1804_ _1805_ _1806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3685_ net7 _0968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2636_ _1576_ _1736_ _1737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_173_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2567_ _1667_ _1668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__2542__A1 _1347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2498_ _1298_ _1598_ _1281_ _1599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_101_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3098__A2 _0276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2196__B _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3119_ _0330_ _0357_ _0361_ _0362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_244_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_proj_example_208 io_oeb[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_104_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xuser_proj_example_219 io_out[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_109_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_238_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2533__A1 _1633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_150_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2834__B _1579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3013__A2 _1493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3665__B net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3470_ _0741_ _0744_ _0748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_155_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2421_ _1303_ _1295_ _1522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_171_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2524__A1 _1213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_237_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2352_ _1290_ _1287_ _1312_ _1314_ _1453_ _1454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_96_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_96_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2283_ dsynth.freeRunCntr\[4\] _1385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_205_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3806_ dsynth.freeRunCntr\[16\] _1083_ _1085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_159_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1998_ _0811_ _0833_ _0877_ _0909_ _0920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_181_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3737_ _0994_ _1019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2763__A1 _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2763__B2 _1838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3668_ _0951_ _0955_ _0957_ net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_88_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2619_ _1150_ _1251_ _1210_ _1720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_134_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3599_ _0806_ _0817_ _0698_ _0890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_6418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_192_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3491__A2 _0761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_216_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2654__B _1368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_243_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_227_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2203__B1 _1211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2506__A1 _1573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3882__CLK net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_234_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2109__I1 _1210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2548__C _1334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_232_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_235_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2970_ _1630_ _0170_ _0198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_245_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1921_ dsynth.csTable.address\[6\] _0074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2588__A4 _0382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_231_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2745__A1 _1569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3522_ _0803_ _0804_ _0805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_155_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_226_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3453_ _1128_ _1668_ _0729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_143_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2404_ _1227_ _1504_ _1505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_130_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3384_ _0240_ _0612_ _0653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_170_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2739__B _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2335_ _1404_ _1436_ _1437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_217_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2266_ _1275_ _1276_ _1166_ _1368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_84_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2197_ _0942_ _1298_ _1299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_187_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2474__B _1574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2433__B1 _1324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_221_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_222_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_6259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_229_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2672__B1 _1670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2672__C2 _1265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_231_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_101_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2975__A1 _1618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2975__B2 _1734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2831__C _1737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_240_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2403__I _1500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_193_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2120_ _1220_ _1221_ _1214_ _1212_ _1222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_120_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2051_ _0558_ _1049_ _1153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_19_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3455__A2 _0730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2953_ _1220_ _1389_ _1291_ _1370_ _0179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_128_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_203_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2884_ _1619_ _1557_ _0103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2313__I _1414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2718__A1 _1682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_219_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_237_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2194__A2 _1295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3505_ _0784_ _0785_ _0786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_117_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1941__A2 _0283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3436_ _1857_ _0707_ _0628_ _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_28_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3367_ _1818_ _1829_ _0633_ _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2318_ _1347_ _1252_ _1349_ _1420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_111_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3298_ _0541_ _0553_ _0559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_3408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2249_ _1146_ _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3446__A2 _1817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_228_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_178_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput22 net22 io_out[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_6001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_107_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_194_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3134__A1 _0346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_244_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_207_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2948__A1 _1707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_199_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_201_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2133__I _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2176__A2 _1274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3221_ _0460_ _0472_ _0473_ _0474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_45_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_234_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3152_ _0321_ _0358_ _0398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_6590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2103_ _0327_ _0272_ _0679_ _1205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__2509__S _1609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3083_ _0311_ _0322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_3_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2034_ _1135_ _1136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_236_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2752__B _1852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_225_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2936_ _1380_ _0159_ _0160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_148_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2867_ _1137_ _1506_ _0084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2798_ _1127_ _0981_ _1898_ _1899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2167__A2 _1229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_85_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3075__S _0252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3419_ _0685_ _0687_ _0691_ _0692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_232_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3419__A2 _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2662__B _1762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_213_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2158__A2 _1258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_218_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3107__A1 _1838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3107__B2 _1704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_231_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_236_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2330__A2 _1197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_224_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_123_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_166_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1967__I _0569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3770_ _1037_ _1051_ _1052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_160_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2721_ _1684_ _1693_ _1822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_203_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2652_ _1244_ _1153_ _1599_ _1752_ _1753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_195_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2149__A2 _0734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_236_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2583_ _1683_ _1532_ _1684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_177_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_234_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3204_ _0090_ _0451_ _0454_ _0455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_210_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3889__RN net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3135_ _0342_ _0343_ _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_132_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout54_I net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3066_ _1548_ _0114_ _0055_ _0303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_243_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2038__I _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_208_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2017_ _1030_ _1087_ _1095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__2085__A1 dsynth.freeRunCntr\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_51_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2388__A2 _1488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3585__A1 _0868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2919_ _0138_ _0141_ _0142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_143_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_218_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2312__A2 _1413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_232_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2076__A1 _1175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2379__A2 _1479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_237_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2303__A2 _1403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_225_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_4292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2067__A1 _1156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3803__A2 _1077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_220_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3822_ _1098_ _0013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_177_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_165_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_222_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3753_ _1035_ _0031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_18_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2704_ _1802_ _1803_ _1805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_229_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3684_ _0966_ _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_88_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2635_ _1594_ _1736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_12_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2566_ _1666_ _1667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_99_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2542__A2 _1538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2497_ _1374_ _1555_ _1598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_229_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_216_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3118_ _0332_ _0356_ _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_23_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_215_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2058__A1 _0569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3049_ _1428_ _0249_ _0285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_227_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_212_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xuser_proj_example_209 io_oeb[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_137_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2230__A1 _1214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2781__A2 _1880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3730__A1 _0994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2533__A2 _1583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2297__A1 _0129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3549__A1 _0832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_174_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2141__I _1242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2420_ _1351_ _1210_ _1213_ _1521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_142_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2524__A2 _1242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2351_ _1341_ _1452_ _1453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_123_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2282_ _1383_ _1384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_215_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2288__A1 _1291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2288__B2 _1152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2460__A1 _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3805_ _1084_ _0007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1997_ _0888_ _0338_ _0899_ _0909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_119_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3736_ _1018_ _0029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_174_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2763__A2 _1492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3667_ net3 net4 net1 _0957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_179_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2618_ _1148_ _1718_ _1719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_161_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3598_ _0879_ _0882_ _0889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_6408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2549_ _1643_ _1645_ _1647_ _1649_ _1650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_87_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2654__C _0789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_197_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2203__A1 _1301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_221_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3482__A3 _0760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_234_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2136__I _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1920_ dsynth.freeRunCntr\[16\] _0063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3521_ _0798_ _0801_ _0804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_183_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3452_ _1702_ _0159_ _0728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_171_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2403_ _1500_ _1504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_237_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3383_ _0647_ _0648_ _0650_ _0651_ _0652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_69_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2334_ _1434_ _1199_ _1368_ _1436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_85_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2265_ _1245_ _1221_ _1367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_152_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2196_ _1171_ _1297_ _1164_ _1298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_226_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_228_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2433__A1 _1198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2433__B2 _1386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2984__A2 _0211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2490__B _1590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3719_ _0998_ _1002_ _1003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_140_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_192_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_216_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2672__A1 _1311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2672__B2 _1339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_232_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_243_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_227_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2424__A1 _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_242_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_212_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_196_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_153_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_234_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2360__B1 _1365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_239_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2050_ _0338_ _1151_ _1152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_208_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2952_ _1241_ _0176_ _0177_ _1411_ _0178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_182_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3612__B1 _0518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2883_ _1918_ _0100_ _0101_ _0102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_206_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3504_ _1634_ _0623_ _0699_ _1596_ _0785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_143_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3435_ _1128_ _0256_ _0708_ _1498_ _0709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_143_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3366_ _1820_ _1828_ _0633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_217_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2317_ dsynth.freeRunCntr\[2\] _1419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3297_ _0244_ _0526_ _0556_ _0557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_246_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2248_ _1342_ _1343_ _1348_ _1349_ _1350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_26_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2654__A1 _1173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2179_ _1271_ _1281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_96_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2406__A1 _1228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3872__CLK net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_161_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_210_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_222_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput23 net23 io_out[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_190_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_235_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_6068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_193_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2893__A1 _0104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_198_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_213_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_207_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2414__I _1514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_200_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3220_ _0469_ _0471_ _0473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_84_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2333__B1 _1433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3151_ _1444_ _0396_ _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_6580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2884__A1 _1619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2102_ _0503_ _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3082_ _0259_ _0319_ _0320_ _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_5890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_212_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2033_ dsynth.freeRunCntr\[13\] _1135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2636__A1 _1576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3061__A1 _0282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2935_ _1484_ _1669_ _0159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_241_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2866_ _0079_ _0082_ _0083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_223_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2797_ _1501_ _1898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3418_ _1465_ _0689_ _0691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3349_ _0081_ _0614_ _0080_ _0615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_165_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_182_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2618__A1 _1148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_209_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_199_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3043__A1 _1736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2144__I _0283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2720_ _0991_ _1676_ _1683_ _1515_ _1706_ _1821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_157_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2651_ _1328_ _1302_ _1752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_220_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3346__B3 _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2582_ _1566_ _1683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_160_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_218_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3203_ _0252_ _0453_ _0454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_25_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2857__A1 _1906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3134_ _0346_ _0355_ _0377_ _0378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3065_ _0300_ _0301_ _0302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__2609__A1 _1498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_242_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2016_ _0800_ _1078_ _0591_ _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_58_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout47_I net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2085__A2 _1186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_224_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3034__A1 _1736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2918_ _0057_ _0139_ _0047_ _0141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_148_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3585__B3 _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2849_ _0044_ _0062_ _0064_ _0065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_121_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_236_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_137_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2938__B _1898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2848__A1 _0060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2076__A2 _1177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output28_I net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3025__A1 _1429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_230_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_224_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_237_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1978__I _0690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2067__A2 _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3264__A1 _0518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_75_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_177_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3821_ _0349_ _1097_ _1098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_53_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3567__A2 _1118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_242_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3752_ _1031_ _1034_ _1035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_203_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2703_ _1802_ _1803_ _1804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_179_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3683_ net10 _0966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2634_ _1732_ _1734_ _1735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_103_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2565_ _1479_ _1666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_126_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2496_ _1594_ _1596_ _1597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3433__I _1655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3117_ _0325_ _0329_ _0359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_243_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3048_ _0282_ _1678_ _0185_ _1549_ _0284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_93_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2058__A2 _0931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2230__A2 _1331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_232_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2297__A2 _1398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_246_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_206_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3246__A1 _0488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_245_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2350_ _1340_ _1339_ _1384_ _1450_ _1365_ _1451_ _1452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_96_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_229_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2281_ dsynth.freeRunCntr\[6\] _1365_ _1381_ _1382_ _1383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_211_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2288__A2 _1386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2460__A2 _1438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3804_ _1131_ _1083_ _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_165_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1996_ _0261_ _0899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2748__B1 _1616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3735_ _1014_ _1017_ _1018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_140_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3428__I _1584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2332__I _1370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3666_ _0955_ _0956_ _0951_ net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_173_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_238_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2617_ _1219_ _1275_ _1276_ _1718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_133_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3597_ _0818_ _0860_ _0887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_133_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2548_ _1149_ _1648_ _1251_ _1274_ _1334_ _1649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_130_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2479_ _1579_ _1580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_5_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_231_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2451__A2 _0646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_211_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2203__A2 _1302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3400__B2 _0585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_182_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_235_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_207_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_223_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2690__A2 _1766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3520_ _0802_ _0803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_196_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2745__A3 _1845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3451_ _0706_ _0716_ _0727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_170_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2402_ _1502_ _1503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_217_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3382_ dsynth.freeRunCntr\[6\] _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_112_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2333_ _1359_ _1432_ _1433_ _1247_ _1434_ _1435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_123_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2264_ _1357_ _1358_ _1366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_111_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3458__A1 _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2195_ _1196_ _1297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_93_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2327__I _1428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_213_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2433__A2 _1205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3630__A1 _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2197__A1 _0942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1979_ _0646_ _0712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3718_ _0999_ _0992_ _1000_ _1002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3649_ _0906_ _0943_ _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_6206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2946__B _1653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_205_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2672__A2 _1667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2237__I _1338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_197_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_223_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_177_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2951_ _1394_ _1277_ _1392_ _1648_ _1355_ _0177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__1986__I _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3612__A1 _0684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3612__B2 _1445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_108_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2882_ _1506_ _1917_ _0101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_30_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2974__I0 _1786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3503_ _0129_ _1902_ _0784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3434_ _1617_ _0707_ _0708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_174_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3365_ _0620_ _0622_ _0631_ _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XTAP_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2316_ _1385_ _1399_ _1416_ _1417_ _1418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3296_ _0452_ _0545_ _0556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2247_ _0206_ _1349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_226_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2178_ _1147_ _1279_ _1059_ _1179_ _1280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_122_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3851__A1 _1485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_187_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2057__I _1158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2406__A2 _1504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_22_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2590__A1 _1636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput24 net24 io_out[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_159_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_6058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2893__A2 _0110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_232_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_227_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3358__B1 _1640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2430__I _1530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2581__A1 _1681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_193_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_234_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2333__A1 _1359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2333__B2 _1247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3150_ _0395_ _0396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_6570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_239_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2101_ _1195_ _1170_ _1199_ _1201_ _1202_ _1203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_3081_ _0290_ _0318_ _0320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_5880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3261__I _0185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2032_ _1110_ _1130_ _1133_ _1134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_94_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_235_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3833__A1 _0112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2636__A2 _1736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2934_ _0156_ _0157_ _0158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__3061__A2 _1527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_206_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2865_ _0080_ _0081_ _0082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2796_ _1895_ _1896_ _1897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_121_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2572__A1 _1639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xuser_proj_example_190 wbs_dat_o[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_132_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3417_ _0672_ _0604_ _0689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_217_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2324__B2 _1260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_232_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3348_ _1897_ _0078_ _0614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3279_ _0534_ _0537_ _0538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_3218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_227_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_181_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_172_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2079__B1 _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_123_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_200_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2650_ _1699_ _1750_ _1751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_185_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2581_ _1681_ _1653_ _1682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_172_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2306__A1 _1143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_86_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3862__CLK net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3202_ _0090_ _0452_ _0243_ _0453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_132_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input1_I io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_214_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3133_ _0335_ _0345_ _0377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3064_ _0298_ _0299_ _0297_ _0301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_167_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2015_ _1069_ _0393_ _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_149_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2917_ _0050_ _0051_ _0139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_176_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2848_ _0060_ _0061_ _0064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_34_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2779_ _1731_ _1787_ _1880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2070__I _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2545__A1 _0822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2848__A2 _0061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3025__A2 _0256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2784__A1 _1883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2536__A1 _1636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3885__CLK net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_232_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3820_ _1093_ _1094_ _1097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3751_ _1032_ _1025_ _1033_ _1034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2224__B1 _1322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2702_ _1711_ _1748_ _1803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_158_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3682_ _0965_ net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_220_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2633_ _1733_ _1734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_146_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2564_ _1664_ _1631_ _1665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_99_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3861__D net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2495_ _1569_ _1595_ _1596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_142_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3116_ _0330_ _0357_ _0358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_7_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3047_ _1579_ _0282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_58_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2065__I _1166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_197_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2766__A1 _1864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_1735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3182__A1 _1416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2280_ dsynth.freeRunCntr\[5\] _1382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_174_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_237_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_226_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3803_ _1081_ _1077_ _1082_ _1083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1995_ _0316_ _0888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_109_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2748__A1 _1838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2748__B2 _1848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3734_ _1015_ _1008_ _1016_ _1017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_14_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3665_ net3 net4 net1 _0956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_173_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2616_ _1347_ _1716_ _1206_ _1717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_133_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3596_ _0660_ _0696_ _0885_ _0886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_157_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2547_ _1140_ _0228_ _1196_ _1648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_86_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2478_ _1578_ _1579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3476__A2 _0753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_229_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2739__A1 _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_240_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_193_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1962__A2 _0514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2911__A1 _1734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2911__B2 _1581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_216_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1953__A2 dsynth.csTable.address\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3450_ _0717_ _0725_ _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_226_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2401_ _1127_ _1501_ _1502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3381_ _0082_ _0649_ _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_170_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2332_ _1370_ _1434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2263_ _1364_ _1365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3458__A2 _0704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2194_ _1293_ _1295_ _1212_ _1296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_225_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2418__B1 _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_207_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3630__A2 _0707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1978_ _0690_ _0701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_140_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_222_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2197__A2 _1298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3717_ _1417_ _0989_ _1000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_146_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3648_ _0902_ _0941_ _0903_ _0925_ _0943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_175_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_235_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_6207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3579_ _1230_ _0868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_6218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_235_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_164_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_200_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_184_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2253__I _0789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_199_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_229_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3084__I _0291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3688__A2 _0970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2360__A2 _1339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_207_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_212_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_223_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2950_ _1406_ _0767_ _1247_ _1298_ _0176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_206_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3612__A2 _0295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_241_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2881_ _0097_ _0099_ _0100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_148_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2163__I _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3502_ _1129_ _1817_ _0730_ _0783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_239_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2974__I1 _1543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3433_ _1655_ _0707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3364_ _0625_ _0630_ _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_170_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2315_ dsynth.freeRunCntr\[3\] _1417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3295_ _0534_ _0537_ _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_246_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2246_ _1345_ _1346_ _1252_ _1347_ _1348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_66_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2103__A2 _0272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_238_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2177_ _1142_ _1155_ _1279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_199_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_181_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2811__B1 _1251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2073__I _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_202_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput25 net25 io_out[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_66_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_6026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_89_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2957__B _0112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_207_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_201_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_158_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3358__A1 _1702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3358__B2 _0623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_236_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2581__A2 _1653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_171_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2333__A2 _1432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2100_ _0393_ _1202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_6593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3080_ _0290_ _0318_ _0319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_5870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_5881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2031_ _1131_ _1132_ _1129_ _1123_ _1133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_75_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_56_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2933_ _0073_ _0075_ _0157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__3061__A3 _1915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2864_ _1895_ _1896_ _0081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_108_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2795_ _1779_ _1804_ _1896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_144_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_example_180 wbs_dat_o[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_105_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2572__A2 _1657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xuser_proj_example_191 wbs_dat_o[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_85_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3416_ _0685_ _0687_ _0688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2324__A2 _1199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3347_ _0587_ _0605_ _0611_ _0238_ _0612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_98_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3278_ _0532_ _0535_ _0537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_3208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2068__I _0294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2229_ _1141_ _1297_ _1331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_22_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2260__A1 _1125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_107_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2079__B2 _1167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_232_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_157_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_199_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2580_ _1637_ _1681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_12_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2306__A2 _1194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3503__A1 _0129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3201_ _0351_ _0452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_234_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_228_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3132_ _0374_ _0375_ _0376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_6390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_227_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3063_ _0297_ _0298_ _0299_ _0300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_114_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2014_ _1059_ _1069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_223_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_149_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2916_ _0128_ _0136_ _0137_ _0138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_31_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2847_ _0060_ _0061_ _0062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_148_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2778_ _1653_ _1877_ _1878_ _1879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_145_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2481__A1 _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_202_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_224_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2784__A2 _1884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2536__A2 _1595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_221_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3750_ dsynth.freeRunCntr\[7\] _1023_ _1033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2224__B2 _1325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_222_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2701_ _1780_ _1800_ _1801_ _1802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_18_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3681_ net43 tgate.clkp _0965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__3267__I _1415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2632_ _1627_ _1628_ _1578_ _1733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_127_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3724__A1 _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2527__A2 _1626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2563_ _1615_ _1664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_86_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2494_ _1236_ _1355_ _1333_ _1595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__2120__B _1212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_229_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_214_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3115_ _0332_ _0356_ _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_82_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout52_I net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3046_ _0277_ _0280_ _0281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_97_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_225_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2766__A2 _1865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3879_ _0008_ net47 net31 dsynth.freeRunCntr\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_109_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3715__A1 dsynth.freeRunCntr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2518__A2 _1200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_238_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_242_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2206__A1 _1218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2206__B2 _1161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_204_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3182__A2 _0396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_244_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3802_ dsynth.freeRunCntr\[15\] _1080_ _1082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1994_ _0844_ _0855_ _0866_ _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_220_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2748__A2 _1491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3733_ dsynth.freeRunCntr\[5\] _1006_ _1016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3664_ net2 _0955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2615_ _1321_ _1177_ _1716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_133_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3595_ _0818_ _0860_ _0867_ _0884_ _0885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_2546_ _1162_ _1292_ _1646_ _1552_ _1153_ _1647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_115_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2477_ _1577_ _1578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_134_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3029_ _0262_ _0131_ _0260_ _0263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2436__A1 _0690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_243_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3875__CLK net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_224_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2739__A2 _1224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2911__A2 _1858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2675__A1 _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_210_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3624__B1 _1730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2400_ _1500_ _1501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_196_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3380_ _0079_ _0240_ _0612_ _0078_ _1897_ _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_170_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2331_ _1239_ _1432_ _1433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2262_ _1363_ _1364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_38_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2193_ _0888_ _0745_ _1294_ _1295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__2666__A1 _1765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_226_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2418__A1 _1374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_225_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2418__B2 _1327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_206_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1949__B _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3091__A1 _0293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_222_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1977_ _0679_ _0690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3716_ dsynth.freeRunCntr\[3\] _0989_ _0999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_147_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3647_ _0684_ _0295_ _0941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_134_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3578_ dsynth.freeRunCntr\[12\] _0861_ _0862_ _0865_ _1232_ _0867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XTAP_6208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_235_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2529_ _1530_ _1630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_5507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2106__B1 _1199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_229_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2409__A1 _1498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2534__I _1609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_212_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_51_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_240_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_137_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_193_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_238_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2896__A1 _1514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3073__A1 _0175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_204_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2820__A1 _1782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2880_ _1630_ _0098_ _0099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3501_ _1129_ _0395_ _0782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_143_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3432_ _0700_ _0704_ _0705_ _0706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_67_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3363_ _0626_ _0629_ _0630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_28_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2887__A1 _1170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2314_ _1415_ _1416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3294_ _0541_ _0553_ _0554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2245_ _0327_ _0228_ _1347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_230_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3300__A2 _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2176_ _1179_ _1274_ _1250_ _1277_ _1278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_228_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_222_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2303__B _1404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput26 net26 io_out[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_227_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2878__A1 _1642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3134__B _0377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2529__I _1530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_244_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3055__A1 _0284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_241_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2802__A1 _1185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_213_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_184_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_199_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_201_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3358__A2 _1863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2869__A1 _1363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2030_ _1030_ _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_5893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_212_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_236_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3046__A1 _0277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_225_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3597__A2 _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2932_ _0126_ _0154_ _0155_ _0156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_225_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2863_ _1751_ _1806_ _0080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_223_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2794_ _1872_ _1893_ _1894_ _1895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_191_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_proj_example_170 wbs_dat_o[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_181 wbs_dat_o[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_171_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_proj_example_192 wbs_dat_o[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_116_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3415_ _0598_ _0686_ _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_171_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_154_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3346_ _0607_ _0608_ _0597_ _0610_ _0599_ _0603_ _0611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai33_4
XTAP_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2349__I dsynth.freeRunCntr\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3277_ _0523_ _0531_ _0535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2228_ _0833_ _1327_ _1329_ _0963_ _1330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_27_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2159_ _0942_ _1204_ _1163_ _1261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_26_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_226_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3037__A1 _0265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_242_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2084__I _1185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_201_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2548__B1 _1251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_202_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_231_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2720__B1 _1683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_191_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2079__A2 _1179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_207_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2251__A2 _1298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_242_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2878__B _1732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3200_ _0243_ _0451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_171_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3503__A2 _1902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2169__I _0679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3131_ _0365_ _0373_ _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_6380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3062_ _1714_ _0098_ _1687_ _0299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_5690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2013_ _1049_ _1059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_242_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_177_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2915_ _0133_ _0135_ _0137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_221_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2846_ _1876_ _1881_ _0061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_136_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2777_ _1609_ _1713_ _1878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_163_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3329_ _0436_ _0441_ _0592_ _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_218_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2466__C1 _1549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2481__A2 _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_241_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2233__A2 _1295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_237_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3733__A2 _1006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_237_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_224_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_220_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3421__A1 _1385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2700_ _1798_ _1799_ _1801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_203_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3680_ tmux.clkpbb net6 tmux.clkapa vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_118_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_199_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2631_ _1731_ _1732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3724__A2 _0994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2562_ _1480_ _1495_ _1663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2493_ _1590_ _1594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3114_ _0346_ _0355_ _0356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_95_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3045_ _0264_ _0279_ _0280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_fanout45_I net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_227_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2362__I _1463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3878_ _0007_ net50 net33 dsynth.freeRunCntr\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_139_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_192_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2829_ _0043_ _0044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_30_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_238_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3479__A1 _1807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_example_90 io_out[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__2151__A1 _1219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_235_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output26_I net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_199_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout50 net51 net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_70_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2447__I _1547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_225_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3642__A1 _1290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_205_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_221_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3801_ dsynth.freeRunCntr\[15\] _1080_ _1081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1993_ _0426_ _0866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_222_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3732_ dsynth.freeRunCntr\[5\] _1006_ _1015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_18_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3663_ _0951_ net14 net15 net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_122_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2614_ _1531_ _1715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_161_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3594_ _0874_ _0879_ _0882_ _0883_ _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_86_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2545_ _0822_ _0360_ _0547_ _0162_ _1646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_126_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2476_ dsynth.freeRunCntr\[30\] _1499_ _1577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_233_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_214_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_205_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_217_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3028_ _0130_ _0262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_83_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2436__A2 _1295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_200_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2092__I _1193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_238_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2124__A1 _1194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_212_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2675__A2 _1498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_234_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3624__A1 _1103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3624__B2 dsynth.freeRunCntr\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_204_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_237_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2330_ _0261_ _1197_ _1432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_111_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2261_ _1188_ _1362_ _1363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_111_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2192_ _1197_ _1294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2666__A2 _1728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2910__I0 _0130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2418__A2 _0459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3615__A1 _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_228_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3091__A2 _0308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1976_ _0360_ _0679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_119_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3715_ dsynth.freeRunCntr\[4\] _0997_ _0998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_3646_ _1123_ _0702_ _1681_ _1131_ _0939_ _0940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_140_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3577_ _0863_ _0864_ _0865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_6209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_235_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2528_ _1627_ _1628_ _1629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2459_ _1303_ _1555_ _1171_ _1560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_170_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2106__A1 _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2106__B2 _1205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_240_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_243_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_227_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_205_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2896__A2 _0114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_245_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2281__B1 _1381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_182_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_108_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3500_ _0771_ _0774_ _0780_ _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_32_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3431_ _1132_ _0256_ _1700_ _0991_ _1095_ _1668_ _0705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_4
XTAP_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3362_ _0627_ _0628_ _0629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2887__A2 _1523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2313_ _1414_ _1415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3293_ _0546_ _0551_ _0552_ _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2244_ _1141_ _1155_ _1346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_226_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2175_ _1275_ _1276_ _1172_ _1277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_39_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2811__A2 _1346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1959_ _0481_ _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3629_ _0916_ _0921_ _0922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xoutput16 net16 io_out[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_190_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput27 net27 io_out[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_134_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_143_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_235_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_245_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_198_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_242_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_212_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_164_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_234_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_240_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_200_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_184_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3888__CLK net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2318__A1 _1347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_218_1733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_238_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_6584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_204_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2931_ _0152_ _0153_ _0155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_143_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_203_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2862_ _1897_ _0078_ _0079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_175_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2793_ _1891_ _1892_ _1894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_129_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2557__A1 _1639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_example_160 la_data_out[62] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_171 wbs_dat_o[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_116_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xuser_proj_example_182 wbs_dat_o[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_172_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_example_193 wbs_dat_o[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_3414_ _0587_ _0604_ _0675_ _0686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_125_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3345_ _0590_ _0595_ _0609_ _0596_ _0610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_97_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3276_ _0524_ _0526_ _0528_ _0451_ _0534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_246_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2227_ _1238_ _1304_ _1328_ _1180_ _1329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_41_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3285__A2 _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_227_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2158_ _0942_ _1258_ _1259_ _1260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_148_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2089_ _1190_ _1191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3037__A2 _0270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_195_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2548__A1 _1149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2548__B2 _1274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_194_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_107_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2720__A1 _0991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2720__B2 _1515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_184_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_92_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_232_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_220_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_148_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_218_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2711__A1 _1665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3130_ _0365_ _0373_ _0374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_6370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_1730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3061_ _0282_ _1527_ _1915_ _0298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_5680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_212_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2012_ _1040_ _1049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_236_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2185__I _1286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2778__A1 _1653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2914_ _0133_ _0135_ _0136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_3894_ _0025_ net50 net34 dsynth.freeRunCntr\[32\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2845_ _0047_ _0058_ _0059_ _0060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_148_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2776_ _1590_ _1713_ _1609_ _1877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_163_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_236_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3328_ _0439_ _0440_ _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_189_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3259_ _0483_ _0484_ _0516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_3018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2466__B1 _1532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2466__C2 _1566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2769__A1 _1860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_202_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2941__A1 _1415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_215_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3603__B _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_218_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_242_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_179_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2630_ _1577_ _1730_ _1731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3185__A1 _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2561_ _1512_ _1660_ _1661_ _1662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3724__A3 _0996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2492_ _1576_ _1581_ _1585_ _1592_ _1593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_9_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3488__A2 _0642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2160__A2 _1260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3113_ _0348_ _0354_ _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_56_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3044_ _0278_ _0170_ _0054_ _0279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_237_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout38_I net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2620__B1 _1720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3877_ _0006_ net50 net38 dsynth.freeRunCntr\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_197_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_149_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2828_ _1918_ _0037_ _0043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_136_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2759_ _1850_ _1856_ _1859_ _1860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2923__A1 _0142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_219_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_132_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2687__B1 _1732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xuser_proj_example_80 io_out[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_150_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2151__A2 _1166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xuser_proj_example_91 io_out[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_232_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_228_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3100__A1 _1687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_227_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output19_I net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3891__RN net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout40 net41 net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_147_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout51 net52 net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_54_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_210_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_237_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2142__A2 _1175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_211_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3642__A2 _1678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_206_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_220_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3882__RN net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3800_ _1075_ _1080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1992_ _0635_ _0855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3731_ dsynth.freeRunCntr\[6\] _1013_ _1014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_202_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3662_ _0954_ net14 net15 net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_146_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2613_ _1713_ _1714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3593_ _1288_ _0881_ _0883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_173_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2544_ _1149_ _1152_ _1644_ _1645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_157_1745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2475_ _1572_ _1575_ _1576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_130_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_243_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3027_ _0201_ _0260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_227_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_212_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3873__RN net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2322__B _1148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_238_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_235_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3624__A2 _1586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_199_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2283__I dsynth.freeRunCntr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3864__RN net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2060__A1 _0822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3560__A1 _0843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2260_ _1125_ _1350_ _1361_ _1362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_78_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2191_ _1167_ _1246_ _1293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2666__A3 _1766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2910__I1 _0131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_238_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3615__A2 _1848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_228_1746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_207_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_221_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1975_ _0624_ _0657_ _0668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_124_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3714_ _0994_ _0996_ _0997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2051__A1 _0558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3645_ _0916_ _0917_ _0939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3576_ _0815_ _0773_ _0780_ _0864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_235_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2527_ _1621_ _1626_ _1564_ _1628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_157_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2458_ _1156_ _1173_ _1253_ _0569_ _1559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_114_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3303__A1 _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_68_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2389_ _1489_ _1490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_217_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3606__A2 _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_213_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_197_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2290__A1 _1323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_200_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_193_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2227__B _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_203_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2281__A1 dsynth.freeRunCntr\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2281__B2 _1382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_223_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_204_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3430_ _0699_ _1824_ _0703_ _0704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_143_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3361_ _1586_ _1549_ _1852_ _0628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_100_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2312_ _1020_ _1413_ _1414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3292_ _0549_ _0550_ _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2243_ _1275_ _1344_ _1345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_152_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2174_ _0745_ _1276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2024__A1 _1125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_202_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1958_ _0316_ _0481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_124_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3628_ _0917_ _0919_ _0921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput17 net17 io_out[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput28 net28 io_out[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_192_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3559_ _0840_ _0846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_6018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_142_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_244_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_112_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_227_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_158_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3657__I net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_205_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2015__A1 _1069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_227_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_153_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_239_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_235_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_245_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2254__A1 _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2930_ _0152_ _0153_ _0154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_225_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_182_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2861_ _0071_ _0076_ _0077_ _0078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_54_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2792_ _1891_ _1892_ _1893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_102_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2557__A2 _1657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_example_150 la_data_out[52] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_144_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xuser_proj_example_161 la_data_out[63] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_89_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_proj_example_172 wbs_dat_o[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_183 wbs_dat_o[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_116_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_example_194 wbs_dat_o[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_171_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3413_ _0684_ _0685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2420__B _1213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_193_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3344_ _0224_ _0225_ _0606_ _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3275_ _0523_ _0531_ _0532_ _0533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3809__A2 _1085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2226_ _1297_ _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_226_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2157_ _0569_ _1259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_53_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2088_ _1189_ _1190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_241_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2548__A2 _1648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_198_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_163_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_172_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2720__A2 _1676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2484__A1 _1579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2667__S _1703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3060_ _1687_ _1618_ _0297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_5670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2011_ _0074_ dsynth.csTable.address\[4\] _1040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_76_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_225_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2913_ _1635_ _0134_ _0135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_3893_ _0024_ net52 net36 dsynth.freeRunCntr\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_176_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2844_ _0050_ _0057_ _0051_ _0059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_34_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2775_ _1875_ _1853_ _1876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_145_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2950__A2 _0767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3327_ _1399_ _0402_ _0590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_154_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_230_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3258_ _0509_ _0513_ _0515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_3008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_227_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2466__A1 _1515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2209_ _1310_ _1311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_160_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3189_ _0218_ _0411_ _0438_ _0412_ _0420_ _0439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_167_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3878__CLK net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2466__B2 _1544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2941__A2 _1666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2457__A1 _1402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_232_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3709__A1 _1464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2560_ _1614_ _1659_ _1661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_182_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3066__B _0055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2491_ _1586_ _1588_ _1591_ _1592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_153_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3112_ _0350_ _0353_ _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_6190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3043_ _1736_ _0111_ _0113_ _0278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_83_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2620__B2 _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3876_ _0005_ net58 net38 dsynth.freeRunCntr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_176_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2827_ _1906_ _0041_ _0042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_164_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2758_ _1857_ _1858_ _1853_ _1855_ _1859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_151_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2689_ _1531_ _1727_ _1790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_236_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2687__A1 _1618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xuser_proj_example_70 io_oeb[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_134_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_example_81 io_out[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_92 io_out[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_74_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2439__A1 _1433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_246_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2439__B2 _1192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_210_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3100__A2 _1714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3239__I0 _0461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout41 net42 net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_74_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout52 net59 net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_141_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_208_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_155_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3627__B1 _1730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2850__A1 _1883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1991_ _0602_ _0844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3730_ _0994_ _1012_ _1013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2602__A1 _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3661_ _0954_ _0953_ net15 net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2612_ _1633_ _1526_ _1713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_103_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3592_ _1288_ _0881_ _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_133_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_155_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2543_ _1190_ _0173_ _1644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_157_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2474_ _1570_ _1571_ _1574_ _1575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_114_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3618__B1 _1858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout50_I net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3026_ _0242_ _0255_ _0258_ _0259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_58_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2841__A1 _1580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_244_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_205_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3859_ tmux.clkbpb net5 tmux.clkpba vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_164_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2832__A1 _0035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3388__A2 _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2060__A2 _0734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2190_ _0437_ _0261_ _1197_ _1292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_120_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_37_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3076__A1 _1707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_241_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2823__A1 _0035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_228_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3379__A2 _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1974_ _0646_ _0657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_109_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_221_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3713_ _0969_ _0995_ _0996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3644_ _0932_ _0937_ _0938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_134_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3575_ _0779_ _0771_ _0774_ _0863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_196_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_235_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_1729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2526_ _1564_ _1621_ _1626_ _1627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_142_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2457_ _1402_ _1393_ _1556_ _1557_ _1558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_4809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2388_ _1484_ _1488_ _1489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_29_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3067__A1 _1414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_227_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3009_ _0115_ _0241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2814__A1 _1636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_225_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_196_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2290__A2 _1243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_213_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_184_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2052__C _1153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_193_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_238_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3164__B _0410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2805__A1 _1185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_188_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2281__A2 _1365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3360_ _1857_ _1655_ _0627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_125_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2311_ _1400_ _1405_ _1408_ _1412_ _1413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_154_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3291_ _0549_ _0550_ _0551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_170_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2242_ _0811_ _1344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_26_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3297__A1 _0244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2173_ _0712_ _1275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3049__A1 _1428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_213_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1957_ _0459_ _0470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_135_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_179_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3627_ _0063_ _1596_ _1730_ dsynth.freeRunCntr\[13\] _0918_ _0919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
Xoutput18 net18 io_out[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_227_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput29 net29 io_out[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_3558_ _0821_ _0802_ _0823_ _0845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_157_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2509_ _1585_ _1584_ _1609_ _1610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_5307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3489_ _0763_ _0768_ _0769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_5318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3288__A1 _0336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_197_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2063__B _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3212__A1 _0461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_197_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_180_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_218_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_218_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1921__I dsynth.csTable.address\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_236_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2254__A2 _0767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2860_ _1872_ _1893_ _0077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_148_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3203__A1 _0252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2791_ _1780_ _1800_ _1892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_50_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_proj_example_140 la_data_out[42] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_171_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xuser_proj_example_151 la_data_out[53] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_116_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xuser_proj_example_162 wbs_ack_o vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_176_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_proj_example_173 wbs_dat_o[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_171_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xuser_proj_example_184 wbs_dat_o[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_116_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3412_ _1419_ _0684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xuser_proj_example_195 io_oeb[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_131_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2199__I _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3343_ _0606_ _0588_ _0608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3274_ _0496_ _0498_ _0488_ _0532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_234_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2225_ _0492_ _0283_ _1239_ _1327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_41_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2156_ _1257_ _1258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_187_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2087_ dsynth.csTable.address\[5\] _0074_ _1189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_59_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1987__B _0789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2245__A2 _0228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2989_ _0212_ _0218_ _0214_ _0219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_124_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_213_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_190_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3681__A1 net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2484__A2 _1584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_232_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2172__A1 _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_6394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2010_ _1020_ _1030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_94_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3672__A1 net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2912_ _0055_ _0052_ _0053_ _0134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_32_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3892_ _0023_ net51 net35 dsynth.freeRunCntr\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_149_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2843_ _0050_ _0051_ _0057_ _0058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_31_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2774_ _1530_ _1851_ _1875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2950__A3 _1247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_217_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3326_ _0160_ _0588_ _0589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_101_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_218_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3257_ _0482_ _0510_ _0511_ _0512_ _0513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XTAP_3009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2208_ _1020_ _1309_ _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_160_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2466__A2 _1528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3663__A1 _0951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3188_ _0210_ _0211_ _0438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_2308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2139_ _1238_ _1240_ _1069_ _1241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_1607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_241_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_230_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2218__A2 _1316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_208_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2392__I _1492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_224_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_172_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2567__I _1667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_237_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2457__A2 _1393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3406__A1 _0672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1968__A1 _0470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_207_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_229_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_13_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3709__A2 _0989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3347__B _0611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2490_ _1563_ _1565_ _1590_ _1591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_175_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2145__A1 _1245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_229_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2477__I _1577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3111_ _1762_ _0352_ _0353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_6180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_68_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3042_ _0262_ _0276_ _0269_ _0054_ _0277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_5490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_212_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_225_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3875_ _0004_ net58 net38 dsynth.freeRunCntr\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_104_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2826_ _0039_ _0040_ _0041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_118_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2161__B _1262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2757_ _1851_ _1858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_145_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2688_ _1782_ _1783_ _1789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_133_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_235_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2687__A2 _1785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xuser_proj_example_60 io_oeb[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_154_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xuser_proj_example_71 io_oeb[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_63_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_example_82 io_out[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_3309_ _0546_ _0551_ _0571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_219_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xuser_proj_example_93 io_out[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_45_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_58_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3100__A3 _0098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2336__B _1239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_199_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3011__I _0186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout31 net32 net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout42 net45 net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_165_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout53 net57 net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_168_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_178_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3627__B2 dsynth.freeRunCntr\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3630__B _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2850__A2 _1884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1990_ _0481_ _0272_ _0822_ _0833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_166_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3856__I net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_222_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3660_ net11 _0954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_105_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2611_ _1709_ _1710_ _1712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_127_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3591_ _0880_ _0769_ _0881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_196_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3868__CLK net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2542_ _1347_ _1538_ _1209_ _1643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_154_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2473_ _1573_ _1574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_87_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_218_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2000__I _0931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_228_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3618__A1 _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3618__B2 _0655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3025_ _1429_ _0256_ _0257_ _0258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_70_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout43_I net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2841__A2 _0033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3858_ tmux.clkpaa net44 tmux.clkpab vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_149_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2809_ _1207_ _1909_ _1360_ _1910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_164_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3789_ _1070_ _0004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_210_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2066__B _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2293__B1 _1327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_242_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_221_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_237_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2520__A1 _1619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2520__B2 _0195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_234_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_222_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1973_ _0635_ _0646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2587__A1 _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3712_ _0978_ _0968_ _0995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_179_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2423__C _1272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3643_ _0933_ _0934_ _0936_ _0937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_134_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_155_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3574_ _0751_ _0781_ _0808_ _0862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2525_ _1622_ _1623_ _1624_ _1625_ _1626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_192_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2456_ _1555_ _1294_ _1557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_190_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2387_ _1481_ _1485_ _1487_ _1488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_28_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_229_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3067__A2 _1898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3008_ _0231_ _0235_ _0238_ _0240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_71_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_224_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_51_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_212_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2578__A1 _1137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_196_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_203_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2502__A1 _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2575__I _1675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2805__A2 _1706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_243_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2524__B _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_243_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2310_ _1409_ _1410_ _1411_ _1412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3290_ _0462_ _0520_ _0550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_234_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2241_ _1328_ _1222_ _1343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_112_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2172_ _0613_ _0734_ _0822_ _1274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__3049__A2 _0249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2418__C _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_206_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1956_ _0448_ _0459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2153__C _1069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_222_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3626_ _1118_ _0702_ _0918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_116_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput19 net19 io_out[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_3557_ _0812_ _0813_ _0842_ _0843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_190_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2508_ _1578_ _1607_ _1608_ _1609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_143_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3488_ _0618_ _0642_ _0762_ _0768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_5308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2439_ _1433_ _1537_ _1539_ _1192_ _1191_ _1540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_130_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3288__A2 _0276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_57_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2799__A1 _1337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_188_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_213_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_184_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_166_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2519__B _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2239__B1 _1339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_186_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2254__A3 _1247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3451__A2 _0716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2790_ _1873_ _1889_ _1890_ _1891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_34_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_190_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xuser_proj_example_130 la_data_out[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_171_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2962__A1 _1707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xuser_proj_example_141 la_data_out[43] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_152 la_data_out[54] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_116_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xuser_proj_example_163 wbs_dat_o[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_156_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xuser_proj_example_174 wbs_dat_o[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_3411_ _1385_ _0681_ _0682_ _1463_ _0683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
Xuser_proj_example_185 wbs_dat_o[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_172_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xuser_proj_example_196 io_oeb[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_217_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3342_ _0606_ _0588_ _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_28_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3273_ _0529_ _0530_ _0531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2224_ _1315_ _1320_ _1322_ _1325_ _1326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_230_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2155_ _1256_ _1257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2086_ _1010_ _1188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_226_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3442__A2 _0716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_228_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2988_ _0210_ _0211_ _0218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_241_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1939_ _0261_ _0272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_135_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2953__A1 _1220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3609_ _0895_ _0683_ _0896_ _0900_ _0901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_150_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2181__A2 _1282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_177_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_160_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2172__A2 _0734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_190_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3125__S _1664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3121__A1 _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2227__A3 _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2911_ _1734_ _1858_ _0132_ _1581_ _0133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_232_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3891_ _0021_ net49 net34 dsynth.freeRunCntr\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_148_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2842_ _0052_ _0054_ _0056_ _1635_ _0057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_148_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2773_ _1850_ _1856_ _1874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_191_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2003__I _0958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3360__A1 _1857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3325_ _0224_ _0225_ _0588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_112_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3035__S _0268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3256_ _0476_ _0477_ _0512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_112_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3112__A1 _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2207_ _1291_ _1300_ _1308_ _1309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_239_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3187_ _0414_ _0434_ _0435_ _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_187_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3663__A2 net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2138_ _1239_ _1146_ _1240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_167_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2069_ _0327_ _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_208_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_194_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_237_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_150_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3351__A1 _1807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3351__B2 _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_182_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_232_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3894__RN net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_220_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1968__A2 _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3590__A1 _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2393__A2 _1493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_141_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2145__A2 _1246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3110_ _1310_ _0312_ _0351_ _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_6170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_191_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3041_ _0182_ _0183_ _0276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_5480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_184_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2493__I _1590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3885__RN net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3874_ _0003_ net58 net37 dsynth.freeRunCntr\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_242_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_203_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2825_ _1866_ _1867_ _0040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_136_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2756_ _1765_ _1857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_195_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3581__A1 _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2687_ _1618_ _1785_ _1732_ _1787_ _1788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_117_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xuser_proj_example_61 io_oeb[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_98_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3308_ _0562_ _0566_ _0568_ _0570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
Xuser_proj_example_72 io_oeb[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_83 io_out[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_94 io_out[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_86_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3239_ _0461_ _0493_ _0490_ _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_132_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2109__S _0844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3876__RN net58 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2336__C _1141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_208_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout32 net36 net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_167_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout43 net44 net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout54 net57 net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_22_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2072__A1 _1170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_150_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_237_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3627__A2 _1596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3630__C _0922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2686__I0 _1543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3867__RN net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_221_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2063__A1 _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_207_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2610_ _1312_ _1700_ _1709_ _1710_ _1711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_122_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3590_ _0755_ _0761_ _0880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3563__A1 _0843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_196_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2541_ _1473_ _1545_ _1641_ _1642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_86_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2472_ _1001_ _1573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_237_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_229_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3618__A2 _1728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3024_ _0248_ _0254_ _0257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_225_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2437__B _0679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout36_I net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_225_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2054__A1 _0514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_205_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2172__B _0822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3857_ tmux.clkapa net43 tmux.clkpaa vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2808_ _1220_ _1402_ _1550_ _0470_ _1909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_3788_ _1066_ _1068_ _1070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_106_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2739_ _1204_ _1224_ _1180_ _1840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_145_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3306__A1 _0306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_232_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_215_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2293__A1 _1394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2293__B2 _1367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2066__C _1167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_231_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_199_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output17_I net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2045__A1 _0239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_204_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2520__A2 _1272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1940__I _0272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2808__B1 _1550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2284__A1 _0844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_228_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2036__A1 _1136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1972_ _0305_ dsynth.csTable.address\[2\] _0635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_222_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3088__B _1507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3711_ _0966_ _0994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2587__A2 _0833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3642_ _1290_ _1678_ _0935_ _0936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_60_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3536__A1 _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3573_ _0807_ _0805_ _0816_ _0861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_115_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2524_ _1213_ _1242_ _1234_ _1625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_142_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2455_ _1172_ _1555_ _1556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_233_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2386_ _1486_ _1474_ dsynth.freeRunCntr\[29\] _1481_ _1487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_111_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3007_ _0236_ _0237_ _0238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_65_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2275__A1 _1292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_240_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3075__I0 _1311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2578__A2 _1491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_205_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_193_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3017__I _1898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2502__A2 _0195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3858__CLK net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_147_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_230_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_223_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2569__A2 _1669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2741__A2 _1840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_174_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2240_ _1271_ _1294_ _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_238_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2171_ _1270_ _1257_ _1272_ _1273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_65_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_202_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1955_ _0437_ _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_198_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3625_ dsynth.freeRunCntr\[14\] _1586_ _0702_ _1118_ _0917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_200_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3556_ _0799_ _0779_ _0770_ _0842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_1_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2507_ _1602_ _1606_ _1573_ _1608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_153_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3487_ _0747_ _0765_ _0766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_48_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2438_ _1274_ _1150_ _1209_ _1538_ _1539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_130_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2369_ _1470_ net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_211_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2248__A1 _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2799__A2 _1489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_246_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_227_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_212_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_36_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2420__A1 _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_218_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_1737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_5821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2239__A1 _1313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_204_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_231_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_example_120 la_data_out[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_144_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_example_131 la_data_out[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_201_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xuser_proj_example_142 la_data_out[44] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_8_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2270__B _1272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_example_153 la_data_out[55] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_171_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xuser_proj_example_164 wbs_dat_o[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_116_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3410_ _0231_ _0677_ _0682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
Xuser_proj_example_175 wbs_dat_o[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_186 wbs_dat_o[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_197 io_oeb[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_98_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3341_ _1381_ _0402_ _0606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2190__A3 _1197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3272_ _0521_ _0522_ _0530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input8_I io_in[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_239_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2223_ _1323_ _1201_ _1324_ _1325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_78_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2154_ _0888_ _0899_ _0866_ _1256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_227_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2085_ dsynth.freeRunCntr\[12\] _1186_ _1187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_19_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3427__C2 _1576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_206_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2987_ _0169_ _0193_ _0216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_166_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1938_ _0151_ _0250_ _0261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_181_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2953__A2 _1389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3608_ _0897_ _0898_ _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3202__I0 _0090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3539_ _0821_ _0802_ _0823_ _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_115_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2469__A1 _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_123_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_244_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_213_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_199_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_164_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2180__I0 _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2880__A1 _1630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2910_ _0130_ _0131_ _1733_ _0132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_31_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3890_ _0020_ net49 net33 dsynth.freeRunCntr\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_189_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2841_ _1580_ _0033_ _0055_ _0056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3188__A2 _0211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_223_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2772_ _1869_ _1870_ _1873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_129_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2935__A2 _1669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2699__A1 _1798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3360__A2 _1655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3324_ _0444_ _0446_ _0450_ _0586_ _0587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_86_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3255_ _0479_ _0480_ _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_246_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_230_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2206_ _1218_ _1305_ _1307_ _1161_ _1308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_6_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3186_ _0417_ _0418_ _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3663__A3 net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2137_ _0866_ _1239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_226_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2068_ _0294_ _1170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_242_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2623__A1 _1161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_241_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3639__B1 _0707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_232_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3695__I net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_159_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2104__I _1192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3590__A2 _0761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_218_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3040_ _0271_ _0273_ _0274_ _0275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_5470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_236_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_176_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3873_ _0002_ net53 net37 dsynth.freeRunCntr\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_182_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2824_ _1918_ _0037_ _0038_ _0039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_158_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3030__A1 _1580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2755_ _1854_ _1855_ _1856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_157_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2014__I _1059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2686_ _1543_ _1786_ _1652_ _1787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_160_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2949__I _1762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3307_ _0491_ _0543_ _0567_ _0568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xuser_proj_example_62 io_oeb[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_73 io_oeb[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_84 io_out[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_100_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_example_95 irq[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_80_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3238_ _0282_ _0461_ _0493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3097__A1 _1642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_228_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3169_ _0384_ _0387_ _0416_ _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_227_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout33 net35 net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout44 net45 net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_147_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2072__A2 _1173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout55 net56 net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_35_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3021__A1 _0175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_237_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3088__A1 _1414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_218_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2835__A1 _1785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2686__I1 _1786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_220_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2063__A2 _0283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_198_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3358__C _1503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3012__A1 _0129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2540_ _1487_ _1641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_142_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2471_ _1569_ _1570_ _1571_ _1572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_141_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_151_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3023_ _1676_ _0256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_243_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_184_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_209_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2009__I _1010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_205_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2453__B _1396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3856_ net43 _1919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_20_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2807_ _1389_ _1394_ _1907_ _1355_ _1908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_30_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3787_ _1057_ _1061_ _1067_ _1068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_101_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2738_ _1148_ _1718_ _1839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_118_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2669_ _1767_ _1769_ _1770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_156_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2817__A1 _1506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2293__A2 _1277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2045__A2 _1146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3242__A1 _0336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2505__B1 _1605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_232_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2808__A1 _1220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_219_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2808__B2 _0470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2284__A2 _0228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_207_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_221_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1971_ _0613_ _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2273__B _1344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3233__A1 _0306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2036__A2 _1137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3710_ _0993_ _0026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_18_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3784__A2 _1063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_197_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3641_ _1233_ _1683_ _1678_ _1288_ _0935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_122_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3536__A2 _0761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3572_ _0848_ _0856_ _0857_ _0859_ _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_220_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2720__C _1706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2523_ _0668_ _1344_ _1276_ _0778_ _1624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_114_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2454_ _0745_ _1555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2385_ dsynth.freeRunCntr\[30\] _1486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_170_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput1 io_in[11] net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3006_ _0158_ _0229_ _0234_ _0237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_83_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_197_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3224__A1 _1444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3839_ _1111_ _0019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_197_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_238_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2266__A2 _1276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3215__A1 _0252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_187_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2112__I _1213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2170_ _1271_ _1176_ _0184_ _1272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_66_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2257__A2 _1358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3454__A1 _1576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3454__B2 _1634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_228_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_107_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1954_ _0426_ _0437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_159_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3624_ _1103_ _1586_ _1730_ dsynth.freeRunCntr\[13\] _0916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_239_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2717__B1 _1700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3555_ _0820_ _0824_ _0840_ _0841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2022__I _0107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2506_ _1573_ _1602_ _1606_ _1607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_142_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3486_ _0749_ _0764_ _0765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_103_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2437_ _1140_ _0855_ _0679_ _1538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_142_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2178__B _1059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2368_ _1457_ _1469_ _1470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__2496__A2 _1596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_244_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2299_ _0712_ _0811_ _1401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3445__A1 _0718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_169_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_240_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_201_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_205_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_177_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_90_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2420__A2 _1210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3028__I _0130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2184__A1 _1010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2816__B _1916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3436__A1 _1857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2239__A2 _1312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_245_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1946__I dsynth.csTable.address\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2411__A2 _1510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xuser_proj_example_110 la_data_out[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_183_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_proj_example_121 la_data_out[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_156_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xuser_proj_example_132 la_data_out[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__2962__A3 _0172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xuser_proj_example_143 la_data_out[45] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__2270__C _1202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_proj_example_154 la_data_out[56] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_165 wbs_dat_o[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_176 wbs_dat_o[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_187 wbs_dat_o[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_171_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_example_198 io_oeb[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_158_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3340_ _0598_ _0604_ _0605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_67_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3271_ _0243_ _0528_ _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_98_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2222_ _0481_ _0855_ _1196_ _0866_ _1324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_80_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3675__A1 net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2153_ _1214_ _1243_ _1224_ _1205_ _1069_ _1255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_226_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3427__A1 _1596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2084_ _1185_ _1186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3427__B2 _0623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_222_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_245_1691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2986_ _0213_ _0214_ _0215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_202_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1937_ dsynth.csTable.address\[0\] _0250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_175_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3607_ _1464_ _0682_ _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_174_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3202__I1 _0452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3538_ _0804_ _0751_ _0823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_103_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3469_ _0740_ _0746_ _0747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_5118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_213_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2469__A2 _0833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_123_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3418__A1 _1465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_241_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3354__B1 _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_190_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_190_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_6353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2180__I1 _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_235_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_224_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2880__A2 _0098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_231_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2840_ _1591_ _0055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_73_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2771_ _1862_ _1871_ _1872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_184_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2148__A1 _1242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2699__A2 _1799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3323_ _0517_ _0585_ _0586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_217_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2300__I _1401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3254_ _0321_ _0358_ _0510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2205_ _1304_ _1201_ _1306_ _1178_ _1307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_26_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3185_ _0417_ _0418_ _0434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_227_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2136_ _1237_ _1238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout59_I net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2871__A2 _1398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2067_ _1156_ _1159_ _1161_ _1168_ _1169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_82_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_206_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2969_ _0196_ _0197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_52_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_159_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2210__I _1311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3639__A1 _0868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3639__B2 _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_4236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2311__A1 _1400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_213_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2378__A1 _1473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_155_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_209_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3872_ _0001_ net53 net37 dsynth.freeRunCntr\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_176_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2823_ _0035_ _0036_ _0038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_223_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2754_ _1679_ _1763_ _1855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_160_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3030__A2 _1528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2685_ _1541_ _1542_ _1577_ _1786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_172_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2541__A1 _1473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2030__I _1030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3306_ _0306_ _0565_ _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_58_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_example_63 io_oeb[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_140_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_example_74 io_oeb[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_115_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xuser_proj_example_85 io_out[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_189_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_example_96 irq[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_230_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3237_ _0490_ _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_171_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3097__A2 _0336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3168_ _0385_ _0386_ _0416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2119_ _0239_ _1221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_15_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3099_ _0337_ _0339_ _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout34 net35 net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout45 net46 net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_211_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout56 net57 net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_168_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3088__A2 _1675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3012__A2 _1442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2470_ _0800_ _1078_ _1333_ _0580_ _1571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_126_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_237_1730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_218_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2523__A1 _0668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3022_ _0248_ _0254_ _0255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_5290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3855_ _1122_ _0000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2806_ _0525_ _1619_ _1211_ _1393_ _1907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_140_1743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3786_ _0697_ _1056_ _1067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_164_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2737_ _1124_ _1309_ _1838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_117_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2668_ _1503_ _1768_ _1769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_145_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_161_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2599_ _1670_ _1700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_87_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2817__A2 _1917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_210_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_227_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_216_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_184_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3242__A2 _0260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_100_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2753__A1 _1630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2505__A1 _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_219_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2505__B2 _1193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_218_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2808__A2 _1402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3481__A2 _0753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1970_ _0602_ _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2273__C _1223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3233__A2 _0452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3640_ _1233_ _1683_ _0048_ _1230_ _0934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_186_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3571_ _0841_ _0858_ _1103_ _0859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_161_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2744__A1 _1396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2522_ _1143_ _1346_ _1396_ _1623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_155_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2453_ _1551_ _1553_ _1396_ _1554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_216_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3881__CLK net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2384_ dsynth.freeRunCntr\[30\] _1474_ _1485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_96_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput2 io_in[12] net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_237_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3005_ _0233_ _0236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_209_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_196_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3224__A2 _0256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_221_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2983__A1 _0208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3838_ dsynth.freeRunCntr\[27\] _1109_ _1111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_137_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3527__A3 _0611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3769_ _1050_ _0988_ _1051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_118_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2735__A1 _1807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output22_I net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2423__B1 _1523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_137_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3151__A1 _1444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3454__A2 _0623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_207_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2284__B _0272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_221_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1953_ _0305_ dsynth.csTable.address\[3\] _0426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_203_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3623_ _1131_ _1681_ _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_190_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2717__A1 _1229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2717__B2 _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3554_ _0825_ _0839_ _0840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_227_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3843__B _1477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2505_ _1159_ _1603_ _1605_ _1193_ _1606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_239_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3485_ _0762_ _0763_ _0764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_142_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2436_ _0690_ _1295_ _1317_ _1537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_115_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2459__B _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2367_ _1269_ _1458_ _1468_ _1469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__2178__C _1179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_243_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2350__C1 _1365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2298_ _1344_ _1198_ _1386_ _1059_ _1400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_56_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2194__B _1212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_197_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_94_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_36_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2956__A1 _0112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_201_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_222_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_197_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_87_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_198_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3436__A2 _0707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_210_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_203_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1998__A2 _0833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2947__A1 _1715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xuser_proj_example_100 la_data_out[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_111 la_data_out[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_117_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_example_122 la_data_out[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_172_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_example_133 la_data_out[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_7_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_example_144 la_data_out[46] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_116_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xuser_proj_example_155 la_data_out[57] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_166 wbs_dat_o[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_109_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xuser_proj_example_177 wbs_dat_o[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_188 wbs_dat_o[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_109_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xuser_proj_example_199 io_oeb[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XANTENNA__2175__A2 _1276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3270_ _0524_ _0526_ _0527_ _0528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_87_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2221_ _1175_ _1323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_26_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2152_ _1250_ _1252_ _1253_ _1254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_38_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2083_ _1184_ _1185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_187_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_234_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_222_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2985_ _0142_ _0143_ _0214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_166_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1936_ _0228_ _0239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2033__I dsynth.freeRunCntr\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3606_ _0685_ _0687_ _0692_ _0897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_174_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3537_ _0799_ _0777_ _0773_ _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_131_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3468_ _0741_ _0744_ _0746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_5108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2419_ _0789_ _1518_ _1519_ _1520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2469__A3 _1161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3399_ _0666_ _0667_ _0669_ _0447_ _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_130_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3418__A2 _0689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_232_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_226_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_181_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3354__A1 _1186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3354__B2 _1229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_218_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3106__A1 _1338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_212_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_229_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2118__I _1219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_216_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1957__I _0459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2770_ _1869_ _1870_ _1871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3593__A1 _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2148__A2 _1158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3322_ _0485_ _0513_ _0582_ _0584_ _0585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_140_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3253_ _0504_ _0507_ _0508_ _0509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2204_ _1221_ _0701_ _1200_ _1306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3184_ _0407_ _0422_ _0432_ _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_67_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_226_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2135_ _0657_ _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3888__RN net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3412__I _1419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_242_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2066_ _0503_ _1163_ _1165_ _1167_ _1168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_241_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3568__B _0854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_224_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2968_ _0169_ _0193_ _0194_ _0196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2387__A2 _1485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2899_ _0117_ _0119_ _0120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_15_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2139__A2 _1240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3639__A2 _1640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3879__RN net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_198_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_230_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_70_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3327__A1 _1399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_191_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_237_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_224_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_223_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_220_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3871_ _0032_ net53 net37 dsynth.freeRunCntr\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_127_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2822_ _0035_ _0036_ _0037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_176_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_203_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2753_ _1630_ _1851_ _1853_ _1854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_199_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2684_ _1594_ _1651_ _1785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_12_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3305_ _0306_ _0565_ _0566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_154_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_proj_example_64 io_oeb[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_98_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xuser_proj_example_75 io_out[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_86 io_out[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_97 irq[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_3236_ _0278_ _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_100_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3167_ _0367_ _0370_ _0413_ _0414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_66_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2118_ _1219_ _1220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_215_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3098_ _1715_ _0276_ _0339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2049_ _1144_ _0250_ _1151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_54_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfanout35 net36 net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_165_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout46 net13 net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout57 net58 net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_195_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3557__A1 _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2780__A2 _1880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2221__I _1175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_207_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3548__A1 _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2220__A1 _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_182_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_237_1742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3020__I0 _1365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2523__A2 _1344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_209_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3021_ _0175_ _0253_ _0254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_5280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_225_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3854_ dsynth.freeRunCntr\[0\] _0972_ _1122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_123_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2805_ _1185_ _1706_ _1901_ _1905_ _1906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_34_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3785_ _1064_ _1065_ _1066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_160_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2736_ _1836_ _1837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_117_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2762__A2 _1488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2667_ _1705_ _1702_ _1703_ _1768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_195_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_236_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2598_ _1511_ _1662_ _1698_ _1699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_113_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2514__A2 _1500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3219_ _0469_ _0471_ _0472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2216__I _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2450__A1 _0701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3047__I _1579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_85_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_226_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2126__I _1227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_187_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3666__B _0951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_204_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3570_ _0853_ _0858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2744__A2 _1843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2521_ _1517_ _1270_ _1622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_154_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2452_ _1240_ _1552_ _1553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_237_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2383_ _1483_ _1484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_64_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput3 io_in[13] net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3004_ _0233_ _0234_ _0235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_52_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_224_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout34_I net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_240_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2983__A2 _0209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3837_ dsynth.freeRunCntr\[26\] _1107_ _1109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_203_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3768_ _1021_ _1050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2719_ _1680_ _1695_ _1819_ _1820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3699_ dsynth.freeRunCntr\[2\] _0982_ _0983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_105_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_216_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2655__B _1210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_243_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2423__A1 _0382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_243_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2423__B2 _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_196_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_221_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2187__B1 _1287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_183_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3151__A2 _0396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_239_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_206_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2662__A1 _1616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1952_ _0206_ _0404_ _0415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_241_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_221_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3622_ _0906_ _0907_ _0908_ _0913_ _0914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_11_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_128_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2717__A2 _1817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3553_ _0788_ _0791_ _0826_ _0838_ _0839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_155_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2504_ _1165_ _1257_ _1604_ _1605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_142_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3484_ _0636_ _0748_ _0763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_143_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2435_ _1191_ _1534_ _1535_ _1536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_174_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2366_ _1446_ _1460_ _1462_ _1467_ _1468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_233_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_229_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2297_ _0129_ _1398_ _1399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_211_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_225_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2653__A1 _1345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3150__I _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2653__B2 _1156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_221_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_218_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_238_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_6569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_204_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3871__CLK net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_203_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2947__A2 _0170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_200_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xuser_proj_example_101 la_data_out[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_201_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_proj_example_112 la_data_out[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_71_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xuser_proj_example_123 la_data_out[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_134 la_data_out[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_116_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_proj_example_145 la_data_out[47] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_8_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xuser_proj_example_156 la_data_out[58] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_137_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_example_167 wbs_dat_o[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_178 wbs_dat_o[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_109_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_example_189 wbs_dat_o[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_217_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3235__I _0461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2220_ _1237_ _1321_ _1177_ _0195_ _1322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_191_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3675__A3 net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2151_ _1219_ _1166_ _1192_ _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_238_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2082_ _1124_ _1183_ _1184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_35_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_228_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_1671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2984_ _0210_ _0211_ _0212_ _0213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_21_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2938__A2 _1228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_241_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1935_ _0217_ _0228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3060__A1 _1687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2314__I _1415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3605_ _1465_ _0689_ _0694_ _0896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_162_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3536_ _0755_ _0761_ _0819_ _0820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_239_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3467_ _0620_ _0742_ _0743_ _0744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_170_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2418_ _1374_ _0459_ _1159_ _1327_ _0778_ _1519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_112_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3398_ _0403_ _0424_ _0445_ _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_130_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2349_ dsynth.freeRunCntr\[6\] _1451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_170_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_244_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input14_I io_in[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_244_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_207_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2425__S _0958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3354__A2 _1817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3106__A2 _0249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_236_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2617__A1 _1219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_229_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3042__B2 _0054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2134__I _1235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_199_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3321_ _0508_ _0583_ _0584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_154_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3252_ _0469_ _0471_ _0460_ _0508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_26_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input6_I io_in[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_234_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2203_ _1301_ _1302_ _1211_ _1304_ _1069_ _1305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_140_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3183_ _0409_ _0421_ _0432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_239_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2134_ _1235_ _1236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_212_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2309__I _1218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2065_ _1166_ _1167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2608__A1 _1702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_226_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2608__B2 _1503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2967_ _0191_ _0192_ _0194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2898_ _1505_ _1917_ _0100_ _0119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_191_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3519_ _0799_ _0801_ _0802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_103_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_24_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2847__A1 _0060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2219__I _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_232_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3327__A2 _0402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_218_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2838__B _1587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2066__A2 _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3263__A1 _0518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3870_ _0031_ net54 net41 dsynth.freeRunCntr\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_32_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2821_ _1615_ _1849_ _0036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__3015__A1 _0244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_242_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2752_ _1527_ _1547_ _1852_ _1853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_173_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2683_ _1782_ _1783_ _1784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_160_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3304_ _0561_ _0564_ _0565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_101_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_proj_example_65 io_oeb[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_76 io_out[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_100_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xuser_proj_example_87 io_out[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_3235_ _0461_ _0489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_140_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_proj_example_98 la_data_out[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_67_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3166_ _1428_ _1667_ _0372_ _0413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_94_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2117_ _0844_ _1219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_214_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3097_ _1642_ _0336_ _1635_ _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_227_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2048_ _1149_ _1150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_208_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout36 net39 net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_22_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout47 net48 net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout58 net59 net58 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_167_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_221_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_237_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_219_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_219_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_173_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_220_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3796__A2 _1071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3548__A2 _0396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2523__A3 _1276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_229_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3020_ _1365_ _0251_ _0252_ _0253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_5270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3853_ _1121_ _0025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_203_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2804_ _1380_ _1902_ _1904_ _1905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_118_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3784_ _1135_ _1063_ _1065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_192_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2735_ _1807_ _1835_ _1836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_246_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2666_ _1765_ _1728_ _1766_ _1767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_161_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2597_ _1672_ _1697_ _1698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_138_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3218_ _0265_ _0270_ _0273_ _0471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_60_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3149_ _1700_ _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_231_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2450__A2 _1550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_191_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2674__C1 _1675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_246_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3218__A1 _0265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_221_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_222_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2441__A2 _1540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_201_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2520_ _1619_ _1272_ _1620_ _0195_ _1234_ _1621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_127_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1952__A1 _0206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2451_ _1140_ _0646_ _0437_ _1552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_142_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1981__I _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_233_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2298__B _1059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2382_ _1481_ _1482_ _1483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_9_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3457__A1 _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput4 io_in[14] net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3003_ _0156_ _0157_ _0234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_225_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_178_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3836_ _1108_ _0018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3767_ _1048_ _0001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2196__A1 _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_238_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2718_ _1682_ _1694_ _1819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_3698_ _0969_ _0966_ _0980_ _0982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_195_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2649_ _1711_ _1748_ _1749_ _1750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_160_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2499__A2 _1432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2120__A1 _1220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_223_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2423__A2 _1316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3058__I _0114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2187__A1 _1233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2187__B2 _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_234_1724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3687__A1 net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_238_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2662__A2 _1761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_241_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1951_ _0294_ _0393_ _0404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_187_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3611__A1 _1463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3621_ _0910_ _0911_ _0912_ _0913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_174_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3552_ _0827_ _0837_ _0838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_239_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2503_ _1303_ _1200_ _1604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3483_ _0638_ _0641_ _0762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_192_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2434_ _0184_ _1271_ _1274_ _1535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_130_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2365_ _1464_ _1416_ _1466_ _1341_ _1467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_111_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2296_ _1390_ _1391_ _1397_ _1398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_110_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2653__A2 _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3850__A1 _1485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_240_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_212_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3819_ _1096_ _0012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_203_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_161_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3669__A1 _0954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2341__A1 _1030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_proj_example_102 la_data_out[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_113 la_data_out[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_156_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_proj_example_124 la_data_out[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_135 la_data_out[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_144_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xuser_proj_example_146 la_data_out[48] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_157 la_data_out[59] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_168 wbs_dat_o[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_179 wbs_dat_o[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_124_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_234_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2150_ _1251_ _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2883__A2 _0100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2081_ _1154_ _1169_ _1182_ _1183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_94_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3832__A1 _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2983_ _0208_ _0209_ _0212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_72_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2399__A1 _1477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1934_ _0151_ dsynth.csTable.address\[2\] _0217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__3060__A2 _1618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3604_ _0661_ _0662_ _0665_ _0895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_159_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3535_ _0799_ _0777_ _0770_ _0819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_137_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3426__I _1857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3466_ _0622_ _0631_ _0743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_83_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2417_ _0756_ _1517_ _1211_ _1281_ _1518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_130_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3397_ _0427_ _0424_ _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2323__A1 _1404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_233_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2348_ _1418_ _1448_ _1449_ _1450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_218_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_211_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2279_ _1380_ _1381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_2_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_213_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_224_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_197_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_6323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_197_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3042__A2 _0276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_200_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_223_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2150__I _1251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3320_ _0504_ _0507_ _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3251_ _0505_ _0506_ _0507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2202_ _1303_ _1304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3182_ _1416_ _0396_ _0431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_230_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2133_ _1234_ _1235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_152_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2064_ _0811_ _1166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2608__A2 _1704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_207_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3033__A2 _1728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2966_ _0191_ _0192_ _0193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_147_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2897_ _1704_ _0116_ _0117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_162_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3156__I _0396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2544__A1 _1149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3518_ _0739_ _0775_ _0801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3449_ _0720_ _0724_ _0725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_76_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2847__A2 _0061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_182_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_207_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_205_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_176_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2820_ _1782_ _0034_ _1848_ _1531_ _0035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_34_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3015__A2 _1493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_158_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2751_ _1590_ _1634_ _1852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_191_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2774__A1 _1530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2682_ _1732_ _1730_ _1733_ _1783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_157_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3884__CLK net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_236_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3303_ _0542_ _0563_ _0564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_152_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xuser_proj_example_66 io_oeb[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_3234_ _0241_ _0487_ _0488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_234_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_example_77 io_out[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_246_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_example_88 io_out[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_189_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xuser_proj_example_99 la_data_out[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_171_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_239_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3165_ _0210_ _0211_ _0411_ _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_228_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2116_ _1217_ _1218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3096_ _0098_ _0336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_fanout57_I net58 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2047_ _0481_ _0646_ _0426_ _1149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_23_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2055__I dsynth.csTable.address\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout37 net38 net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_11_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout48 net52 net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout59 net12 net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_56_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2949_ _1762_ _0175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_210_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2765__A1 _1364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3614__I dsynth.freeRunCntr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_241_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2220__A3 _1177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_202_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1979__I _0646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3852_ _1473_ _1120_ _1121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_242_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_220_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2803_ _1901_ _1903_ _1904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_165_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3783_ _1136_ _1063_ _1064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2603__I _1703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2734_ _1834_ _1832_ _1835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_195_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2665_ _1547_ _1544_ _1597_ _1766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_145_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2596_ _1674_ _1696_ _1697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_160_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3217_ _0466_ _0467_ _0468_ _0469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_41_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3148_ _0321_ _0358_ _0392_ _0394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_227_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3079_ _0309_ _0317_ _0318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_167_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_224_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_223_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2738__A1 _1148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3466__A2 _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_246_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2674__B1 _1670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2674__C2 _1286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_233_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3218__A2 _0270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2450_ _0701_ _1550_ _1551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_127_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2381_ dsynth.freeRunCntr\[29\] _1482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_83_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3457__A2 _0704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput5 io_in[21] net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_211_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3002_ _0232_ _0077_ _0233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_5090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_92_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_227_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_206_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_209_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2417__B1 _1211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_196_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3835_ dsynth.freeRunCntr\[26\] _1107_ _1108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_192_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3766_ _1044_ _1047_ _1048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_119_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2717_ _1229_ _1817_ _1700_ _1266_ _1818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_145_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3697_ _0978_ _0979_ _0980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_161_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2648_ _1746_ _1747_ _1749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_160_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2579_ _1185_ _1676_ _1515_ _1678_ _1679_ _1680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_99_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_236_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3620__A2 _0033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2187__A2 _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_193_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1934__A2 dsynth.csTable.address\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_234_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2619__S _1210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1950_ _0382_ _0393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3611__A2 _0489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_159_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3620_ _1451_ _0033_ _0912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3551_ _0830_ _0836_ _0837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_143_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2502_ _1234_ _0195_ _1321_ _1603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_170_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3482_ _0757_ _0759_ _0760_ _0761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_44_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_131_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2433_ _1198_ _1205_ _1324_ _1386_ _1317_ _1534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_233_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2364_ _1465_ _1444_ _1449_ _1466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_97_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2350__A2 _1339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2295_ _1360_ _1392_ _1353_ _1395_ _1396_ _1397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_42_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2328__I _1429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_181_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_205_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3818_ _1093_ _1094_ _1096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_197_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3749_ dsynth.freeRunCntr\[7\] _1023_ _1032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_179_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_173_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3669__A2 net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_6538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2341__A2 _1442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2238__I dsynth.freeRunCntr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output20_I net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_216_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_223_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_example_103 la_data_out[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_114 la_data_out[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_156_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_example_125 la_data_out[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_136 la_data_out[38] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_7_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xuser_proj_example_147 la_data_out[49] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_158 la_data_out[60] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_125_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xuser_proj_example_169 wbs_dat_o[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_10_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_152_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2080_ _0206_ _1174_ _1181_ _0963_ _1182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_46_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2982_ _0188_ _0189_ _0211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_61_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3596__A1 _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1933_ _0195_ _0206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3603_ _0887_ _0891_ _0893_ _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_239_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3534_ _0698_ _0806_ _0817_ _0818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_85_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2571__A2 _1665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3465_ _0622_ _0631_ _0742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2416_ _1171_ _1172_ _1517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3396_ _0394_ _0400_ _0666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_213_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2323__A2 _0767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2347_ dsynth.freeRunCntr\[4\] _1399_ _1381_ _1382_ _1449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_96_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2278_ _1379_ _1380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_183_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_240_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2562__A2 _1495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_231_1739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_196_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_236_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_235_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2617__A3 _1276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_232_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3578__A1 dsynth.freeRunCntr\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3578__B2 _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3750__A1 dsynth.freeRunCntr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2553__A2 _1653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3250_ _0501_ _0502_ _0506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_65_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2201_ _0371_ _1303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2305__A2 _1301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3181_ _0427_ _0428_ _0429_ _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_78_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2132_ _1190_ _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_227_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2063_ _0492_ _0283_ _1164_ _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_240_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_222_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3281__A3 _0539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3211__B _0260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2606__I _1703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3569__A1 _1136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_210_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2965_ _0092_ _0093_ _0192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_206_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2241__A1 _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2896_ _1514_ _0114_ _0115_ _0116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_147_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3741__A1 _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2544__A2 _1152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3517_ _0798_ _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_235_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3448_ _0721_ _0722_ _0724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_217_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3379_ _1837_ _0616_ _0648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_241_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2516__I _1616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2480__A1 _1566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_224_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2960__B _0186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_119_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_209_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_6154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_89_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2200__B _1213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_204_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_72_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2471__A1 _1569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3015__A3 _1786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2223__A1 _1323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2750_ _1761_ _1851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_223_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_184_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_199_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2681_ _1588_ _1782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_201_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3302_ _0276_ _0493_ _0548_ _0563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_141_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xuser_proj_example_67 io_oeb[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_214_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3233_ _0306_ _0452_ _0486_ _0487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xuser_proj_example_78 io_out[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_230_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_proj_example_89 io_out[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_136_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3164_ _0383_ _0388_ _0410_ _0411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_82_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2115_ _1191_ _1217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3095_ _0333_ _0307_ _0334_ _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_39_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2046_ _1147_ _1148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_223_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout38 net39 net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout49 net51 net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_211_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2214__A1 _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2948_ _1707_ _0116_ _0174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_221_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2765__A2 _1479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2879_ _1574_ _1914_ _0098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_135_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3714__A1 _0994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_219_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_173_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2910__S _1733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_218_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_236_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2156__I _1257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3641__B1 _1678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_244_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3851_ _1485_ _1115_ _1120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_149_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2802_ _1185_ _1705_ _1903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_32_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3782_ _1050_ _1036_ _1005_ _1063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_185_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_160_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2733_ _1833_ _1750_ _1834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_121_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2664_ _1715_ _1765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_173_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2595_ _1680_ _1695_ _1696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_236_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_140_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3216_ _0464_ _0465_ _0468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_228_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3147_ _0359_ _0362_ _0391_ _0392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__2683__A1 _1782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3078_ _0311_ _0315_ _0317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2029_ dsynth.freeRunCntr\[16\] _1131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_184_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_219_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2685__B _1577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2674__A1 _1338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2674__B2 _1364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2426__A1 _1516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3874__CLK net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_214_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_237_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2380_ dsynth.freeRunCntr\[32\] _1481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2901__A2 _1902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_232_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3001_ _0071_ _0076_ _0232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xinput6 io_in[22] net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XTAP_5080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2665__A1 _1547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3834_ _0536_ _0085_ _1574_ _1101_ _1107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_220_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3765_ _1045_ _1041_ _1046_ _1047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2716_ _1668_ _1817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_118_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3696_ _0974_ _0979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2647_ _1746_ _1747_ _1748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_133_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2578_ _1137_ _1491_ _1679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2656__A1 _1538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_216_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2120__A3 _1214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2408__A1 _1503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_145_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2959__A2 _1492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_212_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3384__A2 _0612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_183_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2344__B1 _1444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2895__A1 _1363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3072__A1 _1338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3550_ _0831_ _0835_ _0836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3375__A2 _0642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2501_ _1400_ _1599_ _1600_ _1601_ _1217_ _1602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
X_3481_ _0615_ _0753_ _0760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_127_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2432_ _1001_ _1533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2363_ _1445_ _1465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2886__A1 _1323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2294_ _0558_ _0184_ _1396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_81_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout32_I net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2810__A1 _1207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_221_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3817_ _1090_ _1091_ _1094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_222_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3748_ _1028_ _1029_ _1031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3679_ tmux.clkpab _0964_ tmux.clkbpb vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_133_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_87_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_210_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xuser_proj_example_104 la_data_out[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_115 la_data_out[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_71_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_example_126 la_data_out[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_109_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_example_137 la_data_out[39] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_148 la_data_out[50] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_137_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_proj_example_159 la_data_out[61] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_109_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3109__A2 _1492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_238_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2868__A1 _1615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2096__A2 _1197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_234_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2981_ _0208_ _0209_ _0210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_128_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2164__I _1265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3596__A2 _0696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1932_ _0184_ _0195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_226_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3602_ _0856_ _0892_ _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_190_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3533_ _0807_ _0808_ _0816_ _0817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_115_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3464_ _0721_ _0722_ _0741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2415_ _0096_ _1516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_217_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3395_ _0655_ _0654_ _0656_ _0664_ _0665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_170_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2346_ _1417_ _1416_ _1447_ _1448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_69_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2323__A3 _1302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_244_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2277_ _0118_ _1378_ _1379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_244_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3284__A1 _1429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2074__I _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_244_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_224_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3339__A2 _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_146_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_192_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2249__I _1146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_189_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_223_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_145_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2250__A2 _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_171_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2200_ _1219_ _0514_ _1213_ _1302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3502__A2 _1817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3180_ _0406_ _0423_ _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_234_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2131_ dsynth.freeRunCntr\[10\] _1233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_226_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2062_ _0855_ _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_93_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_240_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3018__A1 _1364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2964_ _0172_ _0174_ _0190_ _0191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_245_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2895_ _1363_ _1504_ _0115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_124_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3516_ _0793_ _0797_ _0798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_103_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3447_ _0718_ _0719_ _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_213_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3378_ _1340_ _0647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2329_ _1419_ _1430_ _1431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_3507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input12_I io_in[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_232_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2480__A2 _1580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_214_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_167_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3732__A2 _1006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_175_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_191_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_6188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3248__A1 _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_210_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_203_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3420__A1 _1464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2680_ _1764_ _1770_ _1781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_157_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2526__A3 _1626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3301_ _0268_ _0542_ _0561_ _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_173_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3232_ _1415_ _0351_ _0486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xuser_proj_example_68 io_oeb[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA_input4_I io_in[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xuser_proj_example_79 io_out[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_214_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3163_ _0380_ _0381_ _0410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_227_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2114_ _1211_ _1215_ _0963_ _1216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3094_ _0296_ _0300_ _0301_ _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_243_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2045_ _0239_ _1146_ _0690_ _1147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_78_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2462__A2 _1562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout39 net46 net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_206_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3411__A1 _1385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2947_ _1715_ _0170_ _0171_ _0172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_143_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3411__B2 _1463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_198_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2878_ _1642_ _1851_ _1732_ _0097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_30_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3714__A2 _0996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_219_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3478__A1 _1834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_198_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2453__A2 _1553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_213_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2262__I _1363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_221_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_1746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_225_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2444__A2 _1485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3641__A1 _1233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3641__B2 _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3850_ _1485_ _1116_ _1119_ _0024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_207_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2801_ _1481_ _1478_ _1902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_3781_ _1062_ _0003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_13_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2732_ _1699_ _1833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_199_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2663_ _1679_ _1763_ _1764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_117_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2594_ _1682_ _1694_ _1695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_160_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3215_ _0252_ _0453_ _0467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_45_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3146_ _0376_ _0390_ _0391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_94_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3077_ _0291_ _0314_ _0315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_83_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2028_ _1123_ _1129_ _1095_ _1103_ _1130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_110_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2435__A2 _1534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3632__A1 _1463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_219_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2123__A1 _1218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_213_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_207_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2674__A2 _1666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3623__A1 _1131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_201_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_204_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3387__B1 _0654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2114__A1 _1211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3000_ _0230_ _0231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_7_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput7 io_in[25] net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2665__A2 _1544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3090__A2 _0329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3833_ _0112_ _1104_ _1106_ _0017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_123_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3764_ dsynth.freeRunCntr\[9\] _1027_ _1038_ _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_9_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_203_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2715_ _1672_ _1697_ _1815_ _1816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3695_ net8 _0978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_173_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2646_ _1512_ _1660_ _1747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_195_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_236_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2577_ _1677_ _1678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_210_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3129_ _0366_ _0372_ _0373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3605__A1 _1465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2408__A2 _1506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_184_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2344__A1 _1419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_219_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2344__B2 _1445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_234_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2895__A2 _1504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3844__A1 _1477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2583__A1 _1683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2500_ _0459_ _1331_ _1270_ _0931_ _1601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_3480_ _0758_ _0643_ _0759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2431_ _1531_ _1532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_237_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2335__A1 _1404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2362_ _1463_ _1464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2886__A2 _1403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2293_ _1394_ _1277_ _1327_ _1367_ _0206_ _1395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_237_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_209_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_220_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2810__A2 _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_165_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3816_ _1157_ _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3747_ dsynth.freeRunCntr\[8\] _1019_ _0970_ _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_192_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3678_ net6 _0964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_137_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2629_ _1001_ _1690_ _1730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_192_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2326__A1 _1030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3864__CLK net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_153_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_216_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_212_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_211_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xuser_proj_example_105 la_data_out[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_116 la_data_out[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_184_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_proj_example_127 la_data_out[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_138 la_data_out[40] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_149 la_data_out[51] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_164_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2203__C _1069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2868__A2 _1706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3045__A2 _0279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2980_ _0128_ _0136_ _0209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1931_ _0173_ _0184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_159_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_187_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_238_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput10 io_in[28] net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3601_ _0857_ _0859_ _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_204_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2556__A1 _1640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3887__CLK net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3532_ _0815_ _0773_ _0779_ _0816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_196_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3463_ _0717_ _0725_ _0740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2308__A1 _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2414_ _1514_ _1515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3394_ _1461_ _0658_ _0663_ _1451_ _0664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_135_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2345_ _1431_ _1446_ _1447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_233_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2276_ _1371_ _1373_ _1376_ _1377_ _1378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_111_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_42_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3284__A2 _0249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_240_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_244_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_189_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_19_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_199_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_11_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_199_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3096__I _0098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2538__A1 _1634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_197_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3502__A3 _0730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2130_ _1230_ _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_66_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2061_ _1162_ _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_234_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3018__A2 _0249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2963_ _0188_ _0189_ _0190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_222_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2777__A1 _1609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2894_ _0111_ _0113_ _0114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3515_ _0795_ _0796_ _0797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_200_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3446_ _0991_ _1817_ _0395_ _1186_ _0721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_143_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3377_ _1459_ _0644_ _0645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2328_ _1429_ _1430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_230_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2259_ _1353_ _1356_ _1359_ _1320_ _1360_ _1361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XTAP_2807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_207_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_228_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2768__A1 _1864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2940__A1 _1381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_216_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_245_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2471__A3 _1571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_232_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_160_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_242_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_117_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3300_ _0491_ _0543_ _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_140_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3231_ _0483_ _0484_ _0485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xuser_proj_example_69 io_oeb[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_100_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3162_ _0376_ _0390_ _0408_ _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2113_ _1212_ _1214_ _1215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3093_ _0300_ _0301_ _0296_ _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_236_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2044_ _1144_ _1145_ _1146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_208_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2998__A1 _0160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_235_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_245_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2633__I _1733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2946_ _1548_ _0045_ _1653_ _0171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_17_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2877_ _0084_ _0088_ _0094_ _0095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_191_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3429_ _0702_ _1549_ _1597_ _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_213_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_241_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3890__RN net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_224_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_181_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3166__A1 _1428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_237_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2913__A1 _1635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_237_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_235_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3641__A2 _1683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2800_ _1865_ _1899_ _1900_ _1901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3881__RN net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3780_ _1057_ _1061_ _1062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_203_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2731_ _1811_ _1831_ _1832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_140_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2662_ _1616_ _1761_ _1762_ _1763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_172_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3157__A1 _1430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_246_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_161_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2593_ _1684_ _1693_ _1694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_160_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3214_ _0464_ _0465_ _0466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_227_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_214_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3145_ _0378_ _0389_ _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_243_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout55_I net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3076_ _1707_ _0313_ _0314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_209_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2027_ _1128_ _1129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_208_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3632__A2 _0489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_211_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2363__I _1445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3872__RN net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2929_ _0042_ _0067_ _0153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_108_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_164_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3623__A2 _1681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2682__I0 _1732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2831__B1 _0045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3387__A1 _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_204_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3387__B2 _0655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3139__A1 _0090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3139__B2 _0175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_233_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_209_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput8 io_in[26] net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_5082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_225_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_221_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_162_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3832_ _1132_ _1104_ _1106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_18_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3763_ _1027_ _1038_ dsynth.freeRunCntr\[9\] _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2714_ _1674_ _1696_ _1815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_3694_ _0977_ _0011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2645_ _1712_ _1744_ _1745_ _1746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_133_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2889__B1 _1301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2576_ _1629_ _1677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_160_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3302__A1 _0276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3128_ _0367_ _0370_ _0372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_228_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3059_ _0282_ _1528_ _0279_ _0295_ _0267_ _0296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XANTENNA__3605__A2 _0689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2307__B _1370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_211_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2093__I _0701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_149_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2041__A1 _1141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2592__A2 _1692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_234_1728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2344__A2 _1430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2268__I _1212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_207_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_246_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_187_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_204_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2583__A2 _1532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2430_ _1530_ _1531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2361_ _1417_ _1463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_48_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3562__I dsynth.freeRunCntr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2292_ _1393_ _1394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_173_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3048__B1 _0185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_244_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_61_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2271__A1 _1125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2810__A3 _1244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3815_ _1092_ _0010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_177_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3737__I _0994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_203_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3746_ _1027_ _0970_ _1313_ _1028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_20_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3771__A1 _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3677_ _0962_ net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_173_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2628_ _1714_ _1715_ _1629_ _1685_ _1728_ _1617_ _1729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_66_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2326__A2 _1427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2559_ _1614_ _1659_ _1660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_5807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_178_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_221_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_proj_example_106 la_data_out[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_example_117 la_data_out[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_32_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_example_128 la_data_out[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_165_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_example_139 la_data_out[41] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__3762__A1 _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3382__I dsynth.freeRunCntr\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2500__B _0931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_234_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1930_ _0162_ _0173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_245_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3600_ _1232_ _0865_ _0874_ _0889_ _0890_ _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
Xinput11 io_in[35] net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_200_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2556__A2 _1642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3531_ _0812_ _0813_ _0814_ _0769_ _0815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_122_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3462_ _0726_ _0738_ _0739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_143_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2308__A2 _1282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2413_ _1513_ _1476_ _1473_ _1514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_174_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3393_ _0082_ _0649_ _0663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_83_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2344_ _1419_ _1430_ _1444_ _1445_ _1446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_229_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2275_ _1292_ _1329_ _1291_ _1377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_226_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2492__A1 _1576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_225_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2619__I0 _1150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_209_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2244__A1 _1141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_224_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2547__A2 _0228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3729_ _0987_ _1011_ _1012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_244_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_216_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2483__A1 _1516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_231_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_244_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_164_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_196_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_106_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_200_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3035__I0 _0131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2538__A2 _1635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_201_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2060_ _0822_ _0734_ _1162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_240_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_235_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_207_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2962_ _1707_ _0116_ _0172_ _0189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_15_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_206_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_241_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2893_ _0104_ _0110_ _0112_ _0113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_147_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3726__A1 _0655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3514_ _0726_ _0738_ _0796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_239_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3445_ _0718_ _0719_ _0720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3376_ _0617_ _0643_ _0644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2327_ _1428_ _1429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_170_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2258_ _0958_ _1360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_2_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2189_ _1235_ _1291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_246_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_240_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2768__A2 _1865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_223_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3717__A1 _1417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_68_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2153__B1 _1224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_89_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3660__I net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_194_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_4700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2456__A1 _1555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_244_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3877__CLK net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_205_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_197_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2225__B _1239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_158_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3230_ _0398_ _0392_ _0397_ _0484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_98_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3161_ _0378_ _0389_ _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2112_ _1213_ _1214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_212_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3092_ _0309_ _0317_ _0331_ _0332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_5990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2043_ _0250_ _1145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_81_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2945_ _0111_ _0113_ _0170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_56_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2876_ _0092_ _0093_ _0094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_148_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_209_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3428_ _1584_ _0702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3478__A3 _0642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3359_ _1823_ _1825_ _0626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_189_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2438__A1 _1274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_245_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2438__B2 _1538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3635__B1 _1544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_226_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2045__B _0690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2610__A1 _1312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3166__A2 _1667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_207_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_204_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2730_ _1814_ _1816_ _1830_ _1831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_220_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2661_ _1286_ _1500_ _1762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_195_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3157__A2 _0402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2592_ _1686_ _1692_ _1693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_154_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_119_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3213_ _0264_ _0263_ _0465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2668__A1 _1503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3144_ _0383_ _0388_ _0389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_228_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3075_ _1311_ _0312_ _0252_ _0313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_227_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2026_ _1127_ _1128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_fanout48_I net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_224_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2928_ _0148_ _0149_ _0150_ _0152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_206_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2859_ _0073_ _0075_ _0076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_3_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2123__A3 _1224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_227_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_157_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2682__I1 _1730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2831__B2 _1532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_202_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2347__B1 _1381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_235_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput9 io_in[27] net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_5083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2822__A1 _0035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_233_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3831_ _1105_ _0016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_221_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3762_ _0873_ _1043_ _1044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2425__I1 _1525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2713_ _1663_ _1812_ _1813_ _1814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3693_ _0973_ _0976_ _0977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_145_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2644_ _1742_ _1743_ _1745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_161_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2338__B1 _1258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2889__A1 _1331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2575_ _1675_ _1676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__2889__B2 _1389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_236_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_214_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3127_ _0368_ _0369_ _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_27_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3058_ _0114_ _0295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_167_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_227_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2009_ _1010_ _1020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_149_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2307__C _1179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_234_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3057__B2 _0277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_221_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_128_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2233__B _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_204_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2360_ _1461_ _1339_ _1365_ _1451_ _1418_ _1462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_233_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2740__B1 _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2291_ _1374_ _1242_ _1393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3296__A1 _0452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3048__A1 _0282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3048__B2 _1549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_213_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_209_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3814_ _1090_ _1091_ _1092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_193_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3745_ _1019_ _1027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_158_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3676_ net43 tmux.clkpab net5 tmux.clkpbb _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_118_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2627_ _1727_ _1728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_133_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2558_ _1632_ _1658_ _1659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_99_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2369__I _1470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_1740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2489_ _1589_ _1590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3287__A1 _0452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3039__A1 _0265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_244_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_223_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xuser_proj_example_107 la_data_out[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_109_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_example_118 la_data_out[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_123_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xuser_proj_example_129 la_data_out[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_197_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_178_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_228_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2005__A2 _0971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput12 io_in[36] net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_168_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3530_ _0766_ _0814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_176_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3461_ _0727_ _0737_ _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_170_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2412_ dsynth.freeRunCntr\[30\] _1513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_100_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3392_ _1459_ _0644_ _0658_ _1461_ _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_48_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2189__I _1235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2343_ dsynth.freeRunCntr\[1\] _1445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_170_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2274_ _1207_ _1369_ _1375_ _1376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_42_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2492__A2 _1581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_226_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2619__I1 _1251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3044__I1 _0170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1989_ _0217_ _0822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_14_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3728_ _1004_ _0979_ _1011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_179_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3659_ _0951_ _0953_ net15 net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_161_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2099__I _1200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_229_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2483__A2 _1583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_243_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_43_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3432__A1 _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3658__I net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_237_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1994__A1 _0844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3035__I1 _0130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_240_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_193_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_234_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2171__A1 _1270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_226_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2474__A2 _1571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2961_ _0175_ _0187_ _0188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_43_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_143_1737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2892_ _1516_ _0112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3726__A2 _1006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3513_ _0794_ _0737_ _0795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_171_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3444_ _0709_ _0714_ _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_83_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3375_ _0619_ _0642_ _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2326_ _1030_ _1427_ _1428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_230_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2257_ _1357_ _1358_ _1359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_22_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2188_ dsynth.freeRunCntr\[9\] _1290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_225_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3662__A1 _0954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_214_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_20_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3414__A1 _0587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_209_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_33_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3717__A2 _0989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2153__A1 _1214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2153__B2 _1205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_237_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_90_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2456__A2 _1294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2208__A2 _1309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2292__I _1393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_214_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3160_ _0374_ _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_136_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2111_ _0371_ _1213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3091_ _0293_ _0308_ _0331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_5980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2042_ dsynth.csTable.address\[1\] _1144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_66_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_207_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_206_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2944_ _0161_ _0165_ _0168_ _0169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_241_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_176_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2875_ _0084_ _0088_ _0093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_175_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2151__B _1192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1990__B _0822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3427_ _1596_ _1685_ _1824_ _0623_ _0699_ _1576_ _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_217_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3358_ _1702_ _1863_ _1640_ _0623_ _1503_ _0625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XTAP_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2309_ _1218_ _1411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_58_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3289_ _0489_ _0268_ _0542_ _0548_ _0549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_3318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input10_I io_in[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2438__A2 _1150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3635__A1 dsynth.freeRunCntr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3635__B2 _1313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2610__A2 _1700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_237_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3626__A1 _1118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_207_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2750__I _1761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2660_ _1759_ _1760_ _1761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2591_ _1687_ _1691_ _1692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2365__A1 _1464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3212_ _0461_ _0462_ _0463_ _0267_ _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_140_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input2_I io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2912__I0 _0055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3143_ _0384_ _0387_ _0388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_94_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3074_ _1310_ _1504_ _0312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_67_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3617__A1 _1465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2025_ _1124_ _1126_ _1127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_36_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2927_ _0146_ _0147_ _0150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2858_ _0069_ _0070_ _0075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_108_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2789_ _1887_ _1888_ _1890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__2356__A1 _1290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3867__CLK net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2659__A2 _1758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2831__A2 _0033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2347__A1 dsynth.freeRunCntr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2347__B2 _1382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2898__A2 _1917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_237_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3847__A1 _1486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_162_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_188_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_244_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_232_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3830_ _0085_ _1104_ _1105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_127_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3761_ _1021_ _0967_ _0980_ _1043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_105_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2712_ _1665_ _1671_ _1813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3692_ dsynth.freeRunCntr\[1\] _0975_ _0976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_146_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2643_ _1742_ _1743_ _1744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__2338__A1 _1224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2574_ _1490_ _1675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__2889__A2 _1202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_228_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3126_ _1399_ _1675_ _0369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_151_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3057_ _0281_ _0291_ _0292_ _0280_ _0277_ _0293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__3066__A2 _0114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_224_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2008_ _0085_ _1001_ _1010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_145_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2329__A1 _1419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_232_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2501__A1 _1400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_219_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2565__I _1479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3057__A2 _0291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2804__A2 _1902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_159_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2568__A1 _1486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2233__C _1334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2740__A1 _0668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2740__B2 _1270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2290_ _1323_ _1243_ _1354_ _1392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_81_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3048__A2 _1678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_206_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_233_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_221_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3813_ _1145_ dsynth.freeRunCntr\[17\] _1085_ _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_14_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3744_ _1026_ _0030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3675_ net11 _0955_ net1 net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_118_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2626_ _1725_ _1726_ _1727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2557_ _1639_ _1657_ _1658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_153_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2488_ _1513_ _1474_ _1471_ _1589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_25_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_214_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_233_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3109_ _0089_ _1492_ _0351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3039__A2 _0270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_proj_example_108 la_data_out[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_71_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3211__A2 _0336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xuser_proj_example_119 la_data_out[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_137_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2970__A1 _1630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2722__A1 _1640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2228__C _0963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_147_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput13 io_in[37] net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_122_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_204_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2961__A1 _0175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3460_ _0732_ _0736_ _0737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_155_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_157_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_217_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2411_ _1496_ _1510_ _1512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_3391_ _1314_ _0644_ _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_87_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2342_ _1443_ _1444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_96_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2273_ _1374_ _1237_ _1344_ _1223_ _1375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_215_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_197_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_193_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1988_ _0437_ _0811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3727_ _1009_ _0028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2952__A1 _1241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3658_ net14 _0953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_164_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2609_ _1498_ _1509_ _1710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_162_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3589_ dsynth.freeRunCntr\[10\] _0876_ _0878_ _0879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_6318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_192_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3680__A2 net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_244_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3432__A2 _0704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_223_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_240_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_19_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2491__I0 _1586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_11_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2171__A2 _1257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_234_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2960_ _1514_ _0185_ _0186_ _0187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2891_ _1636_ _0104_ _0110_ _0111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_179_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_230_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3512_ _0727_ _0794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_176_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3443_ _1823_ _1825_ _0629_ _0630_ _0625_ _0718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_100_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3374_ _0638_ _0641_ _0642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2325_ _1411_ _1423_ _1426_ _1427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2256_ _1220_ _1246_ _1167_ _1358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_239_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3111__A1 _1762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2187_ _1233_ _1266_ _1287_ _1288_ _1289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_168_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3662__A2 net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_226_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_240_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3178__A1 _1430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2153__A2 _1243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_235_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3102__A1 _1734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3893__RN net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_160_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_212_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_32_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_240_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_193_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_239_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3341__A1 _1381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2110_ _1059_ _1212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3090_ _0325_ _0329_ _0330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_5970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_181_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2041_ _1141_ _1142_ _1143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_47_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3579__I _1230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_222_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3884__RN net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2943_ _0166_ _0167_ _0168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_175_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2080__A1 _0206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2874_ _0091_ _0092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_198_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3528__B _0753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2907__A1 _0100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3426_ _1857_ _0699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_98_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3357_ _1617_ _0623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_246_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2308_ _1253_ _1282_ _1410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3288_ _0336_ _0276_ _0266_ _0548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_189_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2239_ _1313_ _1312_ _1339_ _1340_ _1341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_96_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3635__A2 _1528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_241_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_227_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_241_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3875__RN net58 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2071__A1 _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_237_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_159_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3626__A2 _0702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_233_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3866__RN net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_199_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2590_ _1636_ _1690_ _1691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_172_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2365__A2 _1416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3211_ _0266_ _0336_ _0260_ _0463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_214_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3142_ _0385_ _0386_ _0387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_6490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_227_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3073_ _0175_ _0253_ _0310_ _0311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_94_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3617__A2 _0518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2024_ _1125_ _0800_ _1126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_209_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_223_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_225_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2926_ _0095_ _0124_ _0149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_176_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2857_ _1906_ _0041_ _0072_ _0073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_108_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2788_ _1887_ _1888_ _1889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_191_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2356__A2 _1287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3305__A1 _0306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3409_ _0235_ _0680_ _0681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_154_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_196_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2347__A2 _1399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2898__A3 _0100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_162_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_131_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_221_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_207_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2035__A1 _1010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3760_ _1042_ _0032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3783__A1 _1136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2711_ _1665_ _1671_ _1812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_185_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3691_ net8 _0974_ net9 net10 _0975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_9_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2642_ _1568_ _1612_ _1743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_145_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2338__A2 _1205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2573_ _1632_ _1658_ _1673_ _1674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_113_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_236_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3125_ _1265_ _1704_ _1664_ _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_3_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout53_I net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3056_ _0284_ _0285_ _0292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_64_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2007_ dsynth.csTable.address\[7\] _1001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2274__A1 _1207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_227_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_184_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_221_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2909_ _1759_ _1760_ _0131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_3889_ _0019_ net49 net33 dsynth.freeRunCntr\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_109_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2329__A2 _1430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3435__C _1498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_234_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2067__B _1161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2265__A1 _1245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_226_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_230_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2017__A1 _1030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1925__I _0107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_237_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2740__A2 _1258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_238_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3361__B _1852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2756__I _1765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_237_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2256__A1 _1220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3857__CLK net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_244_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_220_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3812_ _1144_ _1090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_159_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3743_ _0647_ _1023_ _1025_ _1026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_203_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3674_ _0955_ _0959_ net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_173_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3508__A1 _0728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2625_ _1633_ _1721_ _1724_ _1726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_12_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2556_ _1640_ _1642_ _1654_ _1656_ _1657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_142_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_1731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2487_ _1572_ _1575_ _1587_ _1588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_141_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_228_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2495__A1 _1569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3108_ _0303_ _0304_ _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3039_ _0265_ _0270_ _0274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_37_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_example_109 la_data_out[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_20_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2970__A2 _0170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2722__A2 _1765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2576__I _1629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_219_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_235_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2789__A2 _1888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput14 io_in[5] net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_128_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_196_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2410_ _1497_ _1510_ _1511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3390_ _0645_ _0659_ _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_108_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2341_ _1030_ _1442_ _1443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_96_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2272_ _0888_ _1374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2229__A1 _1141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_222_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1987_ _0668_ _0701_ _0767_ _0789_ _0800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_33_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3726_ _0655_ _1006_ _1008_ _1009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_119_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_174_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3657_ net11 _0951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_106_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2608_ _1702_ _1704_ _1708_ _1503_ _1709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_161_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3588_ _0869_ _0870_ _0875_ _0878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_6308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2539_ _1607_ _1608_ _1640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_5607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_217_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3432__A3 _0705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_197_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_240_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_137_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3690__I net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_143_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2890_ _1411_ _0106_ _0108_ _1283_ _0109_ _1194_ _0110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XTAP_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_147_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_204_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3511_ _0788_ _0792_ _0793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_128_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3442_ _0706_ _0716_ _0717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_170_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3373_ _1814_ _0639_ _0640_ _0641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2324_ _1349_ _1199_ _1424_ _1425_ _1260_ _1426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XTAP_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2255_ _1175_ _1246_ _1357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_111_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2186_ dsynth.freeRunCntr\[9\] _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3662__A3 net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_228_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2622__A1 _0958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_240_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3178__A2 _0402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3709_ _1464_ _0989_ _0992_ _0993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_134_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_89_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_192_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_216_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_207_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3685__I net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_149_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2129__B1 _1229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1933__I _0195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3341__A2 _0402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_234_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2040_ _0712_ _1142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_5993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_235_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2942_ _0161_ _0165_ _0167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_222_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2080__A2 _1174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2873_ _0090_ _1902_ _0091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_191_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3425_ _0697_ _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_213_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3356_ _1821_ _1827_ _0621_ _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2307_ _1250_ _1252_ _1370_ _1179_ _1409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_189_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3287_ _0452_ _0545_ _0546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2238_ dsynth.freeRunCntr\[7\] _1340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2169_ _0679_ _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3323__A2 _0585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_192_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3087__A1 _1443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2584__I _1642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2834__A1 _0048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3890__CLK net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_198_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_203_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1928__I dsynth.csTable.address\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_158_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3210_ _0266_ _1848_ _0462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3141_ _1762_ _0187_ _0386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_6480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3072_ _1338_ _0241_ _0310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_5790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2023_ _0580_ _1125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_208_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3250__A1 _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2925_ _0146_ _0147_ _0148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_143_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_225_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2856_ _0039_ _0040_ _0072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_15_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2787_ _1781_ _1796_ _1888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_116_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_236_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3408_ _0231_ _0677_ _0678_ _0680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_172_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3339_ _0599_ _0603_ _0604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3069__A1 _0303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2816__A1 _1514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_227_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2667__I1 _1702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_198_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_164_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3241__A1 _0489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_110_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_225_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2807__A1 _1389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2035__A2 _0971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3232__A1 _1415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2710_ _1810_ _1811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_199_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3783__A2 _1063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3690_ net7 _0974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_158_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_145_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2641_ _1729_ _1740_ _1741_ _1742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_12_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2572_ _1639_ _1657_ _1673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_114_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3124_ _0326_ _0328_ _0367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_23_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_215_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3055_ _0284_ _0285_ _0291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_209_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2006_ _0981_ _0991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_227_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_fanout46_I net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2908_ _1759_ _1760_ _1587_ _0130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_137_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3888_ _0018_ net49 net33 dsynth.freeRunCntr\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2839_ _0053_ _0054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_178_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_236_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_207_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3023__I _1676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_187_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3214__A1 _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2017__A2 _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_204_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_233_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_215_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2256__A2 _1246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3453__A1 _1128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_221_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_181_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3811_ _1089_ _0009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3205__A1 _1838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3742_ _1014_ _1017_ _1024_ _1025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_174_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_173_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3673_ _0959_ _0961_ net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_179_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2624_ _1721_ _1724_ _1569_ _1725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2555_ _1638_ _1655_ _1656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_192_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2486_ _1578_ _1587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_141_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3044__S _0054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_210_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2495__A2 _1595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_244_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3107_ _1838_ _0347_ _0313_ _1704_ _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_186_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3038_ _0186_ _0246_ _0273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_110_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_221_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2183__A1 _1235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_219_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_234_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3435__A1 _1128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2806__B _1211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput15 io_in[6] net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1936__I _0228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2410__A2 _1510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_217_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_174_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2340_ _1435_ _1437_ _1441_ _1404_ _1442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_123_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2271_ _1125_ _1372_ _1373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_46_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_237_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3029__I1 _0131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1986_ _0778_ _0789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3725_ _0998_ _1002_ _1007_ _1008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_20_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3656_ _0927_ _0938_ _0950_ net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_173_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2607_ _1706_ _1707_ _1708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_192_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3587_ _0875_ _0869_ _0870_ _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__2165__A1 _1233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2538_ _1634_ _1635_ _1610_ _1638_ _1639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_216_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2469_ _1354_ _0833_ _1161_ _1570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_4907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3665__A1 net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_243_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_232_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3417__A1 _0672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_227_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_244_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_164_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_196_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_106_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_240_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2080__C _0963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_234_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2459__A2 _1555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_219_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3510_ _0790_ _0791_ _0792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_89_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3441_ _0709_ _0714_ _0715_ _0716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_170_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2147__A1 _1241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3372_ _1816_ _1830_ _0640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_170_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2323_ _1404_ _0767_ _1302_ _1425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_112_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2254_ _1354_ _0767_ _1247_ _1355_ _1356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__3647__A1 _0684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2185_ _1286_ _1287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_66_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_225_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_214_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_221_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2622__A2 _1206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2181__B _0931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1969_ dsynth.csTable.address\[6\] dsynth.csTable.address\[1\] _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_198_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2386__A1 _1486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3708_ _0983_ _0985_ _0990_ _0992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_174_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3639_ _0868_ _1640_ _0707_ _0698_ _0933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_108_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2138__A1 _1239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_235_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_157_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3350__A3 _0612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_89_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3638__A1 _0647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_217_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_213_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_197_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_235_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_193_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_197_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2129__A1 dsynth.freeRunCntr\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2129__B2 _1230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2110__I _1059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2266__B _1166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2941_ _1415_ _1666_ _0166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2604__A2 _1491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_203_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2872_ _0089_ _0090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_176_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3097__B _1635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_223_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3317__B1 _0539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3424_ dsynth.freeRunCntr\[12\] _0697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_171_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3355_ _1822_ _1826_ _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_48_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2306_ _1143_ _1194_ _1407_ _1408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3286_ _1429_ _0542_ _0544_ _0545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_246_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2237_ _1338_ _1339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_72_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_241_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2168_ _1223_ _1270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_187_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2099_ _1200_ _1201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_228_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_179_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_5213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2531__A1 _1615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3087__A2 _1666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_244_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2834__A2 _1527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2105__I _1206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2522__A1 _1143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3140_ _0337_ _0339_ _0385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_6470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3071_ _0293_ _0308_ _0309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_5780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2022_ _0107_ _1124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_235_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_224_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2724__B _1782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_245_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2589__A1 _0920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2924_ _0043_ _0062_ _0147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_182_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2855_ _0069_ _0070_ _0071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_206_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2786_ _1874_ _1885_ _1886_ _1887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2761__A1 _1860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_236_1730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_236_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3407_ _0158_ _0229_ _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_193_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3338_ _0431_ _0600_ _0601_ _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3069__A2 _0306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3269_ _0526_ _0304_ _0527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_246_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2816__A2 _1915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2752__A1 _1527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_163_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2504__A1 _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_172_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2809__B _1360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2807__A2 _1394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2544__B _1644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_242_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3232__A2 _0351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_203_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_186_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2640_ _1738_ _1739_ _1741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2571_ _1663_ _1665_ _1671_ _1672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_126_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_206_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3123_ _1428_ _1667_ _0366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_110_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2259__B1 _1359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3054_ _0287_ _0288_ _0289_ _0290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_208_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2005_ _0118_ _0971_ _0981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_188_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2274__A3 _1375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout39_I net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_223_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_225_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2907_ _0100_ _0127_ _0128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3887_ _0017_ net51 net35 dsynth.csTable.address\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_176_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2838_ _1725_ _1726_ _1587_ _0053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_136_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2769_ _1860_ _1861_ _1870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2734__A1 _1834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3880__CLK net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_232_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_230_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_227_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_159_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_186_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_199_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_148_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_243_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2973__A1 _1587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2811__C _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3453__A2 _1668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3810_ _1145_ _1088_ _1089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_177_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3205__A2 _1493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3741_ _0651_ _1019_ _1012_ _1024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_158_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2964__A1 _0172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_201_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3672_ net3 net4 net11 net2 _0961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_31_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2623_ _1161_ _1722_ _1723_ _0404_ _1724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_220_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2554_ _1651_ _1655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2485_ _1572_ _1575_ _1586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_233_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3141__A1 _1762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3106_ _1338_ _0249_ _0347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_231_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3037_ _0265_ _0270_ _0271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_149_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3747__A3 _0970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2955__A1 _1553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2955__B2 _1644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_178_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_210_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2806__C _1393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3435__A2 _0256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_204_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_167_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_239_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3209__I _1915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_217_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2270_ _1301_ _1258_ _1272_ _1202_ _1372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_26_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2269__B _1370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3123__A1 _1428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_226_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1985_ _0173_ _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_193_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2937__A1 _1265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3724_ _0905_ _0994_ _0996_ _1007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_228_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_179_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3655_ _0915_ _0940_ _0924_ _0949_ _0950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_162_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2606_ _1703_ _1707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_3586_ _0814_ _0875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_66_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2165__A2 _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2537_ _1580_ _1637_ _1638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_114_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_192_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2468_ _1533_ _1569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3114__A1 _0346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2399_ _1477_ _1499_ _1500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_197_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_224_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_223_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_244_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_205_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3353__A1 _1834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_234_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_182_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3592__A1 _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2395__A2 _1495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_200_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3440_ _0710_ _0713_ _0715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_100_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3371_ _1816_ _1830_ _0639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_83_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2322_ _1345_ _1403_ _1148_ _1424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2253_ _0789_ _1355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_214_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3647__A2 _0295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_230_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2184_ _1010_ _1285_ _1286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_187_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3887__RN net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2018__I dsynth.freeRunCntr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_206_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_209_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2622__A3 _1402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2462__B _1516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1968_ _0470_ _0525_ _0580_ _0591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_119_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3707_ _1419_ _0982_ _0990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_88_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3638_ _0647_ _1714_ _0929_ _0930_ _0932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__2138__A2 _1146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_108_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3569_ _1136_ _0841_ _0847_ _0857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_103_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3638__A2 _1714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3878__RN net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_232_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2356__C _1139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_227_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_231_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_207_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_164_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_169_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2377__A2 _1477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3326__A1 _0160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2129__A2 _1186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_234_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_181_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_181_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_235_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3869__RN net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2940_ _1381_ _1490_ _0164_ _0165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_188_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_206_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2871_ _1020_ _1398_ _0089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_128_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3565__A1 _0832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2368__A2 _1469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3423_ _0661_ _0662_ _0665_ _0695_ _0696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_132_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2301__I _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_217_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_119_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3354_ _1186_ _1817_ _0395_ _1229_ _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_225_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2305_ _1406_ _1301_ _1358_ _1407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3285_ _0245_ _0543_ _0544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2236_ _1337_ _1338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_241_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2457__B _1556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_230_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2167_ _1232_ _1229_ _1231_ _1268_ _1269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_214_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2098_ _1151_ _1200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_213_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_210_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_235_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_89_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2531__A2 _1631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2295__A1 _1360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2295__B2 _1396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3547__A1 _1681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_180_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2522__A2 _1346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1960__I _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3070_ _0296_ _0302_ _0307_ _0308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XTAP_5770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2021_ _1118_ _1123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_188_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2286__A1 _1218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2589__A2 _1644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2923_ _0142_ _0143_ _0145_ _0146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_147_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2854_ _1873_ _1889_ _0070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_34_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2785_ _1883_ _1884_ _1886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3406_ _0672_ _0673_ _0676_ _0610_ _0677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_113_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3571__B _1103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3337_ _0433_ _0442_ _0601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3268_ _0285_ _0526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2219_ _0448_ _1321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3199_ _0401_ _0425_ _0449_ _0450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_38_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3746__B _1313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2752__A2 _1547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2504__A2 _1257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_162_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_232_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_201_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2116__I _1217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2570_ _1266_ _1668_ _1670_ _1287_ _1671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_154_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_177_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3122_ _0363_ _0354_ _0364_ _0365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_6290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_228_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2259__A1 _1353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3053_ _0275_ _0286_ _0289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_222_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2004_ _0415_ _0591_ _0952_ _0963_ _0971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_224_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3759__A1 _1290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2906_ _0097_ _0099_ _0127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3886_ _0016_ net52 net36 dsynth.csTable.address\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_149_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2470__B _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2837_ _1563_ _1565_ _0052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_136_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2768_ _1864_ _1865_ _1868_ _1869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2699_ _1798_ _1799_ _1800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_104_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2498__A1 _1298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_210_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_167_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_230_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_208_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2422__A1 _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_1733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2661__A1 _1286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_177_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3740_ _1019_ _1022_ _1023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_159_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3610__B1 _0901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2290__B _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3671_ _0959_ _0960_ net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_173_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2622_ _0958_ _1206_ _1402_ _1257_ _1723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_31_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2553_ _1597_ _1653_ _1654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2484_ _1579_ _1584_ _1585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_190_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3105_ _0335_ _0345_ _0346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_68_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout51_I net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3036_ _0267_ _0269_ _0270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_24_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2652__A1 _1244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_212_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2404__A1 _1227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_225_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3869_ _0030_ net56 net39 dsynth.freeRunCntr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_176_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_100_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2891__A1 _1636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_243_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_196_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2946__A2 _0045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3123__A2 _1667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_215_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2882__A1 _1506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2634__A1 _1732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3870__CLK net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1984_ _0756_ _0767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_140_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2937__A2 _1664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_222_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3723_ _0987_ _0967_ _1005_ _1006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_146_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2304__I _0470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_228_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3654_ _0947_ _0937_ _0933_ _0948_ _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_220_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2605_ _1705_ _1706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_196_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3585_ _0868_ _0863_ _0864_ _0871_ _0872_ _0873_ _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai33_1
XFILLER_157_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2536_ _1636_ _1595_ _1637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_115_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2570__B1 _1670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2467_ _1567_ _1568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_87_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2398_ dsynth.freeRunCntr\[31\] _1471_ _1499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_84_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2873__A1 _0090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_228_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2625__A1 _1633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3019_ _1916_ _0252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_77_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2923__B _0145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_184_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2616__A1 _1347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_234_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3893__CLK net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_179_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_230_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_221_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3370_ _0636_ _0637_ _0638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2321_ _1394_ _1420_ _1422_ _1366_ _1423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2252_ _1321_ _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2183_ _1235_ _1273_ _1278_ _1160_ _1284_ _1285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_93_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_226_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_230_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2607__A1 _1706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_240_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2743__B _1322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2622__A4 _1257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_222_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1967_ _0569_ _0580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3706_ _0987_ _0966_ _0988_ _0989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_120_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3637_ _1314_ _1544_ _0930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3568_ _0849_ _0850_ _0853_ _0854_ _0856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XTAP_6108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_89_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2519_ _1256_ _1342_ _1163_ _1620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_5407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_192_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3499_ _0779_ _0780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_5418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_116_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_229_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_229_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_207_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_160_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_212_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_32_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_137_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_158_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_181_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2119__I _0239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3262__A1 _0268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_200_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_204_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2870_ _0086_ _0087_ _0088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_182_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3014__A1 _1786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_198_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3422_ _0683_ _0693_ _0694_ _0695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3353_ _1834_ _1832_ _0618_ _0619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2304_ _0470_ _1406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_234_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3284_ _1429_ _0249_ _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_135_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2235_ _1188_ _1336_ _1337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_239_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3413__I _0684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2166_ _1187_ _1267_ _1268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_227_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2097_ _1198_ _1199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_241_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2999_ _0158_ _0229_ _0230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_33_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_222_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_172_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_192_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2819__A1 _1547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_204_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2047__A2 _0646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_246_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3795__A2 _1022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_199_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3547__A2 _1515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_201_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2522__A3 _1396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_227_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2020_ dsynth.freeRunCntr\[15\] _1118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_5793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_206_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2922_ _0137_ _0144_ _0141_ _0145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_149_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3786__A2 _1056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2853_ _0042_ _0067_ _0068_ _0069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_129_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2740__C _1206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2784_ _1883_ _1884_ _1885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_30_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3405_ _0674_ _0675_ _0676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_217_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3336_ _0433_ _0442_ _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_219_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3267_ _1415_ _0524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_41_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2218_ _0393_ _1316_ _1319_ _1320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_66_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2277__A2 _1378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_230_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3198_ _0427_ _0428_ _0447_ _0429_ _0449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_2408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2149_ _0613_ _0734_ _0360_ _1251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_1707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_89_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_5045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_162_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2892__I _1516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_221_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_207_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2841__B _0055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_220_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_236_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1951__A1 _0294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3672__B net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1971__I _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3121_ _0350_ _0353_ _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_6280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3052_ _0242_ _0255_ _0288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_5590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3456__A1 _0728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2003_ _0958_ _0963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_64_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2905_ _0095_ _0124_ _0125_ _0126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_176_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3885_ _0015_ net48 net32 dsynth.csTable.address\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_34_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2836_ _1878_ _0049_ _1785_ _0051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_164_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2767_ _1866_ _1867_ _1868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_191_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2698_ _1712_ _1744_ _1799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_104_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3319_ _0540_ _0577_ _0581_ _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_100_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3447__A1 _0718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_162_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_203_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2217__I _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_74_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_148_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2422__A2 _0239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_237_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_238_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2836__B _1785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2661__A2 _1500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2127__I _1228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3667__B net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1966__I _0558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3670_ net3 net4 net2 _0960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_158_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2621_ _1243_ _1150_ _1282_ _1538_ _1722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_173_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2552_ _1652_ _1653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_12_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2483_ _1516_ _1583_ _1584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_233_1724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3104_ _0340_ _0344_ _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_116_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2746__B _1574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3429__A1 _0702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_244_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3035_ _0131_ _0130_ _0268_ _0269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_71_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2101__B2 _1202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout44_I net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2652__A2 _1153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2404__A2 _1504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3868_ _0029_ net56 net40 dsynth.freeRunCntr\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_203_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2819_ _1547_ _0033_ _0034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3799_ _1079_ _0006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_152_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3380__A3 _0612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_219_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3668__A1 _0951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2340__B2 _1404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2656__B _1375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2891__A2 _0104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_246_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_41_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2628__C1 _1728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output25_I net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2159__A1 _0942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_174_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3659__A1 _0951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2331__A1 _1239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_237_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_226_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2882__A2 _1917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_206_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2634__A2 _1734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1983_ _0712_ _0745_ _0756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_186_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3722_ _1004_ _0979_ _1005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_158_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3653_ _0935_ _0934_ _0948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_200_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2604_ _1701_ _1491_ _1705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3584_ dsynth.freeRunCntr\[10\] _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_114_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2535_ _1564_ _1636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2570__A1 _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2570__B2 _1287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2466_ _1515_ _1528_ _1532_ _1544_ _1549_ _1566_ _1567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
XFILLER_157_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_229_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2397_ _1494_ _1498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2322__A1 _1345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2873__A2 _1902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3018_ _1364_ _0249_ _0251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2625__A2 _1721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_212_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_58_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3050__A2 _0284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_238_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_191_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_232_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_215_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2001__B1 _0920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2320_ _1215_ _1421_ _1422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2251_ _1352_ _1298_ _1195_ _1353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_215_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_230_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2182_ _1280_ _1283_ _1217_ _1284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_26_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3804__A1 _1131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2607__A2 _1707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1966_ _0558_ _0569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_159_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3705_ _0978_ _0968_ _0988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_146_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_174_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3636_ _0928_ _0929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_146_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3567_ dsynth.freeRunCntr\[16\] _1118_ _0854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_108_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2518_ _1142_ _1200_ _1166_ _1619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_102_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3498_ _0777_ _0779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_5408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2449_ _1176_ _1294_ _1550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_4707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_213_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2653__C _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_242_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_240_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_193_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_165_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3860__CLK net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_181_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_210_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_245_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1974__I _0646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3421_ _1385_ _0681_ _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3352_ _1811_ _1831_ _0618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_97_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2303_ _1402_ _1403_ _1404_ _1405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_174_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3283_ _0245_ _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2234_ _1125_ _1326_ _1330_ _1335_ _1336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_238_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2165_ _1233_ _1266_ _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2096_ _1196_ _1197_ _1198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2998_ _0160_ _0226_ _0227_ _0229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_72_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1949_ _0327_ _0338_ _0371_ _0382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_120_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2764__A1 _1137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3619_ _1382_ _0131_ _0911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_200_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3883__CLK net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2819__A2 _0033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2295__A3 _1353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3492__A2 _0642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_229_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_60_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_233_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_235_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2293__C _0206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_232_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2921_ _0128_ _0136_ _0144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_204_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_231_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2852_ _0065_ _0066_ _0068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_79_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2783_ _1791_ _1793_ _1884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_15_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_157_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3404_ _0599_ _0603_ _0675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_171_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_236_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_119_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3171__A1 _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3335_ _0590_ _0595_ _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_59_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3424__I dsynth.freeRunCntr\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3266_ _0521_ _0522_ _0523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_239_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2217_ _1318_ _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3197_ _0431_ _0433_ _0442_ _0447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XTAP_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_227_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2148_ _1242_ _1158_ _1250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_93_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_198_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2079_ _1178_ _1179_ _1159_ _1167_ _1180_ _1181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_78_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2985__A1 _0142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_206_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3529__A3 _0760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2659__B _1633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_172_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_162_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3465__A2 _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2394__B _1494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2976__A1 _0055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_213_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2440__A3 _1540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_224_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_199_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3672__C net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2288__C _1389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3120_ _0348_ _0363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_151_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3051_ _0275_ _0286_ _0287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_5580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2002_ _0558_ _0958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_212_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_223_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2904_ _0121_ _0123_ _0125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_162_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3884_ _0014_ net48 net32 dsynth.csTable.address\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_137_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2835_ _1785_ _1878_ _0049_ _0050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_192_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2766_ _1864_ _1865_ _1867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_129_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2697_ _1781_ _1796_ _1797_ _1798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_144_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_28_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3318_ _0578_ _0579_ _0581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_86_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3249_ _0251_ _0487_ _0486_ _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_189_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3383__A1 _0647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3383__B2 _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_221_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_207_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2413__A3 _1473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2143__I _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_146_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2620_ _1717_ _1719_ _1720_ _1319_ _1259_ _1721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_86_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_220_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2551_ _1589_ _1651_ _1652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1982__I _0734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2482_ _1235_ _1078_ _1582_ _1583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_173_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3126__A1 _1399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_233_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3103_ _0342_ _0343_ _0344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_3_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3429__A2 _1549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_231_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3034_ _1736_ _0182_ _0183_ _0268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_64_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2101__A2 _1170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_236_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_197_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout37_I net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_224_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3867_ _0028_ net55 net40 dsynth.freeRunCntr\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_108_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3149__I _1700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_197_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2818_ _1725_ _1726_ _0033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_3798_ _1123_ _1075_ _1077_ _1079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_191_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2749_ _1664_ _1849_ _1850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_105_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2656__C _1193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2891__A3 _0110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_234_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2628__B1 _1629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_210_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output18_I net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_187_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_204_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2159__A2 _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_237_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3108__A1 _0303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_215_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2331__A2 _1432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_179_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1977__I _0679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1982_ _0734_ _0745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3721_ _0978_ _1004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_158_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3652_ _0928_ _0930_ _0912_ _0946_ _0947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_146_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3347__A1 _0587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2603_ _1703_ _1704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_200_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3583_ _0869_ _0870_ _0814_ _0872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_115_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2534_ _1609_ _1635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_192_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2570__A2 _1668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_244_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2465_ _1563_ _1565_ _1566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_9_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2396_ _1496_ _1497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_228_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2322__A2 _1403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2048__I _1149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3017_ _1898_ _0249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_240_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_205_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_74_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_245_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2001__B2 _0942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2250_ _1221_ _1351_ _1352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_239_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2181_ _1281_ _1282_ _0931_ _1283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_226_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_225_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_221_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1965_ _0547_ _0558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3704_ _0969_ _0987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_198_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3635_ dsynth.freeRunCntr\[7\] _1528_ _1544_ _1313_ _0928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_31_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3566_ _0827_ _0837_ _0839_ _0825_ _0852_ _0853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_143_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2517_ _1541_ _1542_ _1618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3497_ _0739_ _0776_ _0777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_157_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2448_ _1548_ _1549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2487__B _1587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_229_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2379_ _1286_ _1479_ _1480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_5_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_212_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_164_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_240_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2950__B _1298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_228_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2231__A1 _1245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3731__A1 dsynth.freeRunCntr\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_181_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2298__A1 _1344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_207_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3800__I _1075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3798__A1 _1123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_231_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_203_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_proj_example_220 io_out[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_116_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3420_ _1464_ _0682_ _0688_ _0692_ _0693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_7_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3351_ _1807_ _1832_ _1837_ _0616_ _0617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_124_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2302_ _1360_ _1404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3282_ _0529_ _0530_ _0541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_48_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input9_I io_in[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2233_ _1332_ _1295_ _1333_ _1334_ _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_230_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2289__A1 _1331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_227_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2164_ _1265_ _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_66_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2095_ dsynth.csTable.address\[1\] dsynth.csTable.address\[2\] _1197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_78_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2461__A1 _1194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_181_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2997_ _0224_ _0225_ _0227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1948_ _0360_ _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3618_ _0651_ _1728_ _1858_ _0655_ _0910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_239_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3549_ _0832_ _0834_ _0835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_66_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2236__I _1337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2452__A1 _1240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_240_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_226_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_205_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_125_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_209_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2920_ _0117_ _0119_ _0143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_245_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3640__B1 _0048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2851_ _0065_ _0066_ _0067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_223_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2782_ _1876_ _1881_ _1882_ _1883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2746__A2 _1845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3403_ _0589_ _0597_ _0674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_171_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3334_ _0589_ _0597_ _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3265_ _0262_ _0494_ _0522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2216_ _1317_ _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3196_ _0403_ _0424_ _0443_ _0445_ _0446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_54_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3474__A3 _0611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_226_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2147_ _1241_ _1248_ _1249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_81_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2078_ _0778_ _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_243_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_241_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_148_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2737__A2 _1309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_202_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_200_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_162_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_176_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_241_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_242_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3050_ _0281_ _0284_ _0285_ _0286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_5570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2001_ _0800_ _0404_ _0920_ _0942_ _0952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_222_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_224_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2416__A1 _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_223_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3873__CLK net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_204_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2903_ _0121_ _0123_ _0124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_182_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_220_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3883_ _0013_ net48 net32 dsynth.csTable.address\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_143_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2834_ _0048_ _1527_ _1579_ _0049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_121_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2765_ _1364_ _1479_ _1866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_129_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2696_ _1794_ _1795_ _1797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_145_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2352__B1 _1312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3317_ _0554_ _0560_ _0539_ _0533_ _0555_ _0579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_141_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3248_ _0501_ _0502_ _0504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_246_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_227_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2655__A1 _1245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3179_ _0406_ _0423_ _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_2218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_148_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2407__A1 _1128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_223_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_210_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_132_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_199_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3071__A1 _0293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2550_ _0096_ _1650_ _1651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_127_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2481_ _1180_ _1333_ _1582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3126__A2 _1675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2885__A1 _1174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3102_ _1734_ _0202_ _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_6090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3033_ _0266_ _1728_ _0267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_209_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2637__B2 _1737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2101__A3 _1199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3062__A1 _1714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3866_ _0027_ net55 net40 dsynth.freeRunCntr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_176_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2817_ _1506_ _1917_ _1918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_3797_ _1072_ _1073_ _1076_ _1077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_164_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_178_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2748_ _1838_ _1491_ _1616_ _1848_ _1849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_117_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2679_ _1774_ _1777_ _1780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_86_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3117__A2 _0329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2628__A1 _1714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2953__B _1291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2800__A1 _1865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_211_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2180__S _1176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2159__A3 _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_202_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2316__B1 _1416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3659__A3 net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2867__A1 _1137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2095__A2 dsynth.csTable.address\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1981_ _0723_ _0734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_18_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_226_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3720_ _1003_ _0027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_158_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3595__A2 _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3651_ _0910_ _0945_ _0932_ _0946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_179_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2602_ _1264_ _1501_ _1703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_220_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3582_ _0814_ _0869_ _0870_ _0871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_173_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2533_ _1633_ _1583_ _1634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2103__B _0679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2464_ _1564_ _1554_ _1562_ _1565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_29_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2395_ _1480_ _1495_ _1496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_56_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_231_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3016_ _0243_ _0246_ _0247_ _0248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_25_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_224_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_193_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3849_ _1486_ _1116_ _1476_ _1119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_138_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2546__B1 _1552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_234_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output30_I net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_210_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3813__A3 _1085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_216_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_223_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_204_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_221_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2180_ _0624_ _1164_ _1176_ _1282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3501__A2 _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_239_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_230_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_179_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_222_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1964_ _0536_ _0074_ _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_175_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3703_ _0986_ _0022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_159_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2240__A2 _1294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_198_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3634_ _0902_ _0904_ _0914_ _0926_ _0927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_162_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3565_ _0832_ _0834_ _0851_ _0852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_192_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3740__A2 _1022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2516_ _1616_ _1617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3496_ _0775_ _0750_ _0776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_216_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2447_ _1547_ _1548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2378_ _1473_ _1478_ _1479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_116_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_229_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3599__B _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_205_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_235_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2231__A2 _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_240_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_181_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2298__A2 _1198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_181_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_235_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3798__A2 _1075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xuser_proj_example_210 io_oeb[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_106_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_193_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3350_ _0083_ _0240_ _0612_ _0615_ _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_140_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2301_ _1351_ _1403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3281_ _0533_ _0538_ _0539_ _0540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_151_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2232_ _1189_ _1049_ _1334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_78_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2289__A2 _1202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2163_ _1264_ _1265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_96_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3238__A1 _0282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2094_ _0723_ _1196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_224_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_221_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2996_ _0224_ _0225_ _0226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_9_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1947_ _0151_ _0349_ _0360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_159_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2342__I _1443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3617_ _1465_ _0518_ _0908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_235_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3548_ _1132_ _0396_ _0834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_135_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3479_ _1807_ _1835_ _0758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_233_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_164_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2452__A2 _1552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2204__A2 _0701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_219_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_197_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_175_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_6420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_6486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_125_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2427__I _1527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_225_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3640__A1 _1233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_203_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3640__B2 _1230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2850_ _1883_ _1884_ _1874_ _0066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_176_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2781_ _1879_ _1880_ _1882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_172_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3402_ _0598_ _0604_ _0673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3333_ _0590_ _0595_ _0596_ _0597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3264_ _0518_ _0491_ _0520_ _0462_ _0521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_230_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_227_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2215_ _1040_ _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_152_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3195_ _0406_ _0423_ _0445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_66_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2146_ _1243_ _1244_ _1247_ _0470_ _1248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_215_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2077_ _0877_ _1179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_228_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_81_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2979_ _0200_ _0205_ _0207_ _0208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2198__A1 _1292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2198__B2 _1173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_137_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2247__I _0206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_232_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_231_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_209_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2113__A1 _1212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_236_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2000_ _0931_ _0942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_4870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2157__I _0569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3613__A1 _0684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2902_ _0122_ _1904_ _0123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_56_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3882_ _0012_ net47 net31 dsynth.csTable.address\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_177_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2833_ _1607_ _1608_ _0048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_160_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2764_ _1137_ _1502_ _1865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2695_ _1794_ _1795_ _1796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_144_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_236_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2352__A1 _1290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3316_ _0533_ _0538_ _0539_ _0578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_112_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2776__B _1609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3247_ _0466_ _0467_ _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_73_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3178_ _1430_ _0402_ _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_39_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2655__A2 _0514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3852__A1 _1473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2129_ dsynth.freeRunCntr\[12\] _1186_ _1229_ _1230_ _1231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_242_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_214_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2407__A2 _1507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_74_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2591__A1 _1687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_1737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3071__A2 _0308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2480_ _1566_ _1580_ _1581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_126_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_233_1727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3101_ _0297_ _0299_ _0341_ _0342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_6080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3032_ _1736_ _0266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_5390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2637__A2 _1692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_224_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3062__A2 _0098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3865_ _0026_ net55 net42 dsynth.freeRunCntr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_149_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2816_ _1514_ _1915_ _1916_ _1917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_149_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_176_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3796_ _0849_ _1071_ _1076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_176_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2747_ _1846_ _1847_ _1848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__3365__A3 _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_199_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_160_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2678_ _1774_ _1777_ _1778_ _1779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_132_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3125__I0 _1265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_246_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2628__A2 _1715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2953__C _1370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2564__A1 _1664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_201_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2316__A1 _1385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3863__CLK net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2316__B2 _1417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2867__A2 _1506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1980_ _0305_ dsynth.csTable.address\[0\] _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_1871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3650_ _0944_ _0911_ _0907_ _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_158_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2601_ _1701_ _1702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_228_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3581_ _0812_ _0813_ _0769_ _0870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_173_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2532_ _1533_ _1633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_154_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2463_ _0096_ _1564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_170_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2307__A1 _1250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2394_ _1228_ _1490_ _1494_ _1495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_233_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3015_ _0244_ _1493_ _1786_ _0247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_243_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_225_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout42_I net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_36_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3848_ _1117_ _0023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3779_ _1058_ _1054_ _1060_ _1061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2546__B2 _1153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3886__CLK net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_236_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_179_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_179_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_230_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2785__A1 _1883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2537__A1 _1580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_226_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1963_ dsynth.csTable.address\[5\] _0536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_193_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2776__A1 _1590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3702_ _0983_ _0985_ _0986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_204_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3633_ _0924_ _0925_ _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2114__B _0963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3564_ _0828_ _0829_ _0836_ _0851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_161_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2515_ _1513_ _1475_ _1472_ _1616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_89_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3495_ _0740_ _0746_ _0775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_130_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2446_ _1487_ _1546_ _1547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_237_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2377_ _1476_ _1477_ _1478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_64_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2700__A1 _1798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2075__I _1176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_244_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_240_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2231__A3 _0459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1990__A2 _0272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2298__A3 _1386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_216_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3798__A3 _1077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2758__A1 _1857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_proj_example_200 io_oeb[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
Xuser_proj_example_211 io_oeb[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_157_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_221_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2300_ _1401_ _1402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3280_ _0505_ _0506_ _0539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_193_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_234_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2231_ _1245_ _1237_ _0459_ _1177_ _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_97_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_239_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2162_ _1188_ _1263_ _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_187_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2093_ _0701_ _1195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3238__A2 _0461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2995_ _0126_ _0154_ _0225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2749__A1 _1664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1946_ dsynth.csTable.address\[3\] _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_124_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1972__A2 dsynth.csTable.address\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3616_ _1385_ _0045_ _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_162_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_200_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3547_ _1681_ _1515_ _0832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_85_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3478_ _1834_ _1832_ _0642_ _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_115_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_213_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2429_ _1475_ _1529_ _1530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_83_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_226_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_231_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_241_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2204__A3 _1200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_240_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_192_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_238_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_6498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3640__A2 _1683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_204_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_206_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2443__I _1543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3880__RN net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2780_ _1879_ _1880_ _1881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_156_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_200_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3401_ _0670_ _0449_ _0671_ _0672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_236_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3332_ _0593_ _0594_ _0596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3263_ _0518_ _0490_ _0519_ _0520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3459__A2 _0705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2214_ _0624_ _0657_ _1297_ _1316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_117_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3194_ _0401_ _0425_ _0430_ _0443_ _0444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_94_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_230_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2145_ _1245_ _1246_ _1247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_208_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2076_ _1175_ _1177_ _1178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_241_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2434__A3 _1274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_210_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_223_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3871__RN net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2978_ _0203_ _0204_ _0207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_241_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3395__A1 _0655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1929_ _0151_ dsynth.csTable.address\[4\] _0162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_147_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_235_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_89_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_183_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2263__I _1364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_231_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3862__RN net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2113__A2 _1214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_236_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3613__A2 _0295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2901_ _1380_ _1902_ _0122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_205_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3881_ _0010_ net47 net31 dsynth.csTable.address\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_162_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2832_ _0035_ _0046_ _0047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__2106__C _1207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2763_ _1087_ _1492_ _1863_ _1838_ _1864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_145_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1927__A2 _0129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_172_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2694_ _1729_ _1740_ _1795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_144_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2352__A2 _1287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3315_ _0554_ _0555_ _0574_ _0576_ _0577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_140_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_236_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3246_ _0488_ _0499_ _0500_ _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3301__A1 _0268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3177_ _0403_ _0424_ _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_215_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2128_ dsynth.freeRunCntr\[11\] _1230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_187_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_199_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2059_ _1160_ _1161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2258__I _0958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_181_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2031__A1 _1131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2031__B2 _1123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2334__A2 _1199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3531__A1 _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3100_ _1687_ _1714_ _0098_ _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_1_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2168__I _1223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3031_ _1858_ _0260_ _0263_ _0264_ _0265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XTAP_5380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2270__A1 _1301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3864_ _0022_ net55 net40 dsynth.freeRunCntr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_176_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2815_ _1337_ _1501_ _1916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_242_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3795_ _0967_ _1022_ _1075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_145_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2746_ _1842_ _1845_ _1574_ _1847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_173_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_172_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2677_ _1772_ _1773_ _1778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2078__I _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3125__I1 _1704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_210_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3229_ _0321_ _0358_ _0482_ _0483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_221_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2564__A2 _1631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2316__A2 _1399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_238_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_234_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2716__I _1668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2600_ _1124_ _1087_ _1701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_200_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2004__B2 _0963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3580_ _0772_ _0869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_127_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_155_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2555__A2 _1655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2531_ _1615_ _1631_ _1632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_192_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2462_ _1554_ _1562_ _1516_ _1563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_114_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3504__A1 _1634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3504__B2 _1596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2393_ _0118_ _1493_ _1494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_229_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3807__A2 _1085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_243_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3014_ _1786_ _0245_ _0246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_224_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_92_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout35_I net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3847_ _1486_ _1116_ _1117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_149_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2361__I _1417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3778_ dsynth.freeRunCntr\[11\] _1037_ _1051_ _1060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_88_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3743__A1 _0647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2546__A2 _1292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2729_ _1818_ _1829_ _1830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_133_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_161_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3274__A3 _0488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_243_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_215_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2482__A1 _1235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output16_I net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2234__A1 _1125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_180_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3431__B1 _1700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3431__C2 _1668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2785__A2 _1884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_195_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_178_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3316__B _0539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2220__B _0195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_206_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_221_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2225__A1 _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1962_ _0503_ _0514_ _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_239_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_222_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3701_ _0973_ _0976_ _0984_ _0985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_37_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3632_ _1463_ _0489_ _0925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_174_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3563_ _0843_ _0845_ _0846_ _0850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_143_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2514_ _1184_ _1500_ _1615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_3494_ _0773_ _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_115_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2445_ _1472_ _1545_ _1546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_233_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2376_ dsynth.freeRunCntr\[29\] _1477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2700__A2 _1799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_213_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2305__B _1358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2231__A4 _1177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_166_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2519__A2 _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_181_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_173_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_181_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_181_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2207__A1 _1291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_230_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2758__A2 _1858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_223_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_example_201 io_oeb[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
Xuser_proj_example_212 io_oeb[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_139_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3707__A1 _1419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2230_ _1214_ _1331_ _1332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2885__B _1334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2161_ _1236_ _1249_ _1254_ _1262_ _1263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_93_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2092_ _1193_ _1194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_207_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3876__CLK net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_226_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2994_ _0197_ _0222_ _0223_ _0224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_241_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1945_ _0217_ _0338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3615_ _0905_ _1848_ _0906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3546_ _0784_ _0785_ _0831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_89_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3477_ _0238_ _0752_ _0754_ _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_142_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2428_ _1513_ _1483_ _1529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_4508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2359_ _1340_ _1461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input15_I io_in[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2086__I _1010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2988__A2 _0211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3165__A2 _0211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3625__B1 _0702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_216_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_232_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3400_ _0666_ _0667_ _0517_ _0585_ _0446_ _0671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_236_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3331_ _0593_ _0594_ _0595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XTAP_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_119_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3262_ _0268_ _0490_ _0519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_45_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input7_I io_in[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2213_ _1195_ _1201_ _1315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_239_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3193_ _0431_ _0433_ _0442_ _0443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_132_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2144_ _0283_ _1246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_54_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2419__A1 _0789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2075_ _1176_ _1177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_53_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2977_ _0203_ _0204_ _0205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_210_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3395__A2 _0654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1928_ dsynth.csTable.address\[6\] _0151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_147_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2355__B1 _1139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3529_ _0757_ _0759_ _0760_ _0813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_1_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2658__A1 _1573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_211_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2897__A1 _1704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2900_ _0102_ _0120_ _0121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_204_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3880_ _0009_ net47 net31 dsynth.csTable.address\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__2821__A1 _1615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_242_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2831_ _1548_ _0033_ _0045_ _1532_ _1737_ _0046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_143_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_203_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2762_ _1484_ _1488_ _1863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_203_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2693_ _1784_ _1788_ _1789_ _1791_ _1793_ _1794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_184_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3314_ _0554_ _0555_ _0575_ _0576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_140_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3245_ _0496_ _0498_ _0500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3301__A2 _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_230_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3176_ _0406_ _0423_ _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_55_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2127_ _1228_ _1229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_82_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2058_ _0569_ _0931_ _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_179_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2812__A1 _1236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_223_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2879__A1 _1574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_18_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3056__A1 _0284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_221_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_207_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_199_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2223__B _1324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2031__A2 _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2334__A3 _1368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3030_ _1580_ _1528_ _0264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_5370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2893__B _0112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_231_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3834__A3 _1574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_225_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3863_ _0011_ net54 net41 dsynth.freeRunCntr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__2270__A2 _1258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2814_ _1636_ _1914_ _1915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_192_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3794_ _1074_ _0005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2745_ _1569_ _1842_ _1845_ _1846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_191_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2676_ _1775_ _1776_ _1777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_191_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_173_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_207_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_236_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3228_ _0479_ _0480_ _0482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_189_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3286__A1 _1429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_228_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3159_ _0325_ _0329_ _0405_ _0391_ _0362_ _0406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XTAP_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3038__A1 _0186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_203_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2094__I _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_204_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_183_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2218__B _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2530_ _1617_ _1618_ _1629_ _1630_ _1631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_170_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2888__B _1236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2461_ _1194_ _1558_ _1559_ _1561_ _1562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_244_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3504__A2 _0623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2392_ _1492_ _1493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_174_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_228_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3013_ _0244_ _1493_ _0245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_168_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2243__A2 _1344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3846_ _1114_ _1116_ _0021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_193_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3777_ _1036_ _1051_ dsynth.freeRunCntr\[11\] _1058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_14_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2728_ _1820_ _1828_ _1829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_88_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2798__B _1898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_175_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2659_ _1753_ _1758_ _1633_ _1760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_154_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_210_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_55_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_223_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3431__A1 _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3431__B2 _0991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3670__A1 net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2225__A2 _0283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1961_ _0338_ _0514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3700_ _1445_ _0975_ _0984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_175_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3631_ _0923_ _0924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_200_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3562_ dsynth.freeRunCntr\[14\] _0849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_31_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2513_ _1568_ _1612_ _1613_ _1614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_192_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3493_ _0747_ _0764_ _0766_ _0772_ _0773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_100_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2444_ dsynth.freeRunCntr\[29\] _1485_ _1545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2375_ _1475_ _1476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_229_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2161__A1 _1236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_245_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_216_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3661__A1 _0954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_227_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_212_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1975__A1 _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3829_ _0536_ _1101_ _1104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3716__A2 _0989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2152__A1 _1250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2455__A2 _1555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_231_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_example_202 io_oeb[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_8_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_example_213 io_oeb[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_11_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_151_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_239_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_155_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2160_ _1255_ _1260_ _1261_ _1262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_227_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3062__B _1687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_241_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2091_ _1191_ _1192_ _1193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_130_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_221_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_210_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2993_ _0220_ _0221_ _0223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_206_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2192__I _1197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_222_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1944_ _0316_ _0327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_128_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3614_ dsynth.freeRunCntr\[4\] _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_116_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3545_ _0828_ _0829_ _0830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3476_ _0083_ _0753_ _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_131_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2427_ _1527_ _1528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_233_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2358_ _1459_ _1312_ _1431_ _1383_ _1460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_69_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2289_ _1331_ _1202_ _1349_ _1391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_85_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_240_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_205_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3165__A3 _0411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_6489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_125_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2428__A2 _1483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3625__A1 dsynth.freeRunCntr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3625__B2 _1118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_223_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2600__A2 _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2364__A1 _1465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_236_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3330_ _0196_ _0222_ _0594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_152_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3261_ _0185_ _0518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2212_ _1313_ _1314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_230_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3192_ _0436_ _0441_ _0442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_6_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2143_ _0624_ _1245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_43_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_226_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2074_ _0723_ _1176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__3616__A1 _1385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_228_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2976_ _0055_ _0132_ _0204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_50_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2052__B1 _1150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1927_ _0063_ _0129_ _0140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_175_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2355__A1 _0140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2355__B2 _1456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3528_ _0809_ _0810_ _0753_ _0083_ _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_118_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3459_ _0733_ _0705_ _0735_ _0736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_103_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2097__I _1198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3607__A1 _1464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_240_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2594__A1 _1682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2346__A1 _1417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3866__CLK net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_218_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3074__A2 _1504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_232_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2830_ _1846_ _1847_ _0045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_231_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2761_ _1860_ _1861_ _1862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2692_ _1788_ _1792_ _1793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_177_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3313_ _0561_ _0564_ _0570_ _0571_ _0567_ _0575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_59_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3244_ _0496_ _0498_ _0499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_100_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3175_ _0407_ _0422_ _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_26_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2126_ _1227_ _1228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_227_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout58_I net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_148_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2057_ _1158_ _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_78_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_210_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_206_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2959_ _1379_ _1492_ _0186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_194_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3889__CLK net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2500__A1 _0459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_198_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_241_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_224_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3386__I _1382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_177_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2319__A1 _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_163_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_6094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_204_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3862_ _0000_ net53 net41 dsynth.freeRunCntr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_31_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2813_ _1908_ _1910_ _1911_ _1913_ _1914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_3793_ _1072_ _1073_ _1074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_176_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_176_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2744_ _1396_ _1843_ _1844_ _1845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_118_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_199_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2675_ _1087_ _1498_ _1776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_201_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_173_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3227_ _0259_ _0319_ _0480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_246_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3286__A2 _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3158_ _0362_ _0391_ _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_2008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2109_ _0657_ _1210_ _0844_ _1211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_43_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3089_ _0326_ _0328_ _0329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3210__A2 _1848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_232_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2285__I _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3110__S _0351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2960__A1 _1514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2460_ _1318_ _1438_ _1560_ _1217_ _1561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_142_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2391_ _1491_ _1492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_174_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2712__A1 _1665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_218_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3012_ _0129_ _1442_ _0244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_5190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_209_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3020__S _0252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3845_ _1115_ _1116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_149_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3776_ _0697_ _1056_ _1057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_164_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2727_ _1821_ _1827_ _1828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_175_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2951__A1 _1394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2951__B2 _1648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2658_ _1573_ _1753_ _1758_ _1759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_47_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2589_ _0920_ _1644_ _1646_ _1688_ _1689_ _1690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_160_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_236_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_184_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3431__A2 _0256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2054__B _0690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3664__I net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2501__C _1217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2170__A2 _1176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_218_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1960_ _0492_ _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_226_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_230_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3630_ _0698_ _0707_ _0915_ _0922_ _0923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_159_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3186__A1 _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_239_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3561_ _0841_ _0847_ _1136_ _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_127_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2512_ _1593_ _1611_ _1613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_3492_ _0618_ _0642_ _0763_ _0772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_154_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2443_ _1543_ _1544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2374_ _1474_ _1475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2139__B _1069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2464__A3 _1562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout40_I net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_240_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2621__B1 _1282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_220_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3828_ _1102_ _0015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3759_ _1290_ _1039_ _1041_ _1042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_118_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_165_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_181_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_229_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output21_I net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2563__I _1615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3892__RN net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3404__A2 _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_212_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xuser_proj_example_203 io_oeb[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_106_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_proj_example_214 io_oeb[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_171_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2090_ _1049_ _1192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_47_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_222_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2473__I _1573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3883__RN net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2992_ _0220_ _0221_ _0222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1943_ _0305_ dsynth.csTable.address\[1\] _0316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_175_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3613_ _0684_ _0295_ _0903_ _0904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2422__B _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2906__A1 _0097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3544_ _0782_ _0787_ _0829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_192_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_235_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3475_ _1836_ _0643_ _0753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_157_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2509__I1 _1584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2426_ _1516_ _1526_ _1527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_213_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_229_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2357_ _1314_ _1459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2288_ _1291_ _1386_ _1388_ _1152_ _1389_ _1390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_84_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_212_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2383__I _1483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3874__RN net58 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2125__A2 _1226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_197_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_87_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_235_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3625__A2 _1586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2507__B _1573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3865__RN net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_240_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_193_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2364__A2 _1444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3260_ _0485_ _0515_ _0516_ _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2211_ dsynth.freeRunCntr\[8\] _1313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3191_ _0439_ _0440_ _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_227_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2142_ _0503_ _1175_ _1244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_66_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2073_ _1164_ _1175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_78_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3616__A2 _0045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_223_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_206_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2975_ _1618_ _0201_ _0202_ _1734_ _0203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_37_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2052__A1 _1143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1926_ _0118_ _0129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2052__B2 _1152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2152__B _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3527_ _0231_ _0235_ _0611_ _0810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_104_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3458_ _0700_ _0704_ _0735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_5008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2409_ _1498_ _1509_ _1508_ _1510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_97_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3389_ _1459_ _0644_ _0652_ _0656_ _0658_ _1461_ _0659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
XTAP_4307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2658__A3 _1758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_81_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2291__A1 _1374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2346__A2 _1416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3059__B1 _0295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_223_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2760_ _1775_ _1776_ _1861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_203_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_185_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2585__A2 _1655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2691_ _1588_ _1783_ _1792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_117_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2337__A2 _1438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3534__A1 _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_236_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3312_ _0560_ _0573_ _0574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_112_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3243_ _0054_ _0497_ _0498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_136_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_230_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3174_ _0409_ _0421_ _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_67_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2125_ _1188_ _1226_ _1227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_81_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2056_ _1144_ _1157_ _1158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_228_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2273__A1 _1374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2958_ _0182_ _0183_ _0185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3773__A1 _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2889_ _1331_ _1202_ _1301_ _1389_ _0109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_124_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3289__B1 _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_181_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2500__A2 _1331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_220_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2319__A2 _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_224_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2682__S _1733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2255__A1 _1175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3861_ net6 _1919_ tgate.clkp vdd vss gf180mcu_fd_sc_mcu7t5v0__latq_1
XFILLER_220_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2812_ _1236_ _1912_ _1913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3792_ _1066_ _1068_ _1065_ _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_121_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2743_ _1238_ _1604_ _1322_ _1259_ _1844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_157_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2674_ _1338_ _1666_ _1670_ _1364_ _1675_ _1286_ _1775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_4
XFILLER_160_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3226_ _0476_ _0477_ _0478_ _0479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_210_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2494__A1 _1236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3157_ _1430_ _0402_ _0403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_227_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2108_ _1209_ _1210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_243_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3088_ _1414_ _1675_ _1507_ _0328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_184_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_82_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2039_ _1140_ _1141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2246__A1 _1345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2246__B2 _1347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2391__I _1491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_210_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_218_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2566__I _1666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_198_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2788__A2 _1888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2960__A2 _0185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2390_ _1475_ _1472_ _1482_ _1491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_96_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3011_ _0186_ _0243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_5180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3879__CLK net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_225_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2228__A1 _0833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_225_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3844_ _1477_ dsynth.freeRunCntr\[28\] _1112_ _1115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_162_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3775_ _1050_ _1036_ _0995_ _1056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_164_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_199_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2726_ _1822_ _1826_ _1827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_145_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2951__A2 _1277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2657_ _1259_ _1754_ _1755_ _1757_ _1758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_86_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2588_ _1190_ _1317_ _1401_ _0382_ _1689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_160_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3209_ _1915_ _0461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_219_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2458__A1 _1156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_207_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_199_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2630__A1 _1577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_187_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3560_ _0843_ _0845_ _0846_ _0847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2511_ _1593_ _1611_ _1612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_183_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3491_ _0755_ _0761_ _0770_ _0771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2442_ _1541_ _1542_ _1543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_142_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2146__B1 _1247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2373_ dsynth.freeRunCntr\[31\] _1474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2449__A1 _1176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3646__B1 _1681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3661__A3 net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout33_I net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2621__A1 _1243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2621__B2 _1538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_222_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3827_ _0536_ _1101_ _1102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_197_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_229_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_229_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3758_ _1031_ _1034_ _1029_ _1041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_10_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2709_ _1511_ _1808_ _1809_ _1810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3689_ dsynth.freeRunCntr\[0\] _0972_ _0973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_173_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2688__A1 _1782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_181_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2612__A1 _1633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_230_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_183_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xuser_proj_example_204 io_oeb[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_7_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_example_215 io_oeb[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_128_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_221_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_234_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_206_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2991_ _0148_ _0149_ _0221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_222_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_226_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1942_ dsynth.csTable.address\[6\] _0305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_159_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3159__A2 _0329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3612_ _0684_ _0295_ _0518_ _1445_ _0903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_102_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3543_ _0783_ _0786_ _0828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_200_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3474_ _0230_ _0235_ _0611_ _0752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_171_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2425_ _1520_ _1525_ _0958_ _1526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_237_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2356_ _1290_ _1287_ _1289_ _1139_ _1458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_85_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_229_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2287_ _1304_ _1389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_226_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2664__I _1715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2842__B2 _1635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_225_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_192_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_238_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_192_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_6447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2530__B1 _1629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_125_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_229_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_216_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_229_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_231_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2523__B _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_196_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3010__A1 _1311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2210_ _1311_ _1312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_171_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3190_ _0215_ _0216_ _0440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_67_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2141_ _1242_ _1243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2072_ _1170_ _1173_ _1174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3077__A1 _0291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_208_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_207_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_223_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2974_ _1786_ _1543_ _0201_ _0202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_194_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1925_ _0107_ _0118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2052__A2 _1148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_206_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3526_ _0236_ _0237_ _0809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_235_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3457_ _0700_ _0704_ _0733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_5009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2408_ _1503_ _1506_ _1508_ _1509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3388_ _1836_ _0616_ _0658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_130_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2339_ _1387_ _1357_ _1439_ _1440_ _1441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_242_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input13_I io_in[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2815__A1 _1337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_246_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2291__A2 _1242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2579__B1 _1515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3791__A2 _1071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_155_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_6211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_6233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3059__A1 _0282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2518__B _1166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2806__A1 _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_217_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_182_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_203_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_199_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2690_ _1790_ _1766_ _1791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_12_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2742__B1 _1556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3311_ _0570_ _0571_ _0572_ _0573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2479__I _1579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3242_ _0336_ _0260_ _0463_ _0497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_input5_I io_in[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_112_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3173_ _0412_ _0420_ _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_66_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2124_ _1194_ _1203_ _1208_ _1216_ _1225_ _1226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_215_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2055_ dsynth.csTable.address\[2\] _1157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_35_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2273__A2 _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2957_ _0178_ _0181_ _0112_ _0183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2025__A2 _1126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2888_ _1406_ _1387_ _1236_ _0108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_135_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2389__I _1489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3509_ _0732_ _0736_ _0791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_28_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3289__A1 _0489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2500__A3 _1270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2264__A2 _1358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_207_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2319__A3 _1323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2520__C _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2255__A2 _1246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3452__A1 _1702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3860_ tmux.clkpba net5 tmux.clkpbb vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2811_ _1178_ _1346_ _1251_ _1238_ _1319_ _1912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__3204__A1 _0090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3791_ _0849_ _1071_ _1072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_34_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_160_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_242_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2742_ _1170_ _1316_ _1523_ _1556_ _0668_ _1843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_117_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2673_ _1772_ _1773_ _1774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_117_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_236_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2191__A1 _1167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2002__I _0558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3225_ _0474_ _0475_ _0478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_67_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3156_ _0396_ _0402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_94_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3691__A1 net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_228_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2107_ _0250_ _1157_ _1209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_3_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3087_ _1443_ _1666_ _0326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2038_ _0613_ _1140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2246__A2 _1346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3746__A2 _0970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2954__B1 _1250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_213_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_172_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3678__I net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2582__I _1566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_237_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3010_ _1311_ _0241_ _0242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_5170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_224_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2228__A2 _1327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1987__A1 _0668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3843_ dsynth.freeRunCntr\[28\] _1112_ _1477_ _1114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_203_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3774_ _1055_ _0002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2725_ _1823_ _1825_ _1826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_173_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3029__S _0260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2656_ _1538_ _1756_ _1375_ _1193_ _1757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_12_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2587_ _0448_ _0833_ _1688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_82_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_216_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_232_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3208_ _0455_ _0458_ _0460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_86_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_227_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_216_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3139_ _0090_ _0312_ _0352_ _0175_ _0384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_103_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_243_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2616__B _1206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2458__A2 _1173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3655__A1 _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_222_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3201__I _0351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1969__A1 dsynth.csTable.address\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_239_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2630__A2 _1730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2394__A1 _1228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2510_ _1597_ _1610_ _1611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_154_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_196_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3490_ _0766_ _0769_ _0770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_185_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2441_ _1536_ _1540_ _1533_ _1542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_174_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2146__A1 _1243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2146__B2 _0470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2372_ _1472_ _1473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_233_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_229_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2449__A2 _1294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3646__A1 _1123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_209_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3646__B2 _1131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_225_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2436__B _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_209_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_221_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_240_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2621__A2 _1150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3826_ _0349_ _1093_ dsynth.csTable.address\[4\] _1094_ _1101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_21_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2171__B _1272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3757_ _1037_ _1038_ _1039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2708_ _1662_ _1698_ _1809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_145_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3688_ _0967_ _0970_ _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_106_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2639_ _1738_ _1739_ _1740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_133_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_173_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2397__I _1494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_215_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_204_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_example_205 io_oeb[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_184_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xuser_proj_example_216 io_oeb[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_11_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3869__CLK net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_155_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_189_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2256__B _1167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2990_ _0215_ _0216_ _0219_ _0220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1941_ _0239_ _0283_ _0294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_241_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3611_ _1463_ _0489_ _0902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_174_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3542_ _0788_ _0790_ _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_183_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3473_ _0739_ _0750_ _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2424_ _1318_ _1521_ _1522_ _1524_ _1525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_142_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2355_ _0140_ _1134_ _1139_ _1456_ _1457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_170_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2286_ _1218_ _1387_ _1388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3619__A1 _1382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2842__A2 _0054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_246_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3809_ dsynth.freeRunCntr\[17\] _1085_ _1088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_6426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3322__A3 _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2530__B2 _1630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3686__I net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3849__A1 _1486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_234_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2140_ _0899_ _1242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2071_ _1171_ _1172_ _1173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_93_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_234_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2973_ _1587_ _1846_ _1847_ _0201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_72_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1924_ _0085_ _0096_ _0107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_147_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2433__C _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3525_ _0805_ _0808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_137_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3456_ _0728_ _0731_ _0732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_83_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2407_ _1128_ _1507_ _1508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_3387_ _0651_ _0650_ _0654_ _0655_ _0656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_85_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2338_ _1224_ _1205_ _1258_ _1387_ _1434_ _1440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_6_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2269_ _1366_ _1369_ _1370_ _1371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_226_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_148_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2624__B _1569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2579__A1 _1185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2579__B2 _1678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_224_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2751__A1 _1590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_6212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_6289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3059__A2 _1528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_216_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2806__A2 _1619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_231_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_164_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_200_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2742__A1 _1170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2742__B2 _0668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3310_ _0557_ _0559_ _0572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_153_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3241_ _0489_ _0491_ _0495_ _0496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_141_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3172_ _0414_ _0419_ _0420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_41_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2123_ _1218_ _1222_ _1224_ _1225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_55_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2054_ _0514_ _1155_ _0690_ _1156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_235_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_207_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_194_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2956_ _0112_ _0178_ _0181_ _0182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_124_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_206_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2887_ _1170_ _1523_ _0105_ _1215_ _1421_ _0106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__2981__A1 _0208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_219_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_219_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3508_ _0728_ _0731_ _0790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_131_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3439_ _0710_ _0713_ _0714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_106_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3289__A2 _0268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_217_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_57_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2319__A4 _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput30 net30 io_out[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_107_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_225_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3452__A2 _0159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_205_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2810_ _1207_ _1354_ _1244_ _1911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3790_ _1050_ _1037_ _1011_ _1071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_125_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2741_ _1839_ _1840_ _1841_ _0580_ _1842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_201_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2672_ _1311_ _1667_ _1670_ _1339_ _1676_ _1265_ _1773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_4
XFILLER_172_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2191__A2 _1246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_236_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3224_ _1444_ _0256_ _0455_ _0458_ _0477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
.ends

