magic
tech gf180mcuC
magscale 1 5
timestamp 1670260778
<< metal1 >>
rect 672 6285 7360 6302
rect 672 6259 2259 6285
rect 2285 6259 2311 6285
rect 2337 6259 2363 6285
rect 2389 6259 3911 6285
rect 3937 6259 3963 6285
rect 3989 6259 4015 6285
rect 4041 6259 5563 6285
rect 5589 6259 5615 6285
rect 5641 6259 5667 6285
rect 5693 6259 7215 6285
rect 7241 6259 7267 6285
rect 7293 6259 7319 6285
rect 7345 6259 7360 6285
rect 672 6242 7360 6259
rect 1185 6119 1191 6145
rect 1217 6119 1223 6145
rect 1745 6063 1751 6089
rect 1777 6063 1783 6089
rect 3201 6063 3207 6089
rect 3233 6063 3239 6089
rect 5049 6063 5055 6089
rect 5081 6063 5087 6089
rect 3425 6007 3431 6033
rect 3457 6007 3463 6033
rect 5385 6007 5391 6033
rect 5417 6007 5423 6033
rect 672 5893 7280 5910
rect 672 5867 1433 5893
rect 1459 5867 1485 5893
rect 1511 5867 1537 5893
rect 1563 5867 3085 5893
rect 3111 5867 3137 5893
rect 3163 5867 3189 5893
rect 3215 5867 4737 5893
rect 4763 5867 4789 5893
rect 4815 5867 4841 5893
rect 4867 5867 6389 5893
rect 6415 5867 6441 5893
rect 6467 5867 6493 5893
rect 6519 5867 7280 5893
rect 672 5850 7280 5867
rect 961 5727 967 5753
rect 993 5727 999 5753
rect 6001 5727 6007 5753
rect 6033 5727 6039 5753
rect 1521 5671 1527 5697
rect 1553 5671 1559 5697
rect 5441 5671 5447 5697
rect 5473 5671 5479 5697
rect 672 5501 7360 5518
rect 672 5475 2259 5501
rect 2285 5475 2311 5501
rect 2337 5475 2363 5501
rect 2389 5475 3911 5501
rect 3937 5475 3963 5501
rect 3989 5475 4015 5501
rect 4041 5475 5563 5501
rect 5589 5475 5615 5501
rect 5641 5475 5667 5501
rect 5693 5475 7215 5501
rect 7241 5475 7267 5501
rect 7293 5475 7319 5501
rect 7345 5475 7360 5501
rect 672 5458 7360 5475
rect 672 5109 7280 5126
rect 672 5083 1433 5109
rect 1459 5083 1485 5109
rect 1511 5083 1537 5109
rect 1563 5083 3085 5109
rect 3111 5083 3137 5109
rect 3163 5083 3189 5109
rect 3215 5083 4737 5109
rect 4763 5083 4789 5109
rect 4815 5083 4841 5109
rect 4867 5083 6389 5109
rect 6415 5083 6441 5109
rect 6467 5083 6493 5109
rect 6519 5083 7280 5109
rect 672 5066 7280 5083
rect 672 4717 7360 4734
rect 672 4691 2259 4717
rect 2285 4691 2311 4717
rect 2337 4691 2363 4717
rect 2389 4691 3911 4717
rect 3937 4691 3963 4717
rect 3989 4691 4015 4717
rect 4041 4691 5563 4717
rect 5589 4691 5615 4717
rect 5641 4691 5667 4717
rect 5693 4691 7215 4717
rect 7241 4691 7267 4717
rect 7293 4691 7319 4717
rect 7345 4691 7360 4717
rect 672 4674 7360 4691
rect 672 4325 7280 4342
rect 672 4299 1433 4325
rect 1459 4299 1485 4325
rect 1511 4299 1537 4325
rect 1563 4299 3085 4325
rect 3111 4299 3137 4325
rect 3163 4299 3189 4325
rect 3215 4299 4737 4325
rect 4763 4299 4789 4325
rect 4815 4299 4841 4325
rect 4867 4299 6389 4325
rect 6415 4299 6441 4325
rect 6467 4299 6493 4325
rect 6519 4299 7280 4325
rect 672 4282 7280 4299
rect 672 3933 7360 3950
rect 672 3907 2259 3933
rect 2285 3907 2311 3933
rect 2337 3907 2363 3933
rect 2389 3907 3911 3933
rect 3937 3907 3963 3933
rect 3989 3907 4015 3933
rect 4041 3907 5563 3933
rect 5589 3907 5615 3933
rect 5641 3907 5667 3933
rect 5693 3907 7215 3933
rect 7241 3907 7267 3933
rect 7293 3907 7319 3933
rect 7345 3907 7360 3933
rect 672 3890 7360 3907
rect 2367 3849 2393 3855
rect 2367 3817 2393 3823
rect 3487 3849 3513 3855
rect 3487 3817 3513 3823
rect 3991 3849 4017 3855
rect 3991 3817 4017 3823
rect 2367 3737 2393 3743
rect 2367 3705 2393 3711
rect 2535 3737 2561 3743
rect 2535 3705 2561 3711
rect 3375 3737 3401 3743
rect 3375 3705 3401 3711
rect 3487 3737 3513 3743
rect 3487 3705 3513 3711
rect 3599 3737 3625 3743
rect 4159 3737 4185 3743
rect 3929 3711 3935 3737
rect 3961 3711 3967 3737
rect 3599 3705 3625 3711
rect 4159 3705 4185 3711
rect 2423 3625 2449 3631
rect 2423 3593 2449 3599
rect 4047 3625 4073 3631
rect 4047 3593 4073 3599
rect 672 3541 7280 3558
rect 672 3515 1433 3541
rect 1459 3515 1485 3541
rect 1511 3515 1537 3541
rect 1563 3515 3085 3541
rect 3111 3515 3137 3541
rect 3163 3515 3189 3541
rect 3215 3515 4737 3541
rect 4763 3515 4789 3541
rect 4815 3515 4841 3541
rect 4867 3515 6389 3541
rect 6415 3515 6441 3541
rect 6467 3515 6493 3541
rect 6519 3515 7280 3541
rect 672 3498 7280 3515
rect 2199 3457 2225 3463
rect 2199 3425 2225 3431
rect 2871 3345 2897 3351
rect 2871 3313 2897 3319
rect 3151 3345 3177 3351
rect 3151 3313 3177 3319
rect 3487 3345 3513 3351
rect 3487 3313 3513 3319
rect 2479 3289 2505 3295
rect 2479 3257 2505 3263
rect 2255 3233 2281 3239
rect 2255 3201 2281 3207
rect 2367 3233 2393 3239
rect 2367 3201 2393 3207
rect 3095 3233 3121 3239
rect 3095 3201 3121 3207
rect 3207 3233 3233 3239
rect 3207 3201 3233 3207
rect 672 3149 7360 3166
rect 672 3123 2259 3149
rect 2285 3123 2311 3149
rect 2337 3123 2363 3149
rect 2389 3123 3911 3149
rect 3937 3123 3963 3149
rect 3989 3123 4015 3149
rect 4041 3123 5563 3149
rect 5589 3123 5615 3149
rect 5641 3123 5667 3149
rect 5693 3123 7215 3149
rect 7241 3123 7267 3149
rect 7293 3123 7319 3149
rect 7345 3123 7360 3149
rect 672 3106 7360 3123
rect 3823 3065 3849 3071
rect 3823 3033 3849 3039
rect 3879 3009 3905 3015
rect 3879 2977 3905 2983
rect 4103 3009 4129 3015
rect 4103 2977 4129 2983
rect 2591 2953 2617 2959
rect 2591 2921 2617 2927
rect 2815 2953 2841 2959
rect 2815 2921 2841 2927
rect 672 2757 7280 2774
rect 672 2731 1433 2757
rect 1459 2731 1485 2757
rect 1511 2731 1537 2757
rect 1563 2731 3085 2757
rect 3111 2731 3137 2757
rect 3163 2731 3189 2757
rect 3215 2731 4737 2757
rect 4763 2731 4789 2757
rect 4815 2731 4841 2757
rect 4867 2731 6389 2757
rect 6415 2731 6441 2757
rect 6467 2731 6493 2757
rect 6519 2731 7280 2757
rect 672 2714 7280 2731
rect 3263 2617 3289 2623
rect 3263 2585 3289 2591
rect 2087 2561 2113 2567
rect 2249 2535 2255 2561
rect 2281 2535 2287 2561
rect 2087 2529 2113 2535
rect 2143 2505 2169 2511
rect 2143 2473 2169 2479
rect 2367 2505 2393 2511
rect 2367 2473 2393 2479
rect 3039 2505 3065 2511
rect 3039 2473 3065 2479
rect 3151 2505 3177 2511
rect 3151 2473 3177 2479
rect 3319 2505 3345 2511
rect 3319 2473 3345 2479
rect 911 2449 937 2455
rect 911 2417 937 2423
rect 672 2365 7360 2382
rect 672 2339 2259 2365
rect 2285 2339 2311 2365
rect 2337 2339 2363 2365
rect 2389 2339 3911 2365
rect 3937 2339 3963 2365
rect 3989 2339 4015 2365
rect 4041 2339 5563 2365
rect 5589 2339 5615 2365
rect 5641 2339 5667 2365
rect 5693 2339 7215 2365
rect 7241 2339 7267 2365
rect 7293 2339 7319 2365
rect 7345 2339 7360 2365
rect 672 2322 7360 2339
rect 2199 2281 2225 2287
rect 2199 2249 2225 2255
rect 2535 2281 2561 2287
rect 2535 2249 2561 2255
rect 2703 2281 2729 2287
rect 2703 2249 2729 2255
rect 3263 2281 3289 2287
rect 3263 2249 3289 2255
rect 3767 2281 3793 2287
rect 3767 2249 3793 2255
rect 2647 2225 2673 2231
rect 2647 2193 2673 2199
rect 3207 2225 3233 2231
rect 3207 2193 3233 2199
rect 2759 2169 2785 2175
rect 1521 2143 1527 2169
rect 1553 2143 1559 2169
rect 2081 2143 2087 2169
rect 2113 2143 2119 2169
rect 2759 2137 2785 2143
rect 2983 2169 3009 2175
rect 2983 2137 3009 2143
rect 3319 2169 3345 2175
rect 3319 2137 3345 2143
rect 3599 2169 3625 2175
rect 3599 2137 3625 2143
rect 3767 2169 3793 2175
rect 3767 2137 3793 2143
rect 3935 2169 3961 2175
rect 3935 2137 3961 2143
rect 5727 2113 5753 2119
rect 961 2087 967 2113
rect 993 2087 999 2113
rect 5727 2081 5753 2087
rect 672 1973 7280 1990
rect 672 1947 1433 1973
rect 1459 1947 1485 1973
rect 1511 1947 1537 1973
rect 1563 1947 3085 1973
rect 3111 1947 3137 1973
rect 3163 1947 3189 1973
rect 3215 1947 4737 1973
rect 4763 1947 4789 1973
rect 4815 1947 4841 1973
rect 4867 1947 6389 1973
rect 6415 1947 6441 1973
rect 6467 1947 6493 1973
rect 6519 1947 7280 1973
rect 672 1930 7280 1947
rect 1689 1807 1695 1833
rect 1721 1807 1727 1833
rect 3593 1807 3599 1833
rect 3625 1807 3631 1833
rect 2361 1751 2367 1777
rect 2393 1751 2399 1777
rect 5553 1751 5559 1777
rect 5585 1751 5591 1777
rect 2087 1721 2113 1727
rect 1017 1695 1023 1721
rect 1049 1695 1055 1721
rect 2087 1689 2113 1695
rect 2479 1721 2505 1727
rect 3879 1721 3905 1727
rect 2921 1695 2927 1721
rect 2953 1695 2959 1721
rect 2479 1689 2505 1695
rect 3879 1689 3905 1695
rect 4103 1721 4129 1727
rect 4103 1689 4129 1695
rect 4271 1721 4297 1727
rect 4271 1689 4297 1695
rect 6063 1721 6089 1727
rect 6063 1689 6089 1695
rect 6343 1721 6369 1727
rect 6343 1689 6369 1695
rect 5447 1665 5473 1671
rect 5447 1633 5473 1639
rect 5895 1665 5921 1671
rect 5895 1633 5921 1639
rect 672 1581 7360 1598
rect 672 1555 2259 1581
rect 2285 1555 2311 1581
rect 2337 1555 2363 1581
rect 2389 1555 3911 1581
rect 3937 1555 3963 1581
rect 3989 1555 4015 1581
rect 4041 1555 5563 1581
rect 5589 1555 5615 1581
rect 5641 1555 5667 1581
rect 5693 1555 7215 1581
rect 7241 1555 7267 1581
rect 7293 1555 7319 1581
rect 7345 1555 7360 1581
rect 672 1538 7360 1555
<< via1 >>
rect 2259 6259 2285 6285
rect 2311 6259 2337 6285
rect 2363 6259 2389 6285
rect 3911 6259 3937 6285
rect 3963 6259 3989 6285
rect 4015 6259 4041 6285
rect 5563 6259 5589 6285
rect 5615 6259 5641 6285
rect 5667 6259 5693 6285
rect 7215 6259 7241 6285
rect 7267 6259 7293 6285
rect 7319 6259 7345 6285
rect 1191 6119 1217 6145
rect 1751 6063 1777 6089
rect 3207 6063 3233 6089
rect 5055 6063 5081 6089
rect 3431 6007 3457 6033
rect 5391 6007 5417 6033
rect 1433 5867 1459 5893
rect 1485 5867 1511 5893
rect 1537 5867 1563 5893
rect 3085 5867 3111 5893
rect 3137 5867 3163 5893
rect 3189 5867 3215 5893
rect 4737 5867 4763 5893
rect 4789 5867 4815 5893
rect 4841 5867 4867 5893
rect 6389 5867 6415 5893
rect 6441 5867 6467 5893
rect 6493 5867 6519 5893
rect 967 5727 993 5753
rect 6007 5727 6033 5753
rect 1527 5671 1553 5697
rect 5447 5671 5473 5697
rect 2259 5475 2285 5501
rect 2311 5475 2337 5501
rect 2363 5475 2389 5501
rect 3911 5475 3937 5501
rect 3963 5475 3989 5501
rect 4015 5475 4041 5501
rect 5563 5475 5589 5501
rect 5615 5475 5641 5501
rect 5667 5475 5693 5501
rect 7215 5475 7241 5501
rect 7267 5475 7293 5501
rect 7319 5475 7345 5501
rect 1433 5083 1459 5109
rect 1485 5083 1511 5109
rect 1537 5083 1563 5109
rect 3085 5083 3111 5109
rect 3137 5083 3163 5109
rect 3189 5083 3215 5109
rect 4737 5083 4763 5109
rect 4789 5083 4815 5109
rect 4841 5083 4867 5109
rect 6389 5083 6415 5109
rect 6441 5083 6467 5109
rect 6493 5083 6519 5109
rect 2259 4691 2285 4717
rect 2311 4691 2337 4717
rect 2363 4691 2389 4717
rect 3911 4691 3937 4717
rect 3963 4691 3989 4717
rect 4015 4691 4041 4717
rect 5563 4691 5589 4717
rect 5615 4691 5641 4717
rect 5667 4691 5693 4717
rect 7215 4691 7241 4717
rect 7267 4691 7293 4717
rect 7319 4691 7345 4717
rect 1433 4299 1459 4325
rect 1485 4299 1511 4325
rect 1537 4299 1563 4325
rect 3085 4299 3111 4325
rect 3137 4299 3163 4325
rect 3189 4299 3215 4325
rect 4737 4299 4763 4325
rect 4789 4299 4815 4325
rect 4841 4299 4867 4325
rect 6389 4299 6415 4325
rect 6441 4299 6467 4325
rect 6493 4299 6519 4325
rect 2259 3907 2285 3933
rect 2311 3907 2337 3933
rect 2363 3907 2389 3933
rect 3911 3907 3937 3933
rect 3963 3907 3989 3933
rect 4015 3907 4041 3933
rect 5563 3907 5589 3933
rect 5615 3907 5641 3933
rect 5667 3907 5693 3933
rect 7215 3907 7241 3933
rect 7267 3907 7293 3933
rect 7319 3907 7345 3933
rect 2367 3823 2393 3849
rect 3487 3823 3513 3849
rect 3991 3823 4017 3849
rect 2367 3711 2393 3737
rect 2535 3711 2561 3737
rect 3375 3711 3401 3737
rect 3487 3711 3513 3737
rect 3599 3711 3625 3737
rect 3935 3711 3961 3737
rect 4159 3711 4185 3737
rect 2423 3599 2449 3625
rect 4047 3599 4073 3625
rect 1433 3515 1459 3541
rect 1485 3515 1511 3541
rect 1537 3515 1563 3541
rect 3085 3515 3111 3541
rect 3137 3515 3163 3541
rect 3189 3515 3215 3541
rect 4737 3515 4763 3541
rect 4789 3515 4815 3541
rect 4841 3515 4867 3541
rect 6389 3515 6415 3541
rect 6441 3515 6467 3541
rect 6493 3515 6519 3541
rect 2199 3431 2225 3457
rect 2871 3319 2897 3345
rect 3151 3319 3177 3345
rect 3487 3319 3513 3345
rect 2479 3263 2505 3289
rect 2255 3207 2281 3233
rect 2367 3207 2393 3233
rect 3095 3207 3121 3233
rect 3207 3207 3233 3233
rect 2259 3123 2285 3149
rect 2311 3123 2337 3149
rect 2363 3123 2389 3149
rect 3911 3123 3937 3149
rect 3963 3123 3989 3149
rect 4015 3123 4041 3149
rect 5563 3123 5589 3149
rect 5615 3123 5641 3149
rect 5667 3123 5693 3149
rect 7215 3123 7241 3149
rect 7267 3123 7293 3149
rect 7319 3123 7345 3149
rect 3823 3039 3849 3065
rect 3879 2983 3905 3009
rect 4103 2983 4129 3009
rect 2591 2927 2617 2953
rect 2815 2927 2841 2953
rect 1433 2731 1459 2757
rect 1485 2731 1511 2757
rect 1537 2731 1563 2757
rect 3085 2731 3111 2757
rect 3137 2731 3163 2757
rect 3189 2731 3215 2757
rect 4737 2731 4763 2757
rect 4789 2731 4815 2757
rect 4841 2731 4867 2757
rect 6389 2731 6415 2757
rect 6441 2731 6467 2757
rect 6493 2731 6519 2757
rect 3263 2591 3289 2617
rect 2087 2535 2113 2561
rect 2255 2535 2281 2561
rect 2143 2479 2169 2505
rect 2367 2479 2393 2505
rect 3039 2479 3065 2505
rect 3151 2479 3177 2505
rect 3319 2479 3345 2505
rect 911 2423 937 2449
rect 2259 2339 2285 2365
rect 2311 2339 2337 2365
rect 2363 2339 2389 2365
rect 3911 2339 3937 2365
rect 3963 2339 3989 2365
rect 4015 2339 4041 2365
rect 5563 2339 5589 2365
rect 5615 2339 5641 2365
rect 5667 2339 5693 2365
rect 7215 2339 7241 2365
rect 7267 2339 7293 2365
rect 7319 2339 7345 2365
rect 2199 2255 2225 2281
rect 2535 2255 2561 2281
rect 2703 2255 2729 2281
rect 3263 2255 3289 2281
rect 3767 2255 3793 2281
rect 2647 2199 2673 2225
rect 3207 2199 3233 2225
rect 1527 2143 1553 2169
rect 2087 2143 2113 2169
rect 2759 2143 2785 2169
rect 2983 2143 3009 2169
rect 3319 2143 3345 2169
rect 3599 2143 3625 2169
rect 3767 2143 3793 2169
rect 3935 2143 3961 2169
rect 967 2087 993 2113
rect 5727 2087 5753 2113
rect 1433 1947 1459 1973
rect 1485 1947 1511 1973
rect 1537 1947 1563 1973
rect 3085 1947 3111 1973
rect 3137 1947 3163 1973
rect 3189 1947 3215 1973
rect 4737 1947 4763 1973
rect 4789 1947 4815 1973
rect 4841 1947 4867 1973
rect 6389 1947 6415 1973
rect 6441 1947 6467 1973
rect 6493 1947 6519 1973
rect 1695 1807 1721 1833
rect 3599 1807 3625 1833
rect 2367 1751 2393 1777
rect 5559 1751 5585 1777
rect 1023 1695 1049 1721
rect 2087 1695 2113 1721
rect 2479 1695 2505 1721
rect 2927 1695 2953 1721
rect 3879 1695 3905 1721
rect 4103 1695 4129 1721
rect 4271 1695 4297 1721
rect 6063 1695 6089 1721
rect 6343 1695 6369 1721
rect 5447 1639 5473 1665
rect 5895 1639 5921 1665
rect 2259 1555 2285 1581
rect 2311 1555 2337 1581
rect 2363 1555 2389 1581
rect 3911 1555 3937 1581
rect 3963 1555 3989 1581
rect 4015 1555 4041 1581
rect 5563 1555 5589 1581
rect 5615 1555 5641 1581
rect 5667 1555 5693 1581
rect 7215 1555 7241 1581
rect 7267 1555 7293 1581
rect 7319 1555 7345 1581
<< metal2 >>
rect 1008 7600 1064 8000
rect 2968 7600 3024 8000
rect 4928 7600 4984 8000
rect 6888 7600 6944 8000
rect 1022 6146 1050 7600
rect 2258 6286 2390 6291
rect 2286 6258 2310 6286
rect 2338 6258 2362 6286
rect 2258 6253 2390 6258
rect 1190 6146 1218 6151
rect 1022 6145 1218 6146
rect 1022 6119 1191 6145
rect 1217 6119 1218 6145
rect 1022 6118 1218 6119
rect 1190 6113 1218 6118
rect 1750 6090 1778 6095
rect 1750 6089 2226 6090
rect 1750 6063 1751 6089
rect 1777 6063 2226 6089
rect 1750 6062 2226 6063
rect 1750 6057 1778 6062
rect 966 5978 994 5983
rect 966 5753 994 5950
rect 1432 5894 1564 5899
rect 1460 5866 1484 5894
rect 1512 5866 1536 5894
rect 1432 5861 1564 5866
rect 966 5727 967 5753
rect 993 5727 994 5753
rect 966 5721 994 5727
rect 1526 5698 1554 5703
rect 1526 5697 1666 5698
rect 1526 5671 1527 5697
rect 1553 5671 1666 5697
rect 1526 5670 1666 5671
rect 1526 5665 1554 5670
rect 1432 5110 1564 5115
rect 1460 5082 1484 5110
rect 1512 5082 1536 5110
rect 1432 5077 1564 5082
rect 1638 4914 1666 5670
rect 1638 4881 1666 4886
rect 1432 4326 1564 4331
rect 1460 4298 1484 4326
rect 1512 4298 1536 4326
rect 1432 4293 1564 4298
rect 1432 3542 1564 3547
rect 1460 3514 1484 3542
rect 1512 3514 1536 3542
rect 1432 3509 1564 3514
rect 2198 3457 2226 6062
rect 2982 6034 3010 7600
rect 3910 6286 4042 6291
rect 3938 6258 3962 6286
rect 3990 6258 4014 6286
rect 3910 6253 4042 6258
rect 3206 6090 3234 6095
rect 3206 6089 3290 6090
rect 3206 6063 3207 6089
rect 3233 6063 3290 6089
rect 3206 6062 3290 6063
rect 3206 6057 3234 6062
rect 2982 6001 3010 6006
rect 3084 5894 3216 5899
rect 3112 5866 3136 5894
rect 3164 5866 3188 5894
rect 3084 5861 3216 5866
rect 2258 5502 2390 5507
rect 2286 5474 2310 5502
rect 2338 5474 2362 5502
rect 2258 5469 2390 5474
rect 3084 5110 3216 5115
rect 3112 5082 3136 5110
rect 3164 5082 3188 5110
rect 3084 5077 3216 5082
rect 2422 4914 2450 4919
rect 2258 4718 2390 4723
rect 2286 4690 2310 4718
rect 2338 4690 2362 4718
rect 2258 4685 2390 4690
rect 2258 3934 2390 3939
rect 2286 3906 2310 3934
rect 2338 3906 2362 3934
rect 2258 3901 2390 3906
rect 2366 3850 2394 3855
rect 2422 3850 2450 4886
rect 3084 4326 3216 4331
rect 3112 4298 3136 4326
rect 3164 4298 3188 4326
rect 3084 4293 3216 4298
rect 2366 3849 2450 3850
rect 2366 3823 2367 3849
rect 2393 3823 2450 3849
rect 2366 3822 2450 3823
rect 2366 3817 2394 3822
rect 2366 3738 2394 3743
rect 2534 3738 2562 3743
rect 2366 3737 2506 3738
rect 2366 3711 2367 3737
rect 2393 3711 2506 3737
rect 2366 3710 2506 3711
rect 2366 3705 2394 3710
rect 2478 3682 2506 3710
rect 2534 3691 2562 3710
rect 2422 3626 2450 3631
rect 2198 3431 2199 3457
rect 2225 3431 2226 3457
rect 2198 3425 2226 3431
rect 2366 3625 2450 3626
rect 2366 3599 2423 3625
rect 2449 3599 2450 3625
rect 2366 3598 2450 3599
rect 2254 3234 2282 3239
rect 2142 3233 2282 3234
rect 2142 3207 2255 3233
rect 2281 3207 2282 3233
rect 2142 3206 2282 3207
rect 2142 2954 2170 3206
rect 2254 3201 2282 3206
rect 2366 3234 2394 3598
rect 2422 3593 2450 3598
rect 2478 3514 2506 3654
rect 2366 3201 2394 3206
rect 2422 3486 2506 3514
rect 3084 3542 3216 3547
rect 3112 3514 3136 3542
rect 3164 3514 3188 3542
rect 3084 3509 3216 3514
rect 2258 3150 2390 3155
rect 2286 3122 2310 3150
rect 2338 3122 2362 3150
rect 2258 3117 2390 3122
rect 1432 2758 1564 2763
rect 1460 2730 1484 2758
rect 1512 2730 1536 2758
rect 1432 2725 1564 2730
rect 1526 2562 1554 2567
rect 910 2449 938 2455
rect 910 2423 911 2449
rect 937 2423 938 2449
rect 910 1722 938 2423
rect 1526 2169 1554 2534
rect 2086 2562 2114 2567
rect 2086 2515 2114 2534
rect 2142 2505 2170 2926
rect 2254 3066 2282 3071
rect 2254 2562 2282 3038
rect 2142 2479 2143 2505
rect 2169 2479 2170 2505
rect 2142 2473 2170 2479
rect 2198 2561 2282 2562
rect 2198 2535 2255 2561
rect 2281 2535 2282 2561
rect 2198 2534 2282 2535
rect 2198 2281 2226 2534
rect 2254 2529 2282 2534
rect 2366 2506 2394 2511
rect 2422 2506 2450 3486
rect 2870 3346 2898 3351
rect 2814 3318 2870 3346
rect 2366 2505 2450 2506
rect 2366 2479 2367 2505
rect 2393 2479 2450 2505
rect 2366 2478 2450 2479
rect 2366 2473 2394 2478
rect 2258 2366 2390 2371
rect 2286 2338 2310 2366
rect 2338 2338 2362 2366
rect 2258 2333 2390 2338
rect 2198 2255 2199 2281
rect 2225 2255 2226 2281
rect 2198 2249 2226 2255
rect 1526 2143 1527 2169
rect 1553 2143 1554 2169
rect 1526 2137 1554 2143
rect 2086 2170 2114 2175
rect 2422 2170 2450 2478
rect 2478 3289 2506 3295
rect 2478 3263 2479 3289
rect 2505 3263 2506 3289
rect 2478 2282 2506 3263
rect 2590 2954 2618 2959
rect 2590 2907 2618 2926
rect 2814 2954 2842 3318
rect 2870 3280 2898 3318
rect 3150 3346 3178 3351
rect 3262 3346 3290 6062
rect 3430 6034 3458 6039
rect 3430 5987 3458 6006
rect 4942 6034 4970 7600
rect 5562 6286 5694 6291
rect 5590 6258 5614 6286
rect 5642 6258 5666 6286
rect 5562 6253 5694 6258
rect 4942 6001 4970 6006
rect 5054 6089 5082 6095
rect 5054 6063 5055 6089
rect 5081 6063 5082 6089
rect 4736 5894 4868 5899
rect 4764 5866 4788 5894
rect 4816 5866 4840 5894
rect 4736 5861 4868 5866
rect 3910 5502 4042 5507
rect 3938 5474 3962 5502
rect 3990 5474 4014 5502
rect 3910 5469 4042 5474
rect 4736 5110 4868 5115
rect 4764 5082 4788 5110
rect 4816 5082 4840 5110
rect 4736 5077 4868 5082
rect 3910 4718 4042 4723
rect 3938 4690 3962 4718
rect 3990 4690 4014 4718
rect 3910 4685 4042 4690
rect 4736 4326 4868 4331
rect 4764 4298 4788 4326
rect 4816 4298 4840 4326
rect 4736 4293 4868 4298
rect 3486 4018 3514 4023
rect 3486 3849 3514 3990
rect 5054 4018 5082 6063
rect 5390 6034 5418 6039
rect 5390 5987 5418 6006
rect 6388 5894 6520 5899
rect 6416 5866 6440 5894
rect 6468 5866 6492 5894
rect 6388 5861 6520 5866
rect 6006 5754 6034 5759
rect 6006 5707 6034 5726
rect 6902 5754 6930 7600
rect 7214 6286 7346 6291
rect 7242 6258 7266 6286
rect 7294 6258 7318 6286
rect 7214 6253 7346 6258
rect 6902 5721 6930 5726
rect 5054 3985 5082 3990
rect 5446 5697 5474 5703
rect 5446 5671 5447 5697
rect 5473 5671 5474 5697
rect 3910 3934 4042 3939
rect 3938 3906 3962 3934
rect 3990 3906 4014 3934
rect 3910 3901 4042 3906
rect 3486 3823 3487 3849
rect 3513 3823 3514 3849
rect 3486 3817 3514 3823
rect 3990 3850 4018 3855
rect 3990 3803 4018 3822
rect 5446 3850 5474 5671
rect 5562 5502 5694 5507
rect 5590 5474 5614 5502
rect 5642 5474 5666 5502
rect 5562 5469 5694 5474
rect 7214 5502 7346 5507
rect 7242 5474 7266 5502
rect 7294 5474 7318 5502
rect 7214 5469 7346 5474
rect 6388 5110 6520 5115
rect 6416 5082 6440 5110
rect 6468 5082 6492 5110
rect 6388 5077 6520 5082
rect 5562 4718 5694 4723
rect 5590 4690 5614 4718
rect 5642 4690 5666 4718
rect 5562 4685 5694 4690
rect 7214 4718 7346 4723
rect 7242 4690 7266 4718
rect 7294 4690 7318 4718
rect 7214 4685 7346 4690
rect 6388 4326 6520 4331
rect 6416 4298 6440 4326
rect 6468 4298 6492 4326
rect 6388 4293 6520 4298
rect 5562 3934 5694 3939
rect 5590 3906 5614 3934
rect 5642 3906 5666 3934
rect 5562 3901 5694 3906
rect 7214 3934 7346 3939
rect 7242 3906 7266 3934
rect 7294 3906 7318 3934
rect 7214 3901 7346 3906
rect 5446 3817 5474 3822
rect 3150 3345 3290 3346
rect 3150 3319 3151 3345
rect 3177 3319 3290 3345
rect 3150 3318 3290 3319
rect 3374 3737 3402 3743
rect 3374 3711 3375 3737
rect 3401 3711 3402 3737
rect 3150 3313 3178 3318
rect 3094 3234 3122 3239
rect 3094 3187 3122 3206
rect 3206 3234 3234 3239
rect 3206 3233 3290 3234
rect 3206 3207 3207 3233
rect 3233 3207 3290 3233
rect 3206 3206 3290 3207
rect 3206 3201 3234 3206
rect 2814 2907 2842 2926
rect 3084 2758 3216 2763
rect 3112 2730 3136 2758
rect 3164 2730 3188 2758
rect 3084 2725 3216 2730
rect 3262 2617 3290 3206
rect 3262 2591 3263 2617
rect 3289 2591 3290 2617
rect 3262 2585 3290 2591
rect 3374 2562 3402 3711
rect 3486 3737 3514 3743
rect 3486 3711 3487 3737
rect 3513 3711 3514 3737
rect 3486 3682 3514 3711
rect 3598 3738 3626 3743
rect 3934 3738 3962 3743
rect 3598 3691 3626 3710
rect 3766 3737 3962 3738
rect 3766 3711 3935 3737
rect 3961 3711 3962 3737
rect 3766 3710 3962 3711
rect 3486 3649 3514 3654
rect 3486 3346 3514 3351
rect 3486 3010 3514 3318
rect 3486 2977 3514 2982
rect 3374 2529 3402 2534
rect 2478 2249 2506 2254
rect 2534 2506 2562 2511
rect 2534 2281 2562 2478
rect 3038 2506 3066 2511
rect 3038 2459 3066 2478
rect 3150 2506 3178 2511
rect 3150 2505 3234 2506
rect 3150 2479 3151 2505
rect 3177 2479 3234 2505
rect 3150 2478 3234 2479
rect 3150 2473 3178 2478
rect 2534 2255 2535 2281
rect 2561 2255 2562 2281
rect 2422 2142 2506 2170
rect 2086 2123 2114 2142
rect 966 2113 994 2119
rect 966 2087 967 2113
rect 993 2087 994 2113
rect 966 2002 994 2087
rect 966 1969 994 1974
rect 1432 1974 1564 1979
rect 1460 1946 1484 1974
rect 1512 1946 1536 1974
rect 1432 1941 1564 1946
rect 1694 1833 1722 1839
rect 1694 1807 1695 1833
rect 1721 1807 1722 1833
rect 1694 1778 1722 1807
rect 1694 1745 1722 1750
rect 2366 1778 2394 1783
rect 2366 1731 2394 1750
rect 1022 1722 1050 1727
rect 854 1721 1050 1722
rect 854 1695 1023 1721
rect 1049 1695 1050 1721
rect 854 1694 1050 1695
rect 854 400 882 1694
rect 1022 1689 1050 1694
rect 2086 1722 2114 1727
rect 840 0 896 400
rect 2086 378 2114 1694
rect 2478 1721 2506 2142
rect 2534 1778 2562 2255
rect 2702 2282 2730 2287
rect 2702 2235 2730 2254
rect 2646 2226 2674 2231
rect 2646 2179 2674 2198
rect 3206 2226 3234 2478
rect 3318 2505 3346 2511
rect 3318 2479 3319 2505
rect 3345 2479 3346 2505
rect 3262 2394 3290 2399
rect 3262 2281 3290 2366
rect 3262 2255 3263 2281
rect 3289 2255 3290 2281
rect 3262 2249 3290 2255
rect 3206 2179 3234 2198
rect 2758 2169 2786 2175
rect 2758 2143 2759 2169
rect 2785 2143 2786 2169
rect 2758 2114 2786 2143
rect 2982 2170 3010 2175
rect 2982 2123 3010 2142
rect 3318 2169 3346 2479
rect 3766 2281 3794 3710
rect 3934 3705 3962 3710
rect 4158 3738 4186 3743
rect 4158 3691 4186 3710
rect 3822 3626 3850 3631
rect 3822 3065 3850 3598
rect 4046 3625 4074 3631
rect 4046 3599 4047 3625
rect 4073 3599 4074 3625
rect 4046 3570 4074 3599
rect 4046 3537 4074 3542
rect 4736 3542 4868 3547
rect 4764 3514 4788 3542
rect 4816 3514 4840 3542
rect 4736 3509 4868 3514
rect 6388 3542 6520 3547
rect 6416 3514 6440 3542
rect 6468 3514 6492 3542
rect 6388 3509 6520 3514
rect 3910 3150 4042 3155
rect 3938 3122 3962 3150
rect 3990 3122 4014 3150
rect 3910 3117 4042 3122
rect 5562 3150 5694 3155
rect 5590 3122 5614 3150
rect 5642 3122 5666 3150
rect 5562 3117 5694 3122
rect 7214 3150 7346 3155
rect 7242 3122 7266 3150
rect 7294 3122 7318 3150
rect 7214 3117 7346 3122
rect 3822 3039 3823 3065
rect 3849 3039 3850 3065
rect 3822 3033 3850 3039
rect 3878 3010 3906 3015
rect 3878 2963 3906 2982
rect 4102 3010 4130 3015
rect 4102 2963 4130 2982
rect 5894 2898 5922 2903
rect 4736 2758 4868 2763
rect 4764 2730 4788 2758
rect 4816 2730 4840 2758
rect 4736 2725 4868 2730
rect 3910 2366 4042 2371
rect 3938 2338 3962 2366
rect 3990 2338 4014 2366
rect 3910 2333 4042 2338
rect 5562 2366 5694 2371
rect 5590 2338 5614 2366
rect 5642 2338 5666 2366
rect 5562 2333 5694 2338
rect 3766 2255 3767 2281
rect 3793 2255 3794 2281
rect 3766 2249 3794 2255
rect 3318 2143 3319 2169
rect 3345 2143 3346 2169
rect 2758 2081 2786 2086
rect 3318 2114 3346 2143
rect 3318 2081 3346 2086
rect 3598 2170 3626 2175
rect 3084 1974 3216 1979
rect 3112 1946 3136 1974
rect 3164 1946 3188 1974
rect 3084 1941 3216 1946
rect 3598 1833 3626 2142
rect 3766 2170 3794 2175
rect 3766 2123 3794 2142
rect 3934 2169 3962 2175
rect 3934 2143 3935 2169
rect 3961 2143 3962 2169
rect 3934 2114 3962 2143
rect 3934 2081 3962 2086
rect 4102 2170 4130 2175
rect 3598 1807 3599 1833
rect 3625 1807 3626 1833
rect 3598 1801 3626 1807
rect 2534 1745 2562 1750
rect 2478 1695 2479 1721
rect 2505 1695 2506 1721
rect 2478 1689 2506 1695
rect 2926 1722 2954 1727
rect 3878 1722 3906 1727
rect 2926 1675 2954 1694
rect 3822 1694 3878 1722
rect 2258 1582 2390 1587
rect 2286 1554 2310 1582
rect 2338 1554 2362 1582
rect 2258 1549 2390 1554
rect 3822 1106 3850 1694
rect 3878 1656 3906 1694
rect 4102 1721 4130 2142
rect 5446 2114 5474 2119
rect 4736 1974 4868 1979
rect 4764 1946 4788 1974
rect 4816 1946 4840 1974
rect 4736 1941 4868 1946
rect 4102 1695 4103 1721
rect 4129 1695 4130 1721
rect 4102 1689 4130 1695
rect 4270 1722 4298 1727
rect 4270 1675 4298 1694
rect 5446 1665 5474 2086
rect 5726 2113 5754 2119
rect 5726 2087 5727 2113
rect 5753 2087 5754 2113
rect 5558 1778 5586 1783
rect 5726 1778 5754 2087
rect 5446 1639 5447 1665
rect 5473 1639 5474 1665
rect 5446 1633 5474 1639
rect 5502 1777 5754 1778
rect 5502 1751 5559 1777
rect 5585 1751 5754 1777
rect 5502 1750 5754 1751
rect 3910 1582 4042 1587
rect 3938 1554 3962 1582
rect 3990 1554 4014 1582
rect 3910 1549 4042 1554
rect 5502 1274 5530 1750
rect 5558 1745 5586 1750
rect 5894 1665 5922 2870
rect 6388 2758 6520 2763
rect 6416 2730 6440 2758
rect 6468 2730 6492 2758
rect 6388 2725 6520 2730
rect 7214 2366 7346 2371
rect 7242 2338 7266 2366
rect 7294 2338 7318 2366
rect 7214 2333 7346 2338
rect 6388 1974 6520 1979
rect 6416 1946 6440 1974
rect 6468 1946 6492 1974
rect 6388 1941 6520 1946
rect 6062 1722 6090 1727
rect 6062 1675 6090 1694
rect 6342 1722 6370 1727
rect 6342 1675 6370 1694
rect 7126 1722 7154 1727
rect 5894 1639 5895 1665
rect 5921 1639 5922 1665
rect 5894 1633 5922 1639
rect 5562 1582 5694 1587
rect 5590 1554 5614 1582
rect 5642 1554 5666 1582
rect 5562 1549 5694 1554
rect 5502 1246 5586 1274
rect 3822 1078 4018 1106
rect 2254 462 2450 490
rect 2254 378 2282 462
rect 2422 400 2450 462
rect 3990 400 4018 1078
rect 5558 400 5586 1246
rect 7126 400 7154 1694
rect 7214 1582 7346 1587
rect 7242 1554 7266 1582
rect 7294 1554 7318 1582
rect 7214 1549 7346 1554
rect 2086 350 2282 378
rect 2408 0 2464 400
rect 3976 0 4032 400
rect 5544 0 5600 400
rect 7112 0 7168 400
<< via2 >>
rect 2258 6285 2286 6286
rect 2258 6259 2259 6285
rect 2259 6259 2285 6285
rect 2285 6259 2286 6285
rect 2258 6258 2286 6259
rect 2310 6285 2338 6286
rect 2310 6259 2311 6285
rect 2311 6259 2337 6285
rect 2337 6259 2338 6285
rect 2310 6258 2338 6259
rect 2362 6285 2390 6286
rect 2362 6259 2363 6285
rect 2363 6259 2389 6285
rect 2389 6259 2390 6285
rect 2362 6258 2390 6259
rect 966 5950 994 5978
rect 1432 5893 1460 5894
rect 1432 5867 1433 5893
rect 1433 5867 1459 5893
rect 1459 5867 1460 5893
rect 1432 5866 1460 5867
rect 1484 5893 1512 5894
rect 1484 5867 1485 5893
rect 1485 5867 1511 5893
rect 1511 5867 1512 5893
rect 1484 5866 1512 5867
rect 1536 5893 1564 5894
rect 1536 5867 1537 5893
rect 1537 5867 1563 5893
rect 1563 5867 1564 5893
rect 1536 5866 1564 5867
rect 1432 5109 1460 5110
rect 1432 5083 1433 5109
rect 1433 5083 1459 5109
rect 1459 5083 1460 5109
rect 1432 5082 1460 5083
rect 1484 5109 1512 5110
rect 1484 5083 1485 5109
rect 1485 5083 1511 5109
rect 1511 5083 1512 5109
rect 1484 5082 1512 5083
rect 1536 5109 1564 5110
rect 1536 5083 1537 5109
rect 1537 5083 1563 5109
rect 1563 5083 1564 5109
rect 1536 5082 1564 5083
rect 1638 4886 1666 4914
rect 1432 4325 1460 4326
rect 1432 4299 1433 4325
rect 1433 4299 1459 4325
rect 1459 4299 1460 4325
rect 1432 4298 1460 4299
rect 1484 4325 1512 4326
rect 1484 4299 1485 4325
rect 1485 4299 1511 4325
rect 1511 4299 1512 4325
rect 1484 4298 1512 4299
rect 1536 4325 1564 4326
rect 1536 4299 1537 4325
rect 1537 4299 1563 4325
rect 1563 4299 1564 4325
rect 1536 4298 1564 4299
rect 1432 3541 1460 3542
rect 1432 3515 1433 3541
rect 1433 3515 1459 3541
rect 1459 3515 1460 3541
rect 1432 3514 1460 3515
rect 1484 3541 1512 3542
rect 1484 3515 1485 3541
rect 1485 3515 1511 3541
rect 1511 3515 1512 3541
rect 1484 3514 1512 3515
rect 1536 3541 1564 3542
rect 1536 3515 1537 3541
rect 1537 3515 1563 3541
rect 1563 3515 1564 3541
rect 1536 3514 1564 3515
rect 3910 6285 3938 6286
rect 3910 6259 3911 6285
rect 3911 6259 3937 6285
rect 3937 6259 3938 6285
rect 3910 6258 3938 6259
rect 3962 6285 3990 6286
rect 3962 6259 3963 6285
rect 3963 6259 3989 6285
rect 3989 6259 3990 6285
rect 3962 6258 3990 6259
rect 4014 6285 4042 6286
rect 4014 6259 4015 6285
rect 4015 6259 4041 6285
rect 4041 6259 4042 6285
rect 4014 6258 4042 6259
rect 2982 6006 3010 6034
rect 3084 5893 3112 5894
rect 3084 5867 3085 5893
rect 3085 5867 3111 5893
rect 3111 5867 3112 5893
rect 3084 5866 3112 5867
rect 3136 5893 3164 5894
rect 3136 5867 3137 5893
rect 3137 5867 3163 5893
rect 3163 5867 3164 5893
rect 3136 5866 3164 5867
rect 3188 5893 3216 5894
rect 3188 5867 3189 5893
rect 3189 5867 3215 5893
rect 3215 5867 3216 5893
rect 3188 5866 3216 5867
rect 2258 5501 2286 5502
rect 2258 5475 2259 5501
rect 2259 5475 2285 5501
rect 2285 5475 2286 5501
rect 2258 5474 2286 5475
rect 2310 5501 2338 5502
rect 2310 5475 2311 5501
rect 2311 5475 2337 5501
rect 2337 5475 2338 5501
rect 2310 5474 2338 5475
rect 2362 5501 2390 5502
rect 2362 5475 2363 5501
rect 2363 5475 2389 5501
rect 2389 5475 2390 5501
rect 2362 5474 2390 5475
rect 3084 5109 3112 5110
rect 3084 5083 3085 5109
rect 3085 5083 3111 5109
rect 3111 5083 3112 5109
rect 3084 5082 3112 5083
rect 3136 5109 3164 5110
rect 3136 5083 3137 5109
rect 3137 5083 3163 5109
rect 3163 5083 3164 5109
rect 3136 5082 3164 5083
rect 3188 5109 3216 5110
rect 3188 5083 3189 5109
rect 3189 5083 3215 5109
rect 3215 5083 3216 5109
rect 3188 5082 3216 5083
rect 2422 4886 2450 4914
rect 2258 4717 2286 4718
rect 2258 4691 2259 4717
rect 2259 4691 2285 4717
rect 2285 4691 2286 4717
rect 2258 4690 2286 4691
rect 2310 4717 2338 4718
rect 2310 4691 2311 4717
rect 2311 4691 2337 4717
rect 2337 4691 2338 4717
rect 2310 4690 2338 4691
rect 2362 4717 2390 4718
rect 2362 4691 2363 4717
rect 2363 4691 2389 4717
rect 2389 4691 2390 4717
rect 2362 4690 2390 4691
rect 2258 3933 2286 3934
rect 2258 3907 2259 3933
rect 2259 3907 2285 3933
rect 2285 3907 2286 3933
rect 2258 3906 2286 3907
rect 2310 3933 2338 3934
rect 2310 3907 2311 3933
rect 2311 3907 2337 3933
rect 2337 3907 2338 3933
rect 2310 3906 2338 3907
rect 2362 3933 2390 3934
rect 2362 3907 2363 3933
rect 2363 3907 2389 3933
rect 2389 3907 2390 3933
rect 2362 3906 2390 3907
rect 3084 4325 3112 4326
rect 3084 4299 3085 4325
rect 3085 4299 3111 4325
rect 3111 4299 3112 4325
rect 3084 4298 3112 4299
rect 3136 4325 3164 4326
rect 3136 4299 3137 4325
rect 3137 4299 3163 4325
rect 3163 4299 3164 4325
rect 3136 4298 3164 4299
rect 3188 4325 3216 4326
rect 3188 4299 3189 4325
rect 3189 4299 3215 4325
rect 3215 4299 3216 4325
rect 3188 4298 3216 4299
rect 2534 3737 2562 3738
rect 2534 3711 2535 3737
rect 2535 3711 2561 3737
rect 2561 3711 2562 3737
rect 2534 3710 2562 3711
rect 2478 3654 2506 3682
rect 2366 3233 2394 3234
rect 2366 3207 2367 3233
rect 2367 3207 2393 3233
rect 2393 3207 2394 3233
rect 2366 3206 2394 3207
rect 3084 3541 3112 3542
rect 3084 3515 3085 3541
rect 3085 3515 3111 3541
rect 3111 3515 3112 3541
rect 3084 3514 3112 3515
rect 3136 3541 3164 3542
rect 3136 3515 3137 3541
rect 3137 3515 3163 3541
rect 3163 3515 3164 3541
rect 3136 3514 3164 3515
rect 3188 3541 3216 3542
rect 3188 3515 3189 3541
rect 3189 3515 3215 3541
rect 3215 3515 3216 3541
rect 3188 3514 3216 3515
rect 2258 3149 2286 3150
rect 2258 3123 2259 3149
rect 2259 3123 2285 3149
rect 2285 3123 2286 3149
rect 2258 3122 2286 3123
rect 2310 3149 2338 3150
rect 2310 3123 2311 3149
rect 2311 3123 2337 3149
rect 2337 3123 2338 3149
rect 2310 3122 2338 3123
rect 2362 3149 2390 3150
rect 2362 3123 2363 3149
rect 2363 3123 2389 3149
rect 2389 3123 2390 3149
rect 2362 3122 2390 3123
rect 2142 2926 2170 2954
rect 1432 2757 1460 2758
rect 1432 2731 1433 2757
rect 1433 2731 1459 2757
rect 1459 2731 1460 2757
rect 1432 2730 1460 2731
rect 1484 2757 1512 2758
rect 1484 2731 1485 2757
rect 1485 2731 1511 2757
rect 1511 2731 1512 2757
rect 1484 2730 1512 2731
rect 1536 2757 1564 2758
rect 1536 2731 1537 2757
rect 1537 2731 1563 2757
rect 1563 2731 1564 2757
rect 1536 2730 1564 2731
rect 1526 2534 1554 2562
rect 2086 2561 2114 2562
rect 2086 2535 2087 2561
rect 2087 2535 2113 2561
rect 2113 2535 2114 2561
rect 2086 2534 2114 2535
rect 2254 3038 2282 3066
rect 2870 3345 2898 3346
rect 2870 3319 2871 3345
rect 2871 3319 2897 3345
rect 2897 3319 2898 3345
rect 2870 3318 2898 3319
rect 2258 2365 2286 2366
rect 2258 2339 2259 2365
rect 2259 2339 2285 2365
rect 2285 2339 2286 2365
rect 2258 2338 2286 2339
rect 2310 2365 2338 2366
rect 2310 2339 2311 2365
rect 2311 2339 2337 2365
rect 2337 2339 2338 2365
rect 2310 2338 2338 2339
rect 2362 2365 2390 2366
rect 2362 2339 2363 2365
rect 2363 2339 2389 2365
rect 2389 2339 2390 2365
rect 2362 2338 2390 2339
rect 2086 2169 2114 2170
rect 2086 2143 2087 2169
rect 2087 2143 2113 2169
rect 2113 2143 2114 2169
rect 2086 2142 2114 2143
rect 2590 2953 2618 2954
rect 2590 2927 2591 2953
rect 2591 2927 2617 2953
rect 2617 2927 2618 2953
rect 2590 2926 2618 2927
rect 3430 6033 3458 6034
rect 3430 6007 3431 6033
rect 3431 6007 3457 6033
rect 3457 6007 3458 6033
rect 3430 6006 3458 6007
rect 5562 6285 5590 6286
rect 5562 6259 5563 6285
rect 5563 6259 5589 6285
rect 5589 6259 5590 6285
rect 5562 6258 5590 6259
rect 5614 6285 5642 6286
rect 5614 6259 5615 6285
rect 5615 6259 5641 6285
rect 5641 6259 5642 6285
rect 5614 6258 5642 6259
rect 5666 6285 5694 6286
rect 5666 6259 5667 6285
rect 5667 6259 5693 6285
rect 5693 6259 5694 6285
rect 5666 6258 5694 6259
rect 4942 6006 4970 6034
rect 4736 5893 4764 5894
rect 4736 5867 4737 5893
rect 4737 5867 4763 5893
rect 4763 5867 4764 5893
rect 4736 5866 4764 5867
rect 4788 5893 4816 5894
rect 4788 5867 4789 5893
rect 4789 5867 4815 5893
rect 4815 5867 4816 5893
rect 4788 5866 4816 5867
rect 4840 5893 4868 5894
rect 4840 5867 4841 5893
rect 4841 5867 4867 5893
rect 4867 5867 4868 5893
rect 4840 5866 4868 5867
rect 3910 5501 3938 5502
rect 3910 5475 3911 5501
rect 3911 5475 3937 5501
rect 3937 5475 3938 5501
rect 3910 5474 3938 5475
rect 3962 5501 3990 5502
rect 3962 5475 3963 5501
rect 3963 5475 3989 5501
rect 3989 5475 3990 5501
rect 3962 5474 3990 5475
rect 4014 5501 4042 5502
rect 4014 5475 4015 5501
rect 4015 5475 4041 5501
rect 4041 5475 4042 5501
rect 4014 5474 4042 5475
rect 4736 5109 4764 5110
rect 4736 5083 4737 5109
rect 4737 5083 4763 5109
rect 4763 5083 4764 5109
rect 4736 5082 4764 5083
rect 4788 5109 4816 5110
rect 4788 5083 4789 5109
rect 4789 5083 4815 5109
rect 4815 5083 4816 5109
rect 4788 5082 4816 5083
rect 4840 5109 4868 5110
rect 4840 5083 4841 5109
rect 4841 5083 4867 5109
rect 4867 5083 4868 5109
rect 4840 5082 4868 5083
rect 3910 4717 3938 4718
rect 3910 4691 3911 4717
rect 3911 4691 3937 4717
rect 3937 4691 3938 4717
rect 3910 4690 3938 4691
rect 3962 4717 3990 4718
rect 3962 4691 3963 4717
rect 3963 4691 3989 4717
rect 3989 4691 3990 4717
rect 3962 4690 3990 4691
rect 4014 4717 4042 4718
rect 4014 4691 4015 4717
rect 4015 4691 4041 4717
rect 4041 4691 4042 4717
rect 4014 4690 4042 4691
rect 4736 4325 4764 4326
rect 4736 4299 4737 4325
rect 4737 4299 4763 4325
rect 4763 4299 4764 4325
rect 4736 4298 4764 4299
rect 4788 4325 4816 4326
rect 4788 4299 4789 4325
rect 4789 4299 4815 4325
rect 4815 4299 4816 4325
rect 4788 4298 4816 4299
rect 4840 4325 4868 4326
rect 4840 4299 4841 4325
rect 4841 4299 4867 4325
rect 4867 4299 4868 4325
rect 4840 4298 4868 4299
rect 3486 3990 3514 4018
rect 5390 6033 5418 6034
rect 5390 6007 5391 6033
rect 5391 6007 5417 6033
rect 5417 6007 5418 6033
rect 5390 6006 5418 6007
rect 6388 5893 6416 5894
rect 6388 5867 6389 5893
rect 6389 5867 6415 5893
rect 6415 5867 6416 5893
rect 6388 5866 6416 5867
rect 6440 5893 6468 5894
rect 6440 5867 6441 5893
rect 6441 5867 6467 5893
rect 6467 5867 6468 5893
rect 6440 5866 6468 5867
rect 6492 5893 6520 5894
rect 6492 5867 6493 5893
rect 6493 5867 6519 5893
rect 6519 5867 6520 5893
rect 6492 5866 6520 5867
rect 6006 5753 6034 5754
rect 6006 5727 6007 5753
rect 6007 5727 6033 5753
rect 6033 5727 6034 5753
rect 6006 5726 6034 5727
rect 7214 6285 7242 6286
rect 7214 6259 7215 6285
rect 7215 6259 7241 6285
rect 7241 6259 7242 6285
rect 7214 6258 7242 6259
rect 7266 6285 7294 6286
rect 7266 6259 7267 6285
rect 7267 6259 7293 6285
rect 7293 6259 7294 6285
rect 7266 6258 7294 6259
rect 7318 6285 7346 6286
rect 7318 6259 7319 6285
rect 7319 6259 7345 6285
rect 7345 6259 7346 6285
rect 7318 6258 7346 6259
rect 6902 5726 6930 5754
rect 5054 3990 5082 4018
rect 3910 3933 3938 3934
rect 3910 3907 3911 3933
rect 3911 3907 3937 3933
rect 3937 3907 3938 3933
rect 3910 3906 3938 3907
rect 3962 3933 3990 3934
rect 3962 3907 3963 3933
rect 3963 3907 3989 3933
rect 3989 3907 3990 3933
rect 3962 3906 3990 3907
rect 4014 3933 4042 3934
rect 4014 3907 4015 3933
rect 4015 3907 4041 3933
rect 4041 3907 4042 3933
rect 4014 3906 4042 3907
rect 3990 3849 4018 3850
rect 3990 3823 3991 3849
rect 3991 3823 4017 3849
rect 4017 3823 4018 3849
rect 3990 3822 4018 3823
rect 5562 5501 5590 5502
rect 5562 5475 5563 5501
rect 5563 5475 5589 5501
rect 5589 5475 5590 5501
rect 5562 5474 5590 5475
rect 5614 5501 5642 5502
rect 5614 5475 5615 5501
rect 5615 5475 5641 5501
rect 5641 5475 5642 5501
rect 5614 5474 5642 5475
rect 5666 5501 5694 5502
rect 5666 5475 5667 5501
rect 5667 5475 5693 5501
rect 5693 5475 5694 5501
rect 5666 5474 5694 5475
rect 7214 5501 7242 5502
rect 7214 5475 7215 5501
rect 7215 5475 7241 5501
rect 7241 5475 7242 5501
rect 7214 5474 7242 5475
rect 7266 5501 7294 5502
rect 7266 5475 7267 5501
rect 7267 5475 7293 5501
rect 7293 5475 7294 5501
rect 7266 5474 7294 5475
rect 7318 5501 7346 5502
rect 7318 5475 7319 5501
rect 7319 5475 7345 5501
rect 7345 5475 7346 5501
rect 7318 5474 7346 5475
rect 6388 5109 6416 5110
rect 6388 5083 6389 5109
rect 6389 5083 6415 5109
rect 6415 5083 6416 5109
rect 6388 5082 6416 5083
rect 6440 5109 6468 5110
rect 6440 5083 6441 5109
rect 6441 5083 6467 5109
rect 6467 5083 6468 5109
rect 6440 5082 6468 5083
rect 6492 5109 6520 5110
rect 6492 5083 6493 5109
rect 6493 5083 6519 5109
rect 6519 5083 6520 5109
rect 6492 5082 6520 5083
rect 5562 4717 5590 4718
rect 5562 4691 5563 4717
rect 5563 4691 5589 4717
rect 5589 4691 5590 4717
rect 5562 4690 5590 4691
rect 5614 4717 5642 4718
rect 5614 4691 5615 4717
rect 5615 4691 5641 4717
rect 5641 4691 5642 4717
rect 5614 4690 5642 4691
rect 5666 4717 5694 4718
rect 5666 4691 5667 4717
rect 5667 4691 5693 4717
rect 5693 4691 5694 4717
rect 5666 4690 5694 4691
rect 7214 4717 7242 4718
rect 7214 4691 7215 4717
rect 7215 4691 7241 4717
rect 7241 4691 7242 4717
rect 7214 4690 7242 4691
rect 7266 4717 7294 4718
rect 7266 4691 7267 4717
rect 7267 4691 7293 4717
rect 7293 4691 7294 4717
rect 7266 4690 7294 4691
rect 7318 4717 7346 4718
rect 7318 4691 7319 4717
rect 7319 4691 7345 4717
rect 7345 4691 7346 4717
rect 7318 4690 7346 4691
rect 6388 4325 6416 4326
rect 6388 4299 6389 4325
rect 6389 4299 6415 4325
rect 6415 4299 6416 4325
rect 6388 4298 6416 4299
rect 6440 4325 6468 4326
rect 6440 4299 6441 4325
rect 6441 4299 6467 4325
rect 6467 4299 6468 4325
rect 6440 4298 6468 4299
rect 6492 4325 6520 4326
rect 6492 4299 6493 4325
rect 6493 4299 6519 4325
rect 6519 4299 6520 4325
rect 6492 4298 6520 4299
rect 5562 3933 5590 3934
rect 5562 3907 5563 3933
rect 5563 3907 5589 3933
rect 5589 3907 5590 3933
rect 5562 3906 5590 3907
rect 5614 3933 5642 3934
rect 5614 3907 5615 3933
rect 5615 3907 5641 3933
rect 5641 3907 5642 3933
rect 5614 3906 5642 3907
rect 5666 3933 5694 3934
rect 5666 3907 5667 3933
rect 5667 3907 5693 3933
rect 5693 3907 5694 3933
rect 5666 3906 5694 3907
rect 7214 3933 7242 3934
rect 7214 3907 7215 3933
rect 7215 3907 7241 3933
rect 7241 3907 7242 3933
rect 7214 3906 7242 3907
rect 7266 3933 7294 3934
rect 7266 3907 7267 3933
rect 7267 3907 7293 3933
rect 7293 3907 7294 3933
rect 7266 3906 7294 3907
rect 7318 3933 7346 3934
rect 7318 3907 7319 3933
rect 7319 3907 7345 3933
rect 7345 3907 7346 3933
rect 7318 3906 7346 3907
rect 5446 3822 5474 3850
rect 3094 3233 3122 3234
rect 3094 3207 3095 3233
rect 3095 3207 3121 3233
rect 3121 3207 3122 3233
rect 3094 3206 3122 3207
rect 2814 2953 2842 2954
rect 2814 2927 2815 2953
rect 2815 2927 2841 2953
rect 2841 2927 2842 2953
rect 2814 2926 2842 2927
rect 3084 2757 3112 2758
rect 3084 2731 3085 2757
rect 3085 2731 3111 2757
rect 3111 2731 3112 2757
rect 3084 2730 3112 2731
rect 3136 2757 3164 2758
rect 3136 2731 3137 2757
rect 3137 2731 3163 2757
rect 3163 2731 3164 2757
rect 3136 2730 3164 2731
rect 3188 2757 3216 2758
rect 3188 2731 3189 2757
rect 3189 2731 3215 2757
rect 3215 2731 3216 2757
rect 3188 2730 3216 2731
rect 3598 3737 3626 3738
rect 3598 3711 3599 3737
rect 3599 3711 3625 3737
rect 3625 3711 3626 3737
rect 3598 3710 3626 3711
rect 3486 3654 3514 3682
rect 3486 3345 3514 3346
rect 3486 3319 3487 3345
rect 3487 3319 3513 3345
rect 3513 3319 3514 3345
rect 3486 3318 3514 3319
rect 3486 2982 3514 3010
rect 3374 2534 3402 2562
rect 2478 2254 2506 2282
rect 2534 2478 2562 2506
rect 3038 2505 3066 2506
rect 3038 2479 3039 2505
rect 3039 2479 3065 2505
rect 3065 2479 3066 2505
rect 3038 2478 3066 2479
rect 966 1974 994 2002
rect 1432 1973 1460 1974
rect 1432 1947 1433 1973
rect 1433 1947 1459 1973
rect 1459 1947 1460 1973
rect 1432 1946 1460 1947
rect 1484 1973 1512 1974
rect 1484 1947 1485 1973
rect 1485 1947 1511 1973
rect 1511 1947 1512 1973
rect 1484 1946 1512 1947
rect 1536 1973 1564 1974
rect 1536 1947 1537 1973
rect 1537 1947 1563 1973
rect 1563 1947 1564 1973
rect 1536 1946 1564 1947
rect 1694 1750 1722 1778
rect 2366 1777 2394 1778
rect 2366 1751 2367 1777
rect 2367 1751 2393 1777
rect 2393 1751 2394 1777
rect 2366 1750 2394 1751
rect 2086 1721 2114 1722
rect 2086 1695 2087 1721
rect 2087 1695 2113 1721
rect 2113 1695 2114 1721
rect 2086 1694 2114 1695
rect 2702 2281 2730 2282
rect 2702 2255 2703 2281
rect 2703 2255 2729 2281
rect 2729 2255 2730 2281
rect 2702 2254 2730 2255
rect 2646 2225 2674 2226
rect 2646 2199 2647 2225
rect 2647 2199 2673 2225
rect 2673 2199 2674 2225
rect 2646 2198 2674 2199
rect 3262 2366 3290 2394
rect 3206 2225 3234 2226
rect 3206 2199 3207 2225
rect 3207 2199 3233 2225
rect 3233 2199 3234 2225
rect 3206 2198 3234 2199
rect 2982 2169 3010 2170
rect 2982 2143 2983 2169
rect 2983 2143 3009 2169
rect 3009 2143 3010 2169
rect 2982 2142 3010 2143
rect 4158 3737 4186 3738
rect 4158 3711 4159 3737
rect 4159 3711 4185 3737
rect 4185 3711 4186 3737
rect 4158 3710 4186 3711
rect 3822 3598 3850 3626
rect 4046 3542 4074 3570
rect 4736 3541 4764 3542
rect 4736 3515 4737 3541
rect 4737 3515 4763 3541
rect 4763 3515 4764 3541
rect 4736 3514 4764 3515
rect 4788 3541 4816 3542
rect 4788 3515 4789 3541
rect 4789 3515 4815 3541
rect 4815 3515 4816 3541
rect 4788 3514 4816 3515
rect 4840 3541 4868 3542
rect 4840 3515 4841 3541
rect 4841 3515 4867 3541
rect 4867 3515 4868 3541
rect 4840 3514 4868 3515
rect 6388 3541 6416 3542
rect 6388 3515 6389 3541
rect 6389 3515 6415 3541
rect 6415 3515 6416 3541
rect 6388 3514 6416 3515
rect 6440 3541 6468 3542
rect 6440 3515 6441 3541
rect 6441 3515 6467 3541
rect 6467 3515 6468 3541
rect 6440 3514 6468 3515
rect 6492 3541 6520 3542
rect 6492 3515 6493 3541
rect 6493 3515 6519 3541
rect 6519 3515 6520 3541
rect 6492 3514 6520 3515
rect 3910 3149 3938 3150
rect 3910 3123 3911 3149
rect 3911 3123 3937 3149
rect 3937 3123 3938 3149
rect 3910 3122 3938 3123
rect 3962 3149 3990 3150
rect 3962 3123 3963 3149
rect 3963 3123 3989 3149
rect 3989 3123 3990 3149
rect 3962 3122 3990 3123
rect 4014 3149 4042 3150
rect 4014 3123 4015 3149
rect 4015 3123 4041 3149
rect 4041 3123 4042 3149
rect 4014 3122 4042 3123
rect 5562 3149 5590 3150
rect 5562 3123 5563 3149
rect 5563 3123 5589 3149
rect 5589 3123 5590 3149
rect 5562 3122 5590 3123
rect 5614 3149 5642 3150
rect 5614 3123 5615 3149
rect 5615 3123 5641 3149
rect 5641 3123 5642 3149
rect 5614 3122 5642 3123
rect 5666 3149 5694 3150
rect 5666 3123 5667 3149
rect 5667 3123 5693 3149
rect 5693 3123 5694 3149
rect 5666 3122 5694 3123
rect 7214 3149 7242 3150
rect 7214 3123 7215 3149
rect 7215 3123 7241 3149
rect 7241 3123 7242 3149
rect 7214 3122 7242 3123
rect 7266 3149 7294 3150
rect 7266 3123 7267 3149
rect 7267 3123 7293 3149
rect 7293 3123 7294 3149
rect 7266 3122 7294 3123
rect 7318 3149 7346 3150
rect 7318 3123 7319 3149
rect 7319 3123 7345 3149
rect 7345 3123 7346 3149
rect 7318 3122 7346 3123
rect 3878 3009 3906 3010
rect 3878 2983 3879 3009
rect 3879 2983 3905 3009
rect 3905 2983 3906 3009
rect 3878 2982 3906 2983
rect 4102 3009 4130 3010
rect 4102 2983 4103 3009
rect 4103 2983 4129 3009
rect 4129 2983 4130 3009
rect 4102 2982 4130 2983
rect 5894 2870 5922 2898
rect 4736 2757 4764 2758
rect 4736 2731 4737 2757
rect 4737 2731 4763 2757
rect 4763 2731 4764 2757
rect 4736 2730 4764 2731
rect 4788 2757 4816 2758
rect 4788 2731 4789 2757
rect 4789 2731 4815 2757
rect 4815 2731 4816 2757
rect 4788 2730 4816 2731
rect 4840 2757 4868 2758
rect 4840 2731 4841 2757
rect 4841 2731 4867 2757
rect 4867 2731 4868 2757
rect 4840 2730 4868 2731
rect 3910 2365 3938 2366
rect 3910 2339 3911 2365
rect 3911 2339 3937 2365
rect 3937 2339 3938 2365
rect 3910 2338 3938 2339
rect 3962 2365 3990 2366
rect 3962 2339 3963 2365
rect 3963 2339 3989 2365
rect 3989 2339 3990 2365
rect 3962 2338 3990 2339
rect 4014 2365 4042 2366
rect 4014 2339 4015 2365
rect 4015 2339 4041 2365
rect 4041 2339 4042 2365
rect 4014 2338 4042 2339
rect 5562 2365 5590 2366
rect 5562 2339 5563 2365
rect 5563 2339 5589 2365
rect 5589 2339 5590 2365
rect 5562 2338 5590 2339
rect 5614 2365 5642 2366
rect 5614 2339 5615 2365
rect 5615 2339 5641 2365
rect 5641 2339 5642 2365
rect 5614 2338 5642 2339
rect 5666 2365 5694 2366
rect 5666 2339 5667 2365
rect 5667 2339 5693 2365
rect 5693 2339 5694 2365
rect 5666 2338 5694 2339
rect 2758 2086 2786 2114
rect 3318 2086 3346 2114
rect 3598 2169 3626 2170
rect 3598 2143 3599 2169
rect 3599 2143 3625 2169
rect 3625 2143 3626 2169
rect 3598 2142 3626 2143
rect 3084 1973 3112 1974
rect 3084 1947 3085 1973
rect 3085 1947 3111 1973
rect 3111 1947 3112 1973
rect 3084 1946 3112 1947
rect 3136 1973 3164 1974
rect 3136 1947 3137 1973
rect 3137 1947 3163 1973
rect 3163 1947 3164 1973
rect 3136 1946 3164 1947
rect 3188 1973 3216 1974
rect 3188 1947 3189 1973
rect 3189 1947 3215 1973
rect 3215 1947 3216 1973
rect 3188 1946 3216 1947
rect 3766 2169 3794 2170
rect 3766 2143 3767 2169
rect 3767 2143 3793 2169
rect 3793 2143 3794 2169
rect 3766 2142 3794 2143
rect 3934 2086 3962 2114
rect 4102 2142 4130 2170
rect 2534 1750 2562 1778
rect 2926 1721 2954 1722
rect 2926 1695 2927 1721
rect 2927 1695 2953 1721
rect 2953 1695 2954 1721
rect 2926 1694 2954 1695
rect 3878 1721 3906 1722
rect 3878 1695 3879 1721
rect 3879 1695 3905 1721
rect 3905 1695 3906 1721
rect 3878 1694 3906 1695
rect 2258 1581 2286 1582
rect 2258 1555 2259 1581
rect 2259 1555 2285 1581
rect 2285 1555 2286 1581
rect 2258 1554 2286 1555
rect 2310 1581 2338 1582
rect 2310 1555 2311 1581
rect 2311 1555 2337 1581
rect 2337 1555 2338 1581
rect 2310 1554 2338 1555
rect 2362 1581 2390 1582
rect 2362 1555 2363 1581
rect 2363 1555 2389 1581
rect 2389 1555 2390 1581
rect 2362 1554 2390 1555
rect 5446 2086 5474 2114
rect 4736 1973 4764 1974
rect 4736 1947 4737 1973
rect 4737 1947 4763 1973
rect 4763 1947 4764 1973
rect 4736 1946 4764 1947
rect 4788 1973 4816 1974
rect 4788 1947 4789 1973
rect 4789 1947 4815 1973
rect 4815 1947 4816 1973
rect 4788 1946 4816 1947
rect 4840 1973 4868 1974
rect 4840 1947 4841 1973
rect 4841 1947 4867 1973
rect 4867 1947 4868 1973
rect 4840 1946 4868 1947
rect 4270 1721 4298 1722
rect 4270 1695 4271 1721
rect 4271 1695 4297 1721
rect 4297 1695 4298 1721
rect 4270 1694 4298 1695
rect 3910 1581 3938 1582
rect 3910 1555 3911 1581
rect 3911 1555 3937 1581
rect 3937 1555 3938 1581
rect 3910 1554 3938 1555
rect 3962 1581 3990 1582
rect 3962 1555 3963 1581
rect 3963 1555 3989 1581
rect 3989 1555 3990 1581
rect 3962 1554 3990 1555
rect 4014 1581 4042 1582
rect 4014 1555 4015 1581
rect 4015 1555 4041 1581
rect 4041 1555 4042 1581
rect 4014 1554 4042 1555
rect 6388 2757 6416 2758
rect 6388 2731 6389 2757
rect 6389 2731 6415 2757
rect 6415 2731 6416 2757
rect 6388 2730 6416 2731
rect 6440 2757 6468 2758
rect 6440 2731 6441 2757
rect 6441 2731 6467 2757
rect 6467 2731 6468 2757
rect 6440 2730 6468 2731
rect 6492 2757 6520 2758
rect 6492 2731 6493 2757
rect 6493 2731 6519 2757
rect 6519 2731 6520 2757
rect 6492 2730 6520 2731
rect 7214 2365 7242 2366
rect 7214 2339 7215 2365
rect 7215 2339 7241 2365
rect 7241 2339 7242 2365
rect 7214 2338 7242 2339
rect 7266 2365 7294 2366
rect 7266 2339 7267 2365
rect 7267 2339 7293 2365
rect 7293 2339 7294 2365
rect 7266 2338 7294 2339
rect 7318 2365 7346 2366
rect 7318 2339 7319 2365
rect 7319 2339 7345 2365
rect 7345 2339 7346 2365
rect 7318 2338 7346 2339
rect 6388 1973 6416 1974
rect 6388 1947 6389 1973
rect 6389 1947 6415 1973
rect 6415 1947 6416 1973
rect 6388 1946 6416 1947
rect 6440 1973 6468 1974
rect 6440 1947 6441 1973
rect 6441 1947 6467 1973
rect 6467 1947 6468 1973
rect 6440 1946 6468 1947
rect 6492 1973 6520 1974
rect 6492 1947 6493 1973
rect 6493 1947 6519 1973
rect 6519 1947 6520 1973
rect 6492 1946 6520 1947
rect 6062 1721 6090 1722
rect 6062 1695 6063 1721
rect 6063 1695 6089 1721
rect 6089 1695 6090 1721
rect 6062 1694 6090 1695
rect 6342 1721 6370 1722
rect 6342 1695 6343 1721
rect 6343 1695 6369 1721
rect 6369 1695 6370 1721
rect 6342 1694 6370 1695
rect 7126 1694 7154 1722
rect 5562 1581 5590 1582
rect 5562 1555 5563 1581
rect 5563 1555 5589 1581
rect 5589 1555 5590 1581
rect 5562 1554 5590 1555
rect 5614 1581 5642 1582
rect 5614 1555 5615 1581
rect 5615 1555 5641 1581
rect 5641 1555 5642 1581
rect 5614 1554 5642 1555
rect 5666 1581 5694 1582
rect 5666 1555 5667 1581
rect 5667 1555 5693 1581
rect 5693 1555 5694 1581
rect 5666 1554 5694 1555
rect 7214 1581 7242 1582
rect 7214 1555 7215 1581
rect 7215 1555 7241 1581
rect 7241 1555 7242 1581
rect 7214 1554 7242 1555
rect 7266 1581 7294 1582
rect 7266 1555 7267 1581
rect 7267 1555 7293 1581
rect 7293 1555 7294 1581
rect 7266 1554 7294 1555
rect 7318 1581 7346 1582
rect 7318 1555 7319 1581
rect 7319 1555 7345 1581
rect 7345 1555 7346 1581
rect 7318 1554 7346 1555
<< metal3 >>
rect 2253 6258 2258 6286
rect 2286 6258 2310 6286
rect 2338 6258 2362 6286
rect 2390 6258 2395 6286
rect 3905 6258 3910 6286
rect 3938 6258 3962 6286
rect 3990 6258 4014 6286
rect 4042 6258 4047 6286
rect 5557 6258 5562 6286
rect 5590 6258 5614 6286
rect 5642 6258 5666 6286
rect 5694 6258 5699 6286
rect 7209 6258 7214 6286
rect 7242 6258 7266 6286
rect 7294 6258 7318 6286
rect 7346 6258 7351 6286
rect 2977 6006 2982 6034
rect 3010 6006 3430 6034
rect 3458 6006 3463 6034
rect 4937 6006 4942 6034
rect 4970 6006 5390 6034
rect 5418 6006 5423 6034
rect 0 5978 400 5992
rect 0 5950 966 5978
rect 994 5950 999 5978
rect 0 5936 400 5950
rect 1427 5866 1432 5894
rect 1460 5866 1484 5894
rect 1512 5866 1536 5894
rect 1564 5866 1569 5894
rect 3079 5866 3084 5894
rect 3112 5866 3136 5894
rect 3164 5866 3188 5894
rect 3216 5866 3221 5894
rect 4731 5866 4736 5894
rect 4764 5866 4788 5894
rect 4816 5866 4840 5894
rect 4868 5866 4873 5894
rect 6383 5866 6388 5894
rect 6416 5866 6440 5894
rect 6468 5866 6492 5894
rect 6520 5866 6525 5894
rect 6001 5726 6006 5754
rect 6034 5726 6902 5754
rect 6930 5726 6935 5754
rect 2253 5474 2258 5502
rect 2286 5474 2310 5502
rect 2338 5474 2362 5502
rect 2390 5474 2395 5502
rect 3905 5474 3910 5502
rect 3938 5474 3962 5502
rect 3990 5474 4014 5502
rect 4042 5474 4047 5502
rect 5557 5474 5562 5502
rect 5590 5474 5614 5502
rect 5642 5474 5666 5502
rect 5694 5474 5699 5502
rect 7209 5474 7214 5502
rect 7242 5474 7266 5502
rect 7294 5474 7318 5502
rect 7346 5474 7351 5502
rect 1427 5082 1432 5110
rect 1460 5082 1484 5110
rect 1512 5082 1536 5110
rect 1564 5082 1569 5110
rect 3079 5082 3084 5110
rect 3112 5082 3136 5110
rect 3164 5082 3188 5110
rect 3216 5082 3221 5110
rect 4731 5082 4736 5110
rect 4764 5082 4788 5110
rect 4816 5082 4840 5110
rect 4868 5082 4873 5110
rect 6383 5082 6388 5110
rect 6416 5082 6440 5110
rect 6468 5082 6492 5110
rect 6520 5082 6525 5110
rect 1633 4886 1638 4914
rect 1666 4886 2422 4914
rect 2450 4886 2455 4914
rect 2253 4690 2258 4718
rect 2286 4690 2310 4718
rect 2338 4690 2362 4718
rect 2390 4690 2395 4718
rect 3905 4690 3910 4718
rect 3938 4690 3962 4718
rect 3990 4690 4014 4718
rect 4042 4690 4047 4718
rect 5557 4690 5562 4718
rect 5590 4690 5614 4718
rect 5642 4690 5666 4718
rect 5694 4690 5699 4718
rect 7209 4690 7214 4718
rect 7242 4690 7266 4718
rect 7294 4690 7318 4718
rect 7346 4690 7351 4718
rect 1427 4298 1432 4326
rect 1460 4298 1484 4326
rect 1512 4298 1536 4326
rect 1564 4298 1569 4326
rect 3079 4298 3084 4326
rect 3112 4298 3136 4326
rect 3164 4298 3188 4326
rect 3216 4298 3221 4326
rect 4731 4298 4736 4326
rect 4764 4298 4788 4326
rect 4816 4298 4840 4326
rect 4868 4298 4873 4326
rect 6383 4298 6388 4326
rect 6416 4298 6440 4326
rect 6468 4298 6492 4326
rect 6520 4298 6525 4326
rect 3481 3990 3486 4018
rect 3514 3990 5054 4018
rect 5082 3990 5087 4018
rect 2253 3906 2258 3934
rect 2286 3906 2310 3934
rect 2338 3906 2362 3934
rect 2390 3906 2395 3934
rect 3905 3906 3910 3934
rect 3938 3906 3962 3934
rect 3990 3906 4014 3934
rect 4042 3906 4047 3934
rect 5557 3906 5562 3934
rect 5590 3906 5614 3934
rect 5642 3906 5666 3934
rect 5694 3906 5699 3934
rect 7209 3906 7214 3934
rect 7242 3906 7266 3934
rect 7294 3906 7318 3934
rect 7346 3906 7351 3934
rect 3985 3822 3990 3850
rect 4018 3822 5446 3850
rect 5474 3822 5479 3850
rect 2529 3710 2534 3738
rect 2562 3710 3598 3738
rect 3626 3710 4158 3738
rect 4186 3710 4191 3738
rect 2473 3654 2478 3682
rect 2506 3654 3486 3682
rect 3514 3654 3519 3682
rect 3486 3570 3514 3654
rect 3822 3626 3850 3710
rect 3817 3598 3822 3626
rect 3850 3598 3855 3626
rect 3486 3542 4046 3570
rect 4074 3542 4079 3570
rect 1427 3514 1432 3542
rect 1460 3514 1484 3542
rect 1512 3514 1536 3542
rect 1564 3514 1569 3542
rect 3079 3514 3084 3542
rect 3112 3514 3136 3542
rect 3164 3514 3188 3542
rect 3216 3514 3221 3542
rect 4731 3514 4736 3542
rect 4764 3514 4788 3542
rect 4816 3514 4840 3542
rect 4868 3514 4873 3542
rect 6383 3514 6388 3542
rect 6416 3514 6440 3542
rect 6468 3514 6492 3542
rect 6520 3514 6525 3542
rect 2865 3318 2870 3346
rect 2898 3318 3486 3346
rect 3514 3318 3519 3346
rect 2361 3206 2366 3234
rect 2394 3206 3094 3234
rect 3122 3206 3127 3234
rect 2253 3122 2258 3150
rect 2286 3122 2310 3150
rect 2338 3122 2362 3150
rect 2390 3122 2395 3150
rect 2478 3066 2506 3206
rect 3905 3122 3910 3150
rect 3938 3122 3962 3150
rect 3990 3122 4014 3150
rect 4042 3122 4047 3150
rect 5557 3122 5562 3150
rect 5590 3122 5614 3150
rect 5642 3122 5666 3150
rect 5694 3122 5699 3150
rect 7209 3122 7214 3150
rect 7242 3122 7266 3150
rect 7294 3122 7318 3150
rect 7346 3122 7351 3150
rect 2249 3038 2254 3066
rect 2282 3038 2506 3066
rect 3481 2982 3486 3010
rect 3514 2982 3878 3010
rect 3906 2982 4102 3010
rect 4130 2982 4135 3010
rect 2137 2926 2142 2954
rect 2170 2926 2590 2954
rect 2618 2926 2814 2954
rect 2842 2926 2847 2954
rect 4102 2898 4130 2982
rect 4102 2870 5894 2898
rect 5922 2870 5927 2898
rect 1427 2730 1432 2758
rect 1460 2730 1484 2758
rect 1512 2730 1536 2758
rect 1564 2730 1569 2758
rect 3079 2730 3084 2758
rect 3112 2730 3136 2758
rect 3164 2730 3188 2758
rect 3216 2730 3221 2758
rect 4731 2730 4736 2758
rect 4764 2730 4788 2758
rect 4816 2730 4840 2758
rect 4868 2730 4873 2758
rect 6383 2730 6388 2758
rect 6416 2730 6440 2758
rect 6468 2730 6492 2758
rect 6520 2730 6525 2758
rect 1521 2534 1526 2562
rect 1554 2534 2086 2562
rect 2114 2534 2119 2562
rect 3262 2534 3374 2562
rect 3402 2534 3407 2562
rect 2529 2478 2534 2506
rect 2562 2478 3038 2506
rect 3066 2478 3071 2506
rect 3262 2394 3290 2534
rect 3257 2366 3262 2394
rect 3290 2366 3295 2394
rect 2253 2338 2258 2366
rect 2286 2338 2310 2366
rect 2338 2338 2362 2366
rect 2390 2338 2395 2366
rect 3905 2338 3910 2366
rect 3938 2338 3962 2366
rect 3990 2338 4014 2366
rect 4042 2338 4047 2366
rect 5557 2338 5562 2366
rect 5590 2338 5614 2366
rect 5642 2338 5666 2366
rect 5694 2338 5699 2366
rect 7209 2338 7214 2366
rect 7242 2338 7266 2366
rect 7294 2338 7318 2366
rect 7346 2338 7351 2366
rect 2473 2254 2478 2282
rect 2506 2254 2702 2282
rect 2730 2254 2735 2282
rect 2641 2198 2646 2226
rect 2674 2198 3206 2226
rect 3234 2198 3794 2226
rect 3766 2170 3794 2198
rect 2081 2142 2086 2170
rect 2114 2142 2982 2170
rect 3010 2142 3598 2170
rect 3626 2142 3631 2170
rect 3761 2142 3766 2170
rect 3794 2142 4102 2170
rect 4130 2142 4135 2170
rect 2753 2086 2758 2114
rect 2786 2086 3318 2114
rect 3346 2086 3934 2114
rect 3962 2086 5446 2114
rect 5474 2086 5479 2114
rect 0 2002 400 2016
rect 0 1974 966 2002
rect 994 1974 999 2002
rect 0 1960 400 1974
rect 1427 1946 1432 1974
rect 1460 1946 1484 1974
rect 1512 1946 1536 1974
rect 1564 1946 1569 1974
rect 3079 1946 3084 1974
rect 3112 1946 3136 1974
rect 3164 1946 3188 1974
rect 3216 1946 3221 1974
rect 4731 1946 4736 1974
rect 4764 1946 4788 1974
rect 4816 1946 4840 1974
rect 4868 1946 4873 1974
rect 6383 1946 6388 1974
rect 6416 1946 6440 1974
rect 6468 1946 6492 1974
rect 6520 1946 6525 1974
rect 1689 1750 1694 1778
rect 1722 1750 2366 1778
rect 2394 1750 2534 1778
rect 2562 1750 2567 1778
rect 2081 1694 2086 1722
rect 2114 1694 2926 1722
rect 2954 1694 2959 1722
rect 3873 1694 3878 1722
rect 3906 1694 4270 1722
rect 4298 1694 4303 1722
rect 6057 1694 6062 1722
rect 6090 1694 6342 1722
rect 6370 1694 7126 1722
rect 7154 1694 7159 1722
rect 2253 1554 2258 1582
rect 2286 1554 2310 1582
rect 2338 1554 2362 1582
rect 2390 1554 2395 1582
rect 3905 1554 3910 1582
rect 3938 1554 3962 1582
rect 3990 1554 4014 1582
rect 4042 1554 4047 1582
rect 5557 1554 5562 1582
rect 5590 1554 5614 1582
rect 5642 1554 5666 1582
rect 5694 1554 5699 1582
rect 7209 1554 7214 1582
rect 7242 1554 7266 1582
rect 7294 1554 7318 1582
rect 7346 1554 7351 1582
<< via3 >>
rect 2258 6258 2286 6286
rect 2310 6258 2338 6286
rect 2362 6258 2390 6286
rect 3910 6258 3938 6286
rect 3962 6258 3990 6286
rect 4014 6258 4042 6286
rect 5562 6258 5590 6286
rect 5614 6258 5642 6286
rect 5666 6258 5694 6286
rect 7214 6258 7242 6286
rect 7266 6258 7294 6286
rect 7318 6258 7346 6286
rect 1432 5866 1460 5894
rect 1484 5866 1512 5894
rect 1536 5866 1564 5894
rect 3084 5866 3112 5894
rect 3136 5866 3164 5894
rect 3188 5866 3216 5894
rect 4736 5866 4764 5894
rect 4788 5866 4816 5894
rect 4840 5866 4868 5894
rect 6388 5866 6416 5894
rect 6440 5866 6468 5894
rect 6492 5866 6520 5894
rect 2258 5474 2286 5502
rect 2310 5474 2338 5502
rect 2362 5474 2390 5502
rect 3910 5474 3938 5502
rect 3962 5474 3990 5502
rect 4014 5474 4042 5502
rect 5562 5474 5590 5502
rect 5614 5474 5642 5502
rect 5666 5474 5694 5502
rect 7214 5474 7242 5502
rect 7266 5474 7294 5502
rect 7318 5474 7346 5502
rect 1432 5082 1460 5110
rect 1484 5082 1512 5110
rect 1536 5082 1564 5110
rect 3084 5082 3112 5110
rect 3136 5082 3164 5110
rect 3188 5082 3216 5110
rect 4736 5082 4764 5110
rect 4788 5082 4816 5110
rect 4840 5082 4868 5110
rect 6388 5082 6416 5110
rect 6440 5082 6468 5110
rect 6492 5082 6520 5110
rect 2258 4690 2286 4718
rect 2310 4690 2338 4718
rect 2362 4690 2390 4718
rect 3910 4690 3938 4718
rect 3962 4690 3990 4718
rect 4014 4690 4042 4718
rect 5562 4690 5590 4718
rect 5614 4690 5642 4718
rect 5666 4690 5694 4718
rect 7214 4690 7242 4718
rect 7266 4690 7294 4718
rect 7318 4690 7346 4718
rect 1432 4298 1460 4326
rect 1484 4298 1512 4326
rect 1536 4298 1564 4326
rect 3084 4298 3112 4326
rect 3136 4298 3164 4326
rect 3188 4298 3216 4326
rect 4736 4298 4764 4326
rect 4788 4298 4816 4326
rect 4840 4298 4868 4326
rect 6388 4298 6416 4326
rect 6440 4298 6468 4326
rect 6492 4298 6520 4326
rect 2258 3906 2286 3934
rect 2310 3906 2338 3934
rect 2362 3906 2390 3934
rect 3910 3906 3938 3934
rect 3962 3906 3990 3934
rect 4014 3906 4042 3934
rect 5562 3906 5590 3934
rect 5614 3906 5642 3934
rect 5666 3906 5694 3934
rect 7214 3906 7242 3934
rect 7266 3906 7294 3934
rect 7318 3906 7346 3934
rect 1432 3514 1460 3542
rect 1484 3514 1512 3542
rect 1536 3514 1564 3542
rect 3084 3514 3112 3542
rect 3136 3514 3164 3542
rect 3188 3514 3216 3542
rect 4736 3514 4764 3542
rect 4788 3514 4816 3542
rect 4840 3514 4868 3542
rect 6388 3514 6416 3542
rect 6440 3514 6468 3542
rect 6492 3514 6520 3542
rect 2258 3122 2286 3150
rect 2310 3122 2338 3150
rect 2362 3122 2390 3150
rect 3910 3122 3938 3150
rect 3962 3122 3990 3150
rect 4014 3122 4042 3150
rect 5562 3122 5590 3150
rect 5614 3122 5642 3150
rect 5666 3122 5694 3150
rect 7214 3122 7242 3150
rect 7266 3122 7294 3150
rect 7318 3122 7346 3150
rect 1432 2730 1460 2758
rect 1484 2730 1512 2758
rect 1536 2730 1564 2758
rect 3084 2730 3112 2758
rect 3136 2730 3164 2758
rect 3188 2730 3216 2758
rect 4736 2730 4764 2758
rect 4788 2730 4816 2758
rect 4840 2730 4868 2758
rect 6388 2730 6416 2758
rect 6440 2730 6468 2758
rect 6492 2730 6520 2758
rect 2258 2338 2286 2366
rect 2310 2338 2338 2366
rect 2362 2338 2390 2366
rect 3910 2338 3938 2366
rect 3962 2338 3990 2366
rect 4014 2338 4042 2366
rect 5562 2338 5590 2366
rect 5614 2338 5642 2366
rect 5666 2338 5694 2366
rect 7214 2338 7242 2366
rect 7266 2338 7294 2366
rect 7318 2338 7346 2366
rect 1432 1946 1460 1974
rect 1484 1946 1512 1974
rect 1536 1946 1564 1974
rect 3084 1946 3112 1974
rect 3136 1946 3164 1974
rect 3188 1946 3216 1974
rect 4736 1946 4764 1974
rect 4788 1946 4816 1974
rect 4840 1946 4868 1974
rect 6388 1946 6416 1974
rect 6440 1946 6468 1974
rect 6492 1946 6520 1974
rect 2258 1554 2286 1582
rect 2310 1554 2338 1582
rect 2362 1554 2390 1582
rect 3910 1554 3938 1582
rect 3962 1554 3990 1582
rect 4014 1554 4042 1582
rect 5562 1554 5590 1582
rect 5614 1554 5642 1582
rect 5666 1554 5694 1582
rect 7214 1554 7242 1582
rect 7266 1554 7294 1582
rect 7318 1554 7346 1582
<< metal4 >>
rect 1418 5894 1578 6302
rect 1418 5866 1432 5894
rect 1460 5866 1484 5894
rect 1512 5866 1536 5894
rect 1564 5866 1578 5894
rect 1418 5110 1578 5866
rect 1418 5082 1432 5110
rect 1460 5082 1484 5110
rect 1512 5082 1536 5110
rect 1564 5082 1578 5110
rect 1418 4326 1578 5082
rect 1418 4298 1432 4326
rect 1460 4298 1484 4326
rect 1512 4298 1536 4326
rect 1564 4298 1578 4326
rect 1418 3542 1578 4298
rect 1418 3514 1432 3542
rect 1460 3514 1484 3542
rect 1512 3514 1536 3542
rect 1564 3514 1578 3542
rect 1418 2758 1578 3514
rect 1418 2730 1432 2758
rect 1460 2730 1484 2758
rect 1512 2730 1536 2758
rect 1564 2730 1578 2758
rect 1418 1974 1578 2730
rect 1418 1946 1432 1974
rect 1460 1946 1484 1974
rect 1512 1946 1536 1974
rect 1564 1946 1578 1974
rect 1418 1538 1578 1946
rect 2244 6286 2404 6302
rect 2244 6258 2258 6286
rect 2286 6258 2310 6286
rect 2338 6258 2362 6286
rect 2390 6258 2404 6286
rect 2244 5502 2404 6258
rect 2244 5474 2258 5502
rect 2286 5474 2310 5502
rect 2338 5474 2362 5502
rect 2390 5474 2404 5502
rect 2244 4718 2404 5474
rect 2244 4690 2258 4718
rect 2286 4690 2310 4718
rect 2338 4690 2362 4718
rect 2390 4690 2404 4718
rect 2244 3934 2404 4690
rect 2244 3906 2258 3934
rect 2286 3906 2310 3934
rect 2338 3906 2362 3934
rect 2390 3906 2404 3934
rect 2244 3150 2404 3906
rect 2244 3122 2258 3150
rect 2286 3122 2310 3150
rect 2338 3122 2362 3150
rect 2390 3122 2404 3150
rect 2244 2366 2404 3122
rect 2244 2338 2258 2366
rect 2286 2338 2310 2366
rect 2338 2338 2362 2366
rect 2390 2338 2404 2366
rect 2244 1582 2404 2338
rect 2244 1554 2258 1582
rect 2286 1554 2310 1582
rect 2338 1554 2362 1582
rect 2390 1554 2404 1582
rect 2244 1538 2404 1554
rect 3070 5894 3230 6302
rect 3070 5866 3084 5894
rect 3112 5866 3136 5894
rect 3164 5866 3188 5894
rect 3216 5866 3230 5894
rect 3070 5110 3230 5866
rect 3070 5082 3084 5110
rect 3112 5082 3136 5110
rect 3164 5082 3188 5110
rect 3216 5082 3230 5110
rect 3070 4326 3230 5082
rect 3070 4298 3084 4326
rect 3112 4298 3136 4326
rect 3164 4298 3188 4326
rect 3216 4298 3230 4326
rect 3070 3542 3230 4298
rect 3070 3514 3084 3542
rect 3112 3514 3136 3542
rect 3164 3514 3188 3542
rect 3216 3514 3230 3542
rect 3070 2758 3230 3514
rect 3070 2730 3084 2758
rect 3112 2730 3136 2758
rect 3164 2730 3188 2758
rect 3216 2730 3230 2758
rect 3070 1974 3230 2730
rect 3070 1946 3084 1974
rect 3112 1946 3136 1974
rect 3164 1946 3188 1974
rect 3216 1946 3230 1974
rect 3070 1538 3230 1946
rect 3896 6286 4056 6302
rect 3896 6258 3910 6286
rect 3938 6258 3962 6286
rect 3990 6258 4014 6286
rect 4042 6258 4056 6286
rect 3896 5502 4056 6258
rect 3896 5474 3910 5502
rect 3938 5474 3962 5502
rect 3990 5474 4014 5502
rect 4042 5474 4056 5502
rect 3896 4718 4056 5474
rect 3896 4690 3910 4718
rect 3938 4690 3962 4718
rect 3990 4690 4014 4718
rect 4042 4690 4056 4718
rect 3896 3934 4056 4690
rect 3896 3906 3910 3934
rect 3938 3906 3962 3934
rect 3990 3906 4014 3934
rect 4042 3906 4056 3934
rect 3896 3150 4056 3906
rect 3896 3122 3910 3150
rect 3938 3122 3962 3150
rect 3990 3122 4014 3150
rect 4042 3122 4056 3150
rect 3896 2366 4056 3122
rect 3896 2338 3910 2366
rect 3938 2338 3962 2366
rect 3990 2338 4014 2366
rect 4042 2338 4056 2366
rect 3896 1582 4056 2338
rect 3896 1554 3910 1582
rect 3938 1554 3962 1582
rect 3990 1554 4014 1582
rect 4042 1554 4056 1582
rect 3896 1538 4056 1554
rect 4722 5894 4882 6302
rect 4722 5866 4736 5894
rect 4764 5866 4788 5894
rect 4816 5866 4840 5894
rect 4868 5866 4882 5894
rect 4722 5110 4882 5866
rect 4722 5082 4736 5110
rect 4764 5082 4788 5110
rect 4816 5082 4840 5110
rect 4868 5082 4882 5110
rect 4722 4326 4882 5082
rect 4722 4298 4736 4326
rect 4764 4298 4788 4326
rect 4816 4298 4840 4326
rect 4868 4298 4882 4326
rect 4722 3542 4882 4298
rect 4722 3514 4736 3542
rect 4764 3514 4788 3542
rect 4816 3514 4840 3542
rect 4868 3514 4882 3542
rect 4722 2758 4882 3514
rect 4722 2730 4736 2758
rect 4764 2730 4788 2758
rect 4816 2730 4840 2758
rect 4868 2730 4882 2758
rect 4722 1974 4882 2730
rect 4722 1946 4736 1974
rect 4764 1946 4788 1974
rect 4816 1946 4840 1974
rect 4868 1946 4882 1974
rect 4722 1538 4882 1946
rect 5548 6286 5708 6302
rect 5548 6258 5562 6286
rect 5590 6258 5614 6286
rect 5642 6258 5666 6286
rect 5694 6258 5708 6286
rect 5548 5502 5708 6258
rect 5548 5474 5562 5502
rect 5590 5474 5614 5502
rect 5642 5474 5666 5502
rect 5694 5474 5708 5502
rect 5548 4718 5708 5474
rect 5548 4690 5562 4718
rect 5590 4690 5614 4718
rect 5642 4690 5666 4718
rect 5694 4690 5708 4718
rect 5548 3934 5708 4690
rect 5548 3906 5562 3934
rect 5590 3906 5614 3934
rect 5642 3906 5666 3934
rect 5694 3906 5708 3934
rect 5548 3150 5708 3906
rect 5548 3122 5562 3150
rect 5590 3122 5614 3150
rect 5642 3122 5666 3150
rect 5694 3122 5708 3150
rect 5548 2366 5708 3122
rect 5548 2338 5562 2366
rect 5590 2338 5614 2366
rect 5642 2338 5666 2366
rect 5694 2338 5708 2366
rect 5548 1582 5708 2338
rect 5548 1554 5562 1582
rect 5590 1554 5614 1582
rect 5642 1554 5666 1582
rect 5694 1554 5708 1582
rect 5548 1538 5708 1554
rect 6374 5894 6534 6302
rect 6374 5866 6388 5894
rect 6416 5866 6440 5894
rect 6468 5866 6492 5894
rect 6520 5866 6534 5894
rect 6374 5110 6534 5866
rect 6374 5082 6388 5110
rect 6416 5082 6440 5110
rect 6468 5082 6492 5110
rect 6520 5082 6534 5110
rect 6374 4326 6534 5082
rect 6374 4298 6388 4326
rect 6416 4298 6440 4326
rect 6468 4298 6492 4326
rect 6520 4298 6534 4326
rect 6374 3542 6534 4298
rect 6374 3514 6388 3542
rect 6416 3514 6440 3542
rect 6468 3514 6492 3542
rect 6520 3514 6534 3542
rect 6374 2758 6534 3514
rect 6374 2730 6388 2758
rect 6416 2730 6440 2758
rect 6468 2730 6492 2758
rect 6520 2730 6534 2758
rect 6374 1974 6534 2730
rect 6374 1946 6388 1974
rect 6416 1946 6440 1974
rect 6468 1946 6492 1974
rect 6520 1946 6534 1974
rect 6374 1538 6534 1946
rect 7200 6286 7360 6302
rect 7200 6258 7214 6286
rect 7242 6258 7266 6286
rect 7294 6258 7318 6286
rect 7346 6258 7360 6286
rect 7200 5502 7360 6258
rect 7200 5474 7214 5502
rect 7242 5474 7266 5502
rect 7294 5474 7318 5502
rect 7346 5474 7360 5502
rect 7200 4718 7360 5474
rect 7200 4690 7214 4718
rect 7242 4690 7266 4718
rect 7294 4690 7318 4718
rect 7346 4690 7360 4718
rect 7200 3934 7360 4690
rect 7200 3906 7214 3934
rect 7242 3906 7266 3934
rect 7294 3906 7318 3934
rect 7346 3906 7360 3934
rect 7200 3150 7360 3906
rect 7200 3122 7214 3150
rect 7242 3122 7266 3150
rect 7294 3122 7318 3150
rect 7346 3122 7360 3150
rect 7200 2366 7360 3122
rect 7200 2338 7214 2366
rect 7242 2338 7266 2366
rect 7294 2338 7318 2366
rect 7346 2338 7360 2366
rect 7200 1582 7360 2338
rect 7200 1554 7214 1582
rect 7242 1554 7266 1582
rect 7294 1554 7318 1582
rect 7346 1554 7360 1582
rect 7200 1538 7360 1554
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__09__A1 Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 2800 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__10__I
timestamp 1669390400
transform 1 0 4088 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__17__A1
timestamp 1669390400
transform 1 0 2576 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__19__B
timestamp 1669390400
transform -1 0 3528 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1669390400
transform -1 0 2128 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1669390400
transform -1 0 952 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1669390400
transform 1 0 5712 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1669390400
transform -1 0 3920 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1669390400
transform -1 0 6384 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2 Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 784 0 1 1568
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20 Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 1792 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26
timestamp 1669390400
transform 1 0 2128 0 1 1568
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34 Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 2576 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37
timestamp 1669390400
transform 1 0 2744 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54
timestamp 1669390400
transform 1 0 3696 0 1 1568
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58
timestamp 1669390400
transform 1 0 3920 0 1 1568
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66
timestamp 1669390400
transform 1 0 4368 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_72 Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 4704 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80
timestamp 1669390400
transform 1 0 5152 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90
timestamp 1669390400
transform 1 0 5712 0 1 1568
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_98
timestamp 1669390400
transform 1 0 6160 0 1 1568
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_102
timestamp 1669390400
transform 1 0 6384 0 1 1568
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_104
timestamp 1669390400
transform 1 0 6496 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_107
timestamp 1669390400
transform 1 0 6664 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_115
timestamp 1669390400
transform 1 0 7112 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_2
timestamp 1669390400
transform 1 0 784 0 -1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_17
timestamp 1669390400
transform 1 0 1624 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_21
timestamp 1669390400
transform 1 0 1848 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_29
timestamp 1669390400
transform 1 0 2296 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_39
timestamp 1669390400
transform 1 0 2856 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_49
timestamp 1669390400
transform 1 0 3416 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_59
timestamp 1669390400
transform 1 0 3976 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_67
timestamp 1669390400
transform 1 0 4424 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_73 Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 4760 0 -1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_89
timestamp 1669390400
transform 1 0 5656 0 -1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_92
timestamp 1669390400
transform 1 0 5824 0 -1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_108
timestamp 1669390400
transform 1 0 6720 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_2
timestamp 1669390400
transform 1 0 784 0 1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_5
timestamp 1669390400
transform 1 0 952 0 1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_21
timestamp 1669390400
transform 1 0 1848 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_32
timestamp 1669390400
transform 1 0 2464 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_34
timestamp 1669390400
transform 1 0 2576 0 1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_37
timestamp 1669390400
transform 1 0 2744 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_49 Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 3416 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_81
timestamp 1669390400
transform 1 0 5208 0 1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_97
timestamp 1669390400
transform 1 0 6104 0 1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_105
timestamp 1669390400
transform 1 0 6552 0 1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_108
timestamp 1669390400
transform 1 0 6720 0 1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_2
timestamp 1669390400
transform 1 0 784 0 -1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_36
timestamp 1669390400
transform 1 0 2688 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_40
timestamp 1669390400
transform 1 0 2912 0 -1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_48
timestamp 1669390400
transform 1 0 3360 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_52
timestamp 1669390400
transform 1 0 3584 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_54
timestamp 1669390400
transform 1 0 3696 0 -1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_59
timestamp 1669390400
transform 1 0 3976 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_63
timestamp 1669390400
transform 1 0 4200 0 -1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_73
timestamp 1669390400
transform 1 0 4760 0 -1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_105
timestamp 1669390400
transform 1 0 6552 0 -1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_113
timestamp 1669390400
transform 1 0 7000 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_115
timestamp 1669390400
transform 1 0 7112 0 -1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_2
timestamp 1669390400
transform 1 0 784 0 1 3136
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_18
timestamp 1669390400
transform 1 0 1680 0 1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_26
timestamp 1669390400
transform 1 0 2128 0 1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_34
timestamp 1669390400
transform 1 0 2576 0 1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_37
timestamp 1669390400
transform 1 0 2744 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_47
timestamp 1669390400
transform 1 0 3304 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_51
timestamp 1669390400
transform 1 0 3528 0 1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_83
timestamp 1669390400
transform 1 0 5320 0 1 3136
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_99
timestamp 1669390400
transform 1 0 6216 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_103
timestamp 1669390400
transform 1 0 6440 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_105
timestamp 1669390400
transform 1 0 6552 0 1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_108
timestamp 1669390400
transform 1 0 6720 0 1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_2
timestamp 1669390400
transform 1 0 784 0 -1 3920
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_18
timestamp 1669390400
transform 1 0 1680 0 -1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_26
timestamp 1669390400
transform 1 0 2128 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_36
timestamp 1669390400
transform 1 0 2688 0 -1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_44
timestamp 1669390400
transform 1 0 3136 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_46
timestamp 1669390400
transform 1 0 3248 0 -1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_55
timestamp 1669390400
transform 1 0 3752 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_65
timestamp 1669390400
transform 1 0 4312 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_69
timestamp 1669390400
transform 1 0 4536 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_73
timestamp 1669390400
transform 1 0 4760 0 -1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_105
timestamp 1669390400
transform 1 0 6552 0 -1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_113
timestamp 1669390400
transform 1 0 7000 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_115
timestamp 1669390400
transform 1 0 7112 0 -1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_2
timestamp 1669390400
transform 1 0 784 0 1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_34
timestamp 1669390400
transform 1 0 2576 0 1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_37 Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 2744 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_101
timestamp 1669390400
transform 1 0 6328 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_105
timestamp 1669390400
transform 1 0 6552 0 1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_108
timestamp 1669390400
transform 1 0 6720 0 1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_2
timestamp 1669390400
transform 1 0 784 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_66
timestamp 1669390400
transform 1 0 4368 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_70
timestamp 1669390400
transform 1 0 4592 0 -1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_73
timestamp 1669390400
transform 1 0 4760 0 -1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_105
timestamp 1669390400
transform 1 0 6552 0 -1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_113
timestamp 1669390400
transform 1 0 7000 0 -1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_115
timestamp 1669390400
transform 1 0 7112 0 -1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_2
timestamp 1669390400
transform 1 0 784 0 1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_34
timestamp 1669390400
transform 1 0 2576 0 1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_37
timestamp 1669390400
transform 1 0 2744 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_101
timestamp 1669390400
transform 1 0 6328 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_105
timestamp 1669390400
transform 1 0 6552 0 1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_108
timestamp 1669390400
transform 1 0 6720 0 1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_2
timestamp 1669390400
transform 1 0 784 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_66
timestamp 1669390400
transform 1 0 4368 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_70
timestamp 1669390400
transform 1 0 4592 0 -1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_9_73
timestamp 1669390400
transform 1 0 4760 0 -1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_105
timestamp 1669390400
transform 1 0 6552 0 -1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_113
timestamp 1669390400
transform 1 0 7000 0 -1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_115
timestamp 1669390400
transform 1 0 7112 0 -1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_2
timestamp 1669390400
transform 1 0 784 0 1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_17
timestamp 1669390400
transform 1 0 1624 0 1 5488
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_33
timestamp 1669390400
transform 1 0 2520 0 1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_37
timestamp 1669390400
transform 1 0 2744 0 1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_69
timestamp 1669390400
transform 1 0 4536 0 1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_77
timestamp 1669390400
transform 1 0 4984 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_81
timestamp 1669390400
transform 1 0 5208 0 1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_83
timestamp 1669390400
transform 1 0 5320 0 1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_98
timestamp 1669390400
transform 1 0 6160 0 1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_108
timestamp 1669390400
transform 1 0 6720 0 1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_2
timestamp 1669390400
transform 1 0 784 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_6
timestamp 1669390400
transform 1 0 1008 0 -1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_21
timestamp 1669390400
transform 1 0 1848 0 -1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_29
timestamp 1669390400
transform 1 0 2296 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_33
timestamp 1669390400
transform 1 0 2520 0 -1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_37
timestamp 1669390400
transform 1 0 2744 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_41
timestamp 1669390400
transform 1 0 2968 0 -1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_56
timestamp 1669390400
transform 1 0 3808 0 -1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_64
timestamp 1669390400
transform 1 0 4256 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_68
timestamp 1669390400
transform 1 0 4480 0 -1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_72
timestamp 1669390400
transform 1 0 4704 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_76
timestamp 1669390400
transform 1 0 4928 0 -1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_91
timestamp 1669390400
transform 1 0 5768 0 -1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_99
timestamp 1669390400
transform 1 0 6216 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_103
timestamp 1669390400
transform 1 0 6440 0 -1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_107
timestamp 1669390400
transform 1 0 6664 0 -1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_115
timestamp 1669390400
transform 1 0 7112 0 -1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_0 Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 672 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_1
timestamp 1669390400
transform -1 0 7280 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_2
timestamp 1669390400
transform 1 0 672 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_3
timestamp 1669390400
transform -1 0 7280 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_4
timestamp 1669390400
transform 1 0 672 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_5
timestamp 1669390400
transform -1 0 7280 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_6
timestamp 1669390400
transform 1 0 672 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_7
timestamp 1669390400
transform -1 0 7280 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_8
timestamp 1669390400
transform 1 0 672 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_9
timestamp 1669390400
transform -1 0 7280 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_10
timestamp 1669390400
transform 1 0 672 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_11
timestamp 1669390400
transform -1 0 7280 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_12
timestamp 1669390400
transform 1 0 672 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_13
timestamp 1669390400
transform -1 0 7280 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_14
timestamp 1669390400
transform 1 0 672 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_15
timestamp 1669390400
transform -1 0 7280 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_16
timestamp 1669390400
transform 1 0 672 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_17
timestamp 1669390400
transform -1 0 7280 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_18
timestamp 1669390400
transform 1 0 672 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_19
timestamp 1669390400
transform -1 0 7280 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_20
timestamp 1669390400
transform 1 0 672 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_21
timestamp 1669390400
transform -1 0 7280 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_22
timestamp 1669390400
transform 1 0 672 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_23
timestamp 1669390400
transform -1 0 7280 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_24 Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 2632 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_25
timestamp 1669390400
transform 1 0 4592 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_26
timestamp 1669390400
transform 1 0 6552 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_27
timestamp 1669390400
transform 1 0 4648 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_28
timestamp 1669390400
transform 1 0 2632 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_29
timestamp 1669390400
transform 1 0 6608 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_30
timestamp 1669390400
transform 1 0 4648 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_31
timestamp 1669390400
transform 1 0 2632 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_32
timestamp 1669390400
transform 1 0 6608 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_33
timestamp 1669390400
transform 1 0 4648 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_34
timestamp 1669390400
transform 1 0 2632 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_35
timestamp 1669390400
transform 1 0 6608 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_36
timestamp 1669390400
transform 1 0 4648 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_37
timestamp 1669390400
transform 1 0 2632 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_38
timestamp 1669390400
transform 1 0 6608 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_39
timestamp 1669390400
transform 1 0 4648 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_40
timestamp 1669390400
transform 1 0 2632 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_41
timestamp 1669390400
transform 1 0 6608 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_42
timestamp 1669390400
transform 1 0 2632 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_43
timestamp 1669390400
transform 1 0 4592 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_44
timestamp 1669390400
transform 1 0 6552 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _07_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 1960 0 -1 2352
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _08_
timestamp 1669390400
transform 1 0 2240 0 1 1568
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _09_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 2464 0 1 2352
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _10_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 3976 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _11_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 2240 0 -1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _12_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 3416 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _13_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 3304 0 -1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _14_
timestamp 1669390400
transform -1 0 3976 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _15_
timestamp 1669390400
transform 1 0 3864 0 -1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _16_
timestamp 1669390400
transform -1 0 2856 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _17_
timestamp 1669390400
transform -1 0 2576 0 1 3136
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _18_
timestamp 1669390400
transform -1 0 3416 0 1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _19_
timestamp 1669390400
transform -1 0 3304 0 1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input1 Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 2800 0 1 1568
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input2
timestamp 1669390400
transform 1 0 896 0 1 1568
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input3
timestamp 1669390400
transform -1 0 5712 0 1 1568
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input4
timestamp 1669390400
transform -1 0 4368 0 1 1568
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input5
timestamp 1669390400
transform -1 0 6160 0 1 1568
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output6 Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 1624 0 1 5488
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output7
timestamp 1669390400
transform -1 0 1624 0 -1 2352
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output8
timestamp 1669390400
transform 1 0 5376 0 1 5488
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output9
timestamp 1669390400
transform 1 0 4984 0 -1 6272
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output10
timestamp 1669390400
transform 1 0 3024 0 -1 6272
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output11
timestamp 1669390400
transform -1 0 1848 0 -1 6272
box -43 -43 827 435
<< labels >>
flabel metal2 s 2408 0 2464 400 0 FreeSans 224 90 0 0 INmb
port 0 nsew signal input
flabel metal2 s 840 0 896 400 0 FreeSans 224 90 0 0 INpb
port 1 nsew signal input
flabel metal2 s 5544 0 5600 400 0 FreeSans 224 90 0 0 OUTm
port 2 nsew signal input
flabel metal2 s 3976 0 4032 400 0 FreeSans 224 90 0 0 OUTp
port 3 nsew signal input
flabel metal3 s 0 5936 400 5992 0 FreeSans 224 0 0 0 cmnmos
port 4 nsew signal tristate
flabel metal3 s 0 1960 400 2016 0 FreeSans 224 0 0 0 cmpmos
port 5 nsew signal tristate
flabel metal2 s 7112 0 7168 400 0 FreeSans 224 90 0 0 oe
port 6 nsew signal input
flabel metal2 s 6888 7600 6944 8000 0 FreeSans 224 90 0 0 omnmos
port 7 nsew signal tristate
flabel metal2 s 4928 7600 4984 8000 0 FreeSans 224 90 0 0 ompmos
port 8 nsew signal tristate
flabel metal2 s 2968 7600 3024 8000 0 FreeSans 224 90 0 0 opnmos
port 9 nsew signal tristate
flabel metal2 s 1008 7600 1064 8000 0 FreeSans 224 90 0 0 oppmos
port 10 nsew signal tristate
flabel metal4 s 1418 1538 1578 6302 0 FreeSans 640 90 0 0 vdd
port 11 nsew power bidirectional
flabel metal4 s 3070 1538 3230 6302 0 FreeSans 640 90 0 0 vdd
port 11 nsew power bidirectional
flabel metal4 s 4722 1538 4882 6302 0 FreeSans 640 90 0 0 vdd
port 11 nsew power bidirectional
flabel metal4 s 6374 1538 6534 6302 0 FreeSans 640 90 0 0 vdd
port 11 nsew power bidirectional
flabel metal4 s 2244 1538 2404 6302 0 FreeSans 640 90 0 0 vss
port 12 nsew ground bidirectional
flabel metal4 s 3896 1538 4056 6302 0 FreeSans 640 90 0 0 vss
port 12 nsew ground bidirectional
flabel metal4 s 5548 1538 5708 6302 0 FreeSans 640 90 0 0 vss
port 12 nsew ground bidirectional
flabel metal4 s 7200 1538 7360 6302 0 FreeSans 640 90 0 0 vss
port 12 nsew ground bidirectional
rlabel metal1 3976 5880 3976 5880 0 vdd
rlabel via1 4016 6272 4016 6272 0 vss
rlabel metal2 2100 1036 2100 1036 0 INmb
rlabel metal2 952 1708 952 1708 0 INpb
rlabel metal2 5544 1764 5544 1764 0 OUTm
rlabel metal2 3864 1708 3864 1708 0 OUTp
rlabel metal3 2744 3220 2744 3220 0 _00_
rlabel metal2 2408 2492 2408 2492 0 _01_
rlabel metal3 3080 3724 3080 3724 0 _02_
rlabel metal2 3276 2324 3276 2324 0 _03_
rlabel metal2 3780 2996 3780 2996 0 _04_
rlabel metal3 2604 2268 2604 2268 0 _05_
rlabel metal2 3276 2912 3276 2912 0 _06_
rlabel metal3 679 5964 679 5964 0 cmnmos
rlabel metal3 679 1988 679 1988 0 cmpmos
rlabel metal3 2548 2156 2548 2156 0 net1
rlabel metal2 3220 3332 3220 3332 0 net10
rlabel metal2 1988 6076 1988 6076 0 net11
rlabel metal2 2548 2380 2548 2380 0 net2
rlabel metal2 3948 2128 3948 2128 0 net3
rlabel metal3 3948 2156 3948 2156 0 net4
rlabel metal2 2212 3220 2212 3220 0 net5
rlabel metal2 2408 3836 2408 3836 0 net6
rlabel metal2 1540 2352 1540 2352 0 net7
rlabel metal3 4732 3836 4732 3836 0 net8
rlabel metal2 3500 3920 3500 3920 0 net9
rlabel metal3 6748 1708 6748 1708 0 oe
rlabel metal3 6468 5740 6468 5740 0 omnmos
rlabel metal3 5180 6020 5180 6020 0 ompmos
rlabel metal3 3220 6020 3220 6020 0 opnmos
rlabel metal2 1120 6132 1120 6132 0 oppmos
<< properties >>
string FIXED_BBOX 0 0 8000 8000
<< end >>
