magic
tech gf180mcuC
magscale 1 5
timestamp 1670265865
<< obsm1 >>
rect 672 855 99288 98422
<< metal2 >>
rect 1904 99600 1960 100000
rect 5600 99600 5656 100000
rect 9296 99600 9352 100000
rect 12992 99600 13048 100000
rect 16688 99600 16744 100000
rect 20384 99600 20440 100000
rect 24080 99600 24136 100000
rect 27776 99600 27832 100000
rect 31472 99600 31528 100000
rect 35168 99600 35224 100000
rect 38864 99600 38920 100000
rect 42560 99600 42616 100000
rect 46256 99600 46312 100000
rect 49952 99600 50008 100000
rect 53648 99600 53704 100000
rect 57344 99600 57400 100000
rect 61040 99600 61096 100000
rect 64736 99600 64792 100000
rect 68432 99600 68488 100000
rect 72128 99600 72184 100000
rect 75824 99600 75880 100000
rect 79520 99600 79576 100000
rect 83216 99600 83272 100000
rect 86912 99600 86968 100000
rect 90608 99600 90664 100000
rect 94304 99600 94360 100000
rect 98000 99600 98056 100000
rect 7952 0 8008 400
rect 8232 0 8288 400
rect 8512 0 8568 400
rect 8792 0 8848 400
rect 9072 0 9128 400
rect 9352 0 9408 400
rect 9632 0 9688 400
rect 9912 0 9968 400
rect 10192 0 10248 400
rect 10472 0 10528 400
rect 10752 0 10808 400
rect 11032 0 11088 400
rect 11312 0 11368 400
rect 11592 0 11648 400
rect 11872 0 11928 400
rect 12152 0 12208 400
rect 12432 0 12488 400
rect 12712 0 12768 400
rect 12992 0 13048 400
rect 13272 0 13328 400
rect 13552 0 13608 400
rect 13832 0 13888 400
rect 14112 0 14168 400
rect 14392 0 14448 400
rect 14672 0 14728 400
rect 14952 0 15008 400
rect 15232 0 15288 400
rect 15512 0 15568 400
rect 15792 0 15848 400
rect 16072 0 16128 400
rect 16352 0 16408 400
rect 16632 0 16688 400
rect 16912 0 16968 400
rect 17192 0 17248 400
rect 17472 0 17528 400
rect 17752 0 17808 400
rect 18032 0 18088 400
rect 18312 0 18368 400
rect 18592 0 18648 400
rect 18872 0 18928 400
rect 19152 0 19208 400
rect 19432 0 19488 400
rect 19712 0 19768 400
rect 19992 0 20048 400
rect 20272 0 20328 400
rect 20552 0 20608 400
rect 20832 0 20888 400
rect 21112 0 21168 400
rect 21392 0 21448 400
rect 21672 0 21728 400
rect 21952 0 22008 400
rect 22232 0 22288 400
rect 22512 0 22568 400
rect 22792 0 22848 400
rect 23072 0 23128 400
rect 23352 0 23408 400
rect 23632 0 23688 400
rect 23912 0 23968 400
rect 24192 0 24248 400
rect 24472 0 24528 400
rect 24752 0 24808 400
rect 25032 0 25088 400
rect 25312 0 25368 400
rect 25592 0 25648 400
rect 25872 0 25928 400
rect 26152 0 26208 400
rect 26432 0 26488 400
rect 26712 0 26768 400
rect 26992 0 27048 400
rect 27272 0 27328 400
rect 27552 0 27608 400
rect 27832 0 27888 400
rect 28112 0 28168 400
rect 28392 0 28448 400
rect 28672 0 28728 400
rect 28952 0 29008 400
rect 29232 0 29288 400
rect 29512 0 29568 400
rect 29792 0 29848 400
rect 30072 0 30128 400
rect 30352 0 30408 400
rect 30632 0 30688 400
rect 30912 0 30968 400
rect 31192 0 31248 400
rect 31472 0 31528 400
rect 31752 0 31808 400
rect 32032 0 32088 400
rect 32312 0 32368 400
rect 32592 0 32648 400
rect 32872 0 32928 400
rect 33152 0 33208 400
rect 33432 0 33488 400
rect 33712 0 33768 400
rect 33992 0 34048 400
rect 34272 0 34328 400
rect 34552 0 34608 400
rect 34832 0 34888 400
rect 35112 0 35168 400
rect 35392 0 35448 400
rect 35672 0 35728 400
rect 35952 0 36008 400
rect 36232 0 36288 400
rect 36512 0 36568 400
rect 36792 0 36848 400
rect 37072 0 37128 400
rect 37352 0 37408 400
rect 37632 0 37688 400
rect 37912 0 37968 400
rect 38192 0 38248 400
rect 38472 0 38528 400
rect 38752 0 38808 400
rect 39032 0 39088 400
rect 39312 0 39368 400
rect 39592 0 39648 400
rect 39872 0 39928 400
rect 40152 0 40208 400
rect 40432 0 40488 400
rect 40712 0 40768 400
rect 40992 0 41048 400
rect 41272 0 41328 400
rect 41552 0 41608 400
rect 41832 0 41888 400
rect 42112 0 42168 400
rect 42392 0 42448 400
rect 42672 0 42728 400
rect 42952 0 43008 400
rect 43232 0 43288 400
rect 43512 0 43568 400
rect 43792 0 43848 400
rect 44072 0 44128 400
rect 44352 0 44408 400
rect 44632 0 44688 400
rect 44912 0 44968 400
rect 45192 0 45248 400
rect 45472 0 45528 400
rect 45752 0 45808 400
rect 46032 0 46088 400
rect 46312 0 46368 400
rect 46592 0 46648 400
rect 46872 0 46928 400
rect 47152 0 47208 400
rect 47432 0 47488 400
rect 47712 0 47768 400
rect 47992 0 48048 400
rect 48272 0 48328 400
rect 48552 0 48608 400
rect 48832 0 48888 400
rect 49112 0 49168 400
rect 49392 0 49448 400
rect 49672 0 49728 400
rect 49952 0 50008 400
rect 50232 0 50288 400
rect 50512 0 50568 400
rect 50792 0 50848 400
rect 51072 0 51128 400
rect 51352 0 51408 400
rect 51632 0 51688 400
rect 51912 0 51968 400
rect 52192 0 52248 400
rect 52472 0 52528 400
rect 52752 0 52808 400
rect 53032 0 53088 400
rect 53312 0 53368 400
rect 53592 0 53648 400
rect 53872 0 53928 400
rect 54152 0 54208 400
rect 54432 0 54488 400
rect 54712 0 54768 400
rect 54992 0 55048 400
rect 55272 0 55328 400
rect 55552 0 55608 400
rect 55832 0 55888 400
rect 56112 0 56168 400
rect 56392 0 56448 400
rect 56672 0 56728 400
rect 56952 0 57008 400
rect 57232 0 57288 400
rect 57512 0 57568 400
rect 57792 0 57848 400
rect 58072 0 58128 400
rect 58352 0 58408 400
rect 58632 0 58688 400
rect 58912 0 58968 400
rect 59192 0 59248 400
rect 59472 0 59528 400
rect 59752 0 59808 400
rect 60032 0 60088 400
rect 60312 0 60368 400
rect 60592 0 60648 400
rect 60872 0 60928 400
rect 61152 0 61208 400
rect 61432 0 61488 400
rect 61712 0 61768 400
rect 61992 0 62048 400
rect 62272 0 62328 400
rect 62552 0 62608 400
rect 62832 0 62888 400
rect 63112 0 63168 400
rect 63392 0 63448 400
rect 63672 0 63728 400
rect 63952 0 64008 400
rect 64232 0 64288 400
rect 64512 0 64568 400
rect 64792 0 64848 400
rect 65072 0 65128 400
rect 65352 0 65408 400
rect 65632 0 65688 400
rect 65912 0 65968 400
rect 66192 0 66248 400
rect 66472 0 66528 400
rect 66752 0 66808 400
rect 67032 0 67088 400
rect 67312 0 67368 400
rect 67592 0 67648 400
rect 67872 0 67928 400
rect 68152 0 68208 400
rect 68432 0 68488 400
rect 68712 0 68768 400
rect 68992 0 69048 400
rect 69272 0 69328 400
rect 69552 0 69608 400
rect 69832 0 69888 400
rect 70112 0 70168 400
rect 70392 0 70448 400
rect 70672 0 70728 400
rect 70952 0 71008 400
rect 71232 0 71288 400
rect 71512 0 71568 400
rect 71792 0 71848 400
rect 72072 0 72128 400
rect 72352 0 72408 400
rect 72632 0 72688 400
rect 72912 0 72968 400
rect 73192 0 73248 400
rect 73472 0 73528 400
rect 73752 0 73808 400
rect 74032 0 74088 400
rect 74312 0 74368 400
rect 74592 0 74648 400
rect 74872 0 74928 400
rect 75152 0 75208 400
rect 75432 0 75488 400
rect 75712 0 75768 400
rect 75992 0 76048 400
rect 76272 0 76328 400
rect 76552 0 76608 400
rect 76832 0 76888 400
rect 77112 0 77168 400
rect 77392 0 77448 400
rect 77672 0 77728 400
rect 77952 0 78008 400
rect 78232 0 78288 400
rect 78512 0 78568 400
rect 78792 0 78848 400
rect 79072 0 79128 400
rect 79352 0 79408 400
rect 79632 0 79688 400
rect 79912 0 79968 400
rect 80192 0 80248 400
rect 80472 0 80528 400
rect 80752 0 80808 400
rect 81032 0 81088 400
rect 81312 0 81368 400
rect 81592 0 81648 400
rect 81872 0 81928 400
rect 82152 0 82208 400
rect 82432 0 82488 400
rect 82712 0 82768 400
rect 82992 0 83048 400
rect 83272 0 83328 400
rect 83552 0 83608 400
rect 83832 0 83888 400
rect 84112 0 84168 400
rect 84392 0 84448 400
rect 84672 0 84728 400
rect 84952 0 85008 400
rect 85232 0 85288 400
rect 85512 0 85568 400
rect 85792 0 85848 400
rect 86072 0 86128 400
rect 86352 0 86408 400
rect 86632 0 86688 400
rect 86912 0 86968 400
rect 87192 0 87248 400
rect 87472 0 87528 400
rect 87752 0 87808 400
rect 88032 0 88088 400
rect 88312 0 88368 400
rect 88592 0 88648 400
rect 88872 0 88928 400
rect 89152 0 89208 400
rect 89432 0 89488 400
rect 89712 0 89768 400
rect 89992 0 90048 400
rect 90272 0 90328 400
rect 90552 0 90608 400
rect 90832 0 90888 400
rect 91112 0 91168 400
rect 91392 0 91448 400
rect 91672 0 91728 400
rect 91952 0 92008 400
<< obsm2 >>
rect 798 99570 1874 99666
rect 1990 99570 5570 99666
rect 5686 99570 9266 99666
rect 9382 99570 12962 99666
rect 13078 99570 16658 99666
rect 16774 99570 20354 99666
rect 20470 99570 24050 99666
rect 24166 99570 27746 99666
rect 27862 99570 31442 99666
rect 31558 99570 35138 99666
rect 35254 99570 38834 99666
rect 38950 99570 42530 99666
rect 42646 99570 46226 99666
rect 46342 99570 49922 99666
rect 50038 99570 53618 99666
rect 53734 99570 57314 99666
rect 57430 99570 61010 99666
rect 61126 99570 64706 99666
rect 64822 99570 68402 99666
rect 68518 99570 72098 99666
rect 72214 99570 75794 99666
rect 75910 99570 79490 99666
rect 79606 99570 83186 99666
rect 83302 99570 86882 99666
rect 86998 99570 90578 99666
rect 90694 99570 94274 99666
rect 94390 99570 97970 99666
rect 98086 99570 99162 99666
rect 798 430 99162 99570
rect 798 400 7922 430
rect 8038 400 8202 430
rect 8318 400 8482 430
rect 8598 400 8762 430
rect 8878 400 9042 430
rect 9158 400 9322 430
rect 9438 400 9602 430
rect 9718 400 9882 430
rect 9998 400 10162 430
rect 10278 400 10442 430
rect 10558 400 10722 430
rect 10838 400 11002 430
rect 11118 400 11282 430
rect 11398 400 11562 430
rect 11678 400 11842 430
rect 11958 400 12122 430
rect 12238 400 12402 430
rect 12518 400 12682 430
rect 12798 400 12962 430
rect 13078 400 13242 430
rect 13358 400 13522 430
rect 13638 400 13802 430
rect 13918 400 14082 430
rect 14198 400 14362 430
rect 14478 400 14642 430
rect 14758 400 14922 430
rect 15038 400 15202 430
rect 15318 400 15482 430
rect 15598 400 15762 430
rect 15878 400 16042 430
rect 16158 400 16322 430
rect 16438 400 16602 430
rect 16718 400 16882 430
rect 16998 400 17162 430
rect 17278 400 17442 430
rect 17558 400 17722 430
rect 17838 400 18002 430
rect 18118 400 18282 430
rect 18398 400 18562 430
rect 18678 400 18842 430
rect 18958 400 19122 430
rect 19238 400 19402 430
rect 19518 400 19682 430
rect 19798 400 19962 430
rect 20078 400 20242 430
rect 20358 400 20522 430
rect 20638 400 20802 430
rect 20918 400 21082 430
rect 21198 400 21362 430
rect 21478 400 21642 430
rect 21758 400 21922 430
rect 22038 400 22202 430
rect 22318 400 22482 430
rect 22598 400 22762 430
rect 22878 400 23042 430
rect 23158 400 23322 430
rect 23438 400 23602 430
rect 23718 400 23882 430
rect 23998 400 24162 430
rect 24278 400 24442 430
rect 24558 400 24722 430
rect 24838 400 25002 430
rect 25118 400 25282 430
rect 25398 400 25562 430
rect 25678 400 25842 430
rect 25958 400 26122 430
rect 26238 400 26402 430
rect 26518 400 26682 430
rect 26798 400 26962 430
rect 27078 400 27242 430
rect 27358 400 27522 430
rect 27638 400 27802 430
rect 27918 400 28082 430
rect 28198 400 28362 430
rect 28478 400 28642 430
rect 28758 400 28922 430
rect 29038 400 29202 430
rect 29318 400 29482 430
rect 29598 400 29762 430
rect 29878 400 30042 430
rect 30158 400 30322 430
rect 30438 400 30602 430
rect 30718 400 30882 430
rect 30998 400 31162 430
rect 31278 400 31442 430
rect 31558 400 31722 430
rect 31838 400 32002 430
rect 32118 400 32282 430
rect 32398 400 32562 430
rect 32678 400 32842 430
rect 32958 400 33122 430
rect 33238 400 33402 430
rect 33518 400 33682 430
rect 33798 400 33962 430
rect 34078 400 34242 430
rect 34358 400 34522 430
rect 34638 400 34802 430
rect 34918 400 35082 430
rect 35198 400 35362 430
rect 35478 400 35642 430
rect 35758 400 35922 430
rect 36038 400 36202 430
rect 36318 400 36482 430
rect 36598 400 36762 430
rect 36878 400 37042 430
rect 37158 400 37322 430
rect 37438 400 37602 430
rect 37718 400 37882 430
rect 37998 400 38162 430
rect 38278 400 38442 430
rect 38558 400 38722 430
rect 38838 400 39002 430
rect 39118 400 39282 430
rect 39398 400 39562 430
rect 39678 400 39842 430
rect 39958 400 40122 430
rect 40238 400 40402 430
rect 40518 400 40682 430
rect 40798 400 40962 430
rect 41078 400 41242 430
rect 41358 400 41522 430
rect 41638 400 41802 430
rect 41918 400 42082 430
rect 42198 400 42362 430
rect 42478 400 42642 430
rect 42758 400 42922 430
rect 43038 400 43202 430
rect 43318 400 43482 430
rect 43598 400 43762 430
rect 43878 400 44042 430
rect 44158 400 44322 430
rect 44438 400 44602 430
rect 44718 400 44882 430
rect 44998 400 45162 430
rect 45278 400 45442 430
rect 45558 400 45722 430
rect 45838 400 46002 430
rect 46118 400 46282 430
rect 46398 400 46562 430
rect 46678 400 46842 430
rect 46958 400 47122 430
rect 47238 400 47402 430
rect 47518 400 47682 430
rect 47798 400 47962 430
rect 48078 400 48242 430
rect 48358 400 48522 430
rect 48638 400 48802 430
rect 48918 400 49082 430
rect 49198 400 49362 430
rect 49478 400 49642 430
rect 49758 400 49922 430
rect 50038 400 50202 430
rect 50318 400 50482 430
rect 50598 400 50762 430
rect 50878 400 51042 430
rect 51158 400 51322 430
rect 51438 400 51602 430
rect 51718 400 51882 430
rect 51998 400 52162 430
rect 52278 400 52442 430
rect 52558 400 52722 430
rect 52838 400 53002 430
rect 53118 400 53282 430
rect 53398 400 53562 430
rect 53678 400 53842 430
rect 53958 400 54122 430
rect 54238 400 54402 430
rect 54518 400 54682 430
rect 54798 400 54962 430
rect 55078 400 55242 430
rect 55358 400 55522 430
rect 55638 400 55802 430
rect 55918 400 56082 430
rect 56198 400 56362 430
rect 56478 400 56642 430
rect 56758 400 56922 430
rect 57038 400 57202 430
rect 57318 400 57482 430
rect 57598 400 57762 430
rect 57878 400 58042 430
rect 58158 400 58322 430
rect 58438 400 58602 430
rect 58718 400 58882 430
rect 58998 400 59162 430
rect 59278 400 59442 430
rect 59558 400 59722 430
rect 59838 400 60002 430
rect 60118 400 60282 430
rect 60398 400 60562 430
rect 60678 400 60842 430
rect 60958 400 61122 430
rect 61238 400 61402 430
rect 61518 400 61682 430
rect 61798 400 61962 430
rect 62078 400 62242 430
rect 62358 400 62522 430
rect 62638 400 62802 430
rect 62918 400 63082 430
rect 63198 400 63362 430
rect 63478 400 63642 430
rect 63758 400 63922 430
rect 64038 400 64202 430
rect 64318 400 64482 430
rect 64598 400 64762 430
rect 64878 400 65042 430
rect 65158 400 65322 430
rect 65438 400 65602 430
rect 65718 400 65882 430
rect 65998 400 66162 430
rect 66278 400 66442 430
rect 66558 400 66722 430
rect 66838 400 67002 430
rect 67118 400 67282 430
rect 67398 400 67562 430
rect 67678 400 67842 430
rect 67958 400 68122 430
rect 68238 400 68402 430
rect 68518 400 68682 430
rect 68798 400 68962 430
rect 69078 400 69242 430
rect 69358 400 69522 430
rect 69638 400 69802 430
rect 69918 400 70082 430
rect 70198 400 70362 430
rect 70478 400 70642 430
rect 70758 400 70922 430
rect 71038 400 71202 430
rect 71318 400 71482 430
rect 71598 400 71762 430
rect 71878 400 72042 430
rect 72158 400 72322 430
rect 72438 400 72602 430
rect 72718 400 72882 430
rect 72998 400 73162 430
rect 73278 400 73442 430
rect 73558 400 73722 430
rect 73838 400 74002 430
rect 74118 400 74282 430
rect 74398 400 74562 430
rect 74678 400 74842 430
rect 74958 400 75122 430
rect 75238 400 75402 430
rect 75518 400 75682 430
rect 75798 400 75962 430
rect 76078 400 76242 430
rect 76358 400 76522 430
rect 76638 400 76802 430
rect 76918 400 77082 430
rect 77198 400 77362 430
rect 77478 400 77642 430
rect 77758 400 77922 430
rect 78038 400 78202 430
rect 78318 400 78482 430
rect 78598 400 78762 430
rect 78878 400 79042 430
rect 79158 400 79322 430
rect 79438 400 79602 430
rect 79718 400 79882 430
rect 79998 400 80162 430
rect 80278 400 80442 430
rect 80558 400 80722 430
rect 80838 400 81002 430
rect 81118 400 81282 430
rect 81398 400 81562 430
rect 81678 400 81842 430
rect 81958 400 82122 430
rect 82238 400 82402 430
rect 82518 400 82682 430
rect 82798 400 82962 430
rect 83078 400 83242 430
rect 83358 400 83522 430
rect 83638 400 83802 430
rect 83918 400 84082 430
rect 84198 400 84362 430
rect 84478 400 84642 430
rect 84758 400 84922 430
rect 85038 400 85202 430
rect 85318 400 85482 430
rect 85598 400 85762 430
rect 85878 400 86042 430
rect 86158 400 86322 430
rect 86438 400 86602 430
rect 86718 400 86882 430
rect 86998 400 87162 430
rect 87278 400 87442 430
rect 87558 400 87722 430
rect 87838 400 88002 430
rect 88118 400 88282 430
rect 88398 400 88562 430
rect 88678 400 88842 430
rect 88958 400 89122 430
rect 89238 400 89402 430
rect 89518 400 89682 430
rect 89798 400 89962 430
rect 90078 400 90242 430
rect 90358 400 90522 430
rect 90638 400 90802 430
rect 90918 400 91082 430
rect 91198 400 91362 430
rect 91478 400 91642 430
rect 91758 400 91922 430
rect 92038 400 99162 430
<< metal3 >>
rect 0 98168 400 98224
rect 99600 98000 100000 98056
rect 0 95816 400 95872
rect 99600 95816 100000 95872
rect 99600 93632 100000 93688
rect 0 93464 400 93520
rect 99600 91448 100000 91504
rect 0 91112 400 91168
rect 99600 89264 100000 89320
rect 0 88760 400 88816
rect 99600 87080 100000 87136
rect 0 86408 400 86464
rect 99600 84896 100000 84952
rect 0 84056 400 84112
rect 99600 82712 100000 82768
rect 0 81704 400 81760
rect 99600 80528 100000 80584
rect 0 79352 400 79408
rect 99600 78344 100000 78400
rect 0 77000 400 77056
rect 99600 76160 100000 76216
rect 0 74648 400 74704
rect 99600 73976 100000 74032
rect 0 72296 400 72352
rect 99600 71792 100000 71848
rect 0 69944 400 70000
rect 99600 69608 100000 69664
rect 0 67592 400 67648
rect 99600 67424 100000 67480
rect 0 65240 400 65296
rect 99600 65240 100000 65296
rect 99600 63056 100000 63112
rect 0 62888 400 62944
rect 99600 60872 100000 60928
rect 0 60536 400 60592
rect 99600 58688 100000 58744
rect 0 58184 400 58240
rect 99600 56504 100000 56560
rect 0 55832 400 55888
rect 99600 54320 100000 54376
rect 0 53480 400 53536
rect 99600 52136 100000 52192
rect 0 51128 400 51184
rect 99600 49952 100000 50008
rect 0 48776 400 48832
rect 99600 47768 100000 47824
rect 0 46424 400 46480
rect 99600 45584 100000 45640
rect 0 44072 400 44128
rect 99600 43400 100000 43456
rect 0 41720 400 41776
rect 99600 41216 100000 41272
rect 0 39368 400 39424
rect 99600 39032 100000 39088
rect 0 37016 400 37072
rect 99600 36848 100000 36904
rect 0 34664 400 34720
rect 99600 34664 100000 34720
rect 99600 32480 100000 32536
rect 0 32312 400 32368
rect 99600 30296 100000 30352
rect 0 29960 400 30016
rect 99600 28112 100000 28168
rect 0 27608 400 27664
rect 99600 25928 100000 25984
rect 0 25256 400 25312
rect 99600 23744 100000 23800
rect 0 22904 400 22960
rect 99600 21560 100000 21616
rect 0 20552 400 20608
rect 99600 19376 100000 19432
rect 0 18200 400 18256
rect 99600 17192 100000 17248
rect 0 15848 400 15904
rect 99600 15008 100000 15064
rect 0 13496 400 13552
rect 99600 12824 100000 12880
rect 0 11144 400 11200
rect 99600 10640 100000 10696
rect 0 8792 400 8848
rect 99600 8456 100000 8512
rect 0 6440 400 6496
rect 99600 6272 100000 6328
rect 0 4088 400 4144
rect 99600 4088 100000 4144
rect 99600 1904 100000 1960
rect 0 1736 400 1792
<< obsm3 >>
rect 400 98254 99666 98406
rect 430 98138 99666 98254
rect 400 98086 99666 98138
rect 400 97970 99570 98086
rect 400 95902 99666 97970
rect 430 95786 99570 95902
rect 400 93718 99666 95786
rect 400 93602 99570 93718
rect 400 93550 99666 93602
rect 430 93434 99666 93550
rect 400 91534 99666 93434
rect 400 91418 99570 91534
rect 400 91198 99666 91418
rect 430 91082 99666 91198
rect 400 89350 99666 91082
rect 400 89234 99570 89350
rect 400 88846 99666 89234
rect 430 88730 99666 88846
rect 400 87166 99666 88730
rect 400 87050 99570 87166
rect 400 86494 99666 87050
rect 430 86378 99666 86494
rect 400 84982 99666 86378
rect 400 84866 99570 84982
rect 400 84142 99666 84866
rect 430 84026 99666 84142
rect 400 82798 99666 84026
rect 400 82682 99570 82798
rect 400 81790 99666 82682
rect 430 81674 99666 81790
rect 400 80614 99666 81674
rect 400 80498 99570 80614
rect 400 79438 99666 80498
rect 430 79322 99666 79438
rect 400 78430 99666 79322
rect 400 78314 99570 78430
rect 400 77086 99666 78314
rect 430 76970 99666 77086
rect 400 76246 99666 76970
rect 400 76130 99570 76246
rect 400 74734 99666 76130
rect 430 74618 99666 74734
rect 400 74062 99666 74618
rect 400 73946 99570 74062
rect 400 72382 99666 73946
rect 430 72266 99666 72382
rect 400 71878 99666 72266
rect 400 71762 99570 71878
rect 400 70030 99666 71762
rect 430 69914 99666 70030
rect 400 69694 99666 69914
rect 400 69578 99570 69694
rect 400 67678 99666 69578
rect 430 67562 99666 67678
rect 400 67510 99666 67562
rect 400 67394 99570 67510
rect 400 65326 99666 67394
rect 430 65210 99570 65326
rect 400 63142 99666 65210
rect 400 63026 99570 63142
rect 400 62974 99666 63026
rect 430 62858 99666 62974
rect 400 60958 99666 62858
rect 400 60842 99570 60958
rect 400 60622 99666 60842
rect 430 60506 99666 60622
rect 400 58774 99666 60506
rect 400 58658 99570 58774
rect 400 58270 99666 58658
rect 430 58154 99666 58270
rect 400 56590 99666 58154
rect 400 56474 99570 56590
rect 400 55918 99666 56474
rect 430 55802 99666 55918
rect 400 54406 99666 55802
rect 400 54290 99570 54406
rect 400 53566 99666 54290
rect 430 53450 99666 53566
rect 400 52222 99666 53450
rect 400 52106 99570 52222
rect 400 51214 99666 52106
rect 430 51098 99666 51214
rect 400 50038 99666 51098
rect 400 49922 99570 50038
rect 400 48862 99666 49922
rect 430 48746 99666 48862
rect 400 47854 99666 48746
rect 400 47738 99570 47854
rect 400 46510 99666 47738
rect 430 46394 99666 46510
rect 400 45670 99666 46394
rect 400 45554 99570 45670
rect 400 44158 99666 45554
rect 430 44042 99666 44158
rect 400 43486 99666 44042
rect 400 43370 99570 43486
rect 400 41806 99666 43370
rect 430 41690 99666 41806
rect 400 41302 99666 41690
rect 400 41186 99570 41302
rect 400 39454 99666 41186
rect 430 39338 99666 39454
rect 400 39118 99666 39338
rect 400 39002 99570 39118
rect 400 37102 99666 39002
rect 430 36986 99666 37102
rect 400 36934 99666 36986
rect 400 36818 99570 36934
rect 400 34750 99666 36818
rect 430 34634 99570 34750
rect 400 32566 99666 34634
rect 400 32450 99570 32566
rect 400 32398 99666 32450
rect 430 32282 99666 32398
rect 400 30382 99666 32282
rect 400 30266 99570 30382
rect 400 30046 99666 30266
rect 430 29930 99666 30046
rect 400 28198 99666 29930
rect 400 28082 99570 28198
rect 400 27694 99666 28082
rect 430 27578 99666 27694
rect 400 26014 99666 27578
rect 400 25898 99570 26014
rect 400 25342 99666 25898
rect 430 25226 99666 25342
rect 400 23830 99666 25226
rect 400 23714 99570 23830
rect 400 22990 99666 23714
rect 430 22874 99666 22990
rect 400 21646 99666 22874
rect 400 21530 99570 21646
rect 400 20638 99666 21530
rect 430 20522 99666 20638
rect 400 19462 99666 20522
rect 400 19346 99570 19462
rect 400 18286 99666 19346
rect 430 18170 99666 18286
rect 400 17278 99666 18170
rect 400 17162 99570 17278
rect 400 15934 99666 17162
rect 430 15818 99666 15934
rect 400 15094 99666 15818
rect 400 14978 99570 15094
rect 400 13582 99666 14978
rect 430 13466 99666 13582
rect 400 12910 99666 13466
rect 400 12794 99570 12910
rect 400 11230 99666 12794
rect 430 11114 99666 11230
rect 400 10726 99666 11114
rect 400 10610 99570 10726
rect 400 8878 99666 10610
rect 430 8762 99666 8878
rect 400 8542 99666 8762
rect 400 8426 99570 8542
rect 400 6526 99666 8426
rect 430 6410 99666 6526
rect 400 6358 99666 6410
rect 400 6242 99570 6358
rect 400 4174 99666 6242
rect 430 4058 99570 4174
rect 400 1990 99666 4058
rect 400 1874 99570 1990
rect 400 1822 99666 1874
rect 430 1706 99666 1822
rect 400 1554 99666 1706
<< metal4 >>
rect 2224 1538 2384 98422
rect 9904 1538 10064 98422
rect 17584 1538 17744 98422
rect 25264 1538 25424 98422
rect 32944 1538 33104 98422
rect 40624 1538 40784 98422
rect 48304 1538 48464 98422
rect 55984 1538 56144 98422
rect 63664 1538 63824 98422
rect 71344 1538 71504 98422
rect 79024 1538 79184 98422
rect 86704 1538 86864 98422
rect 94384 1538 94544 98422
<< obsm4 >>
rect 3318 31873 9874 69375
rect 10094 31873 17554 69375
rect 17774 31873 25234 69375
rect 25454 31873 25522 69375
<< labels >>
rlabel metal3 s 99600 1904 100000 1960 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 99600 67424 100000 67480 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 99600 73976 100000 74032 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 99600 80528 100000 80584 6 io_in[12]
port 4 nsew signal input
rlabel metal3 s 99600 87080 100000 87136 6 io_in[13]
port 5 nsew signal input
rlabel metal3 s 99600 93632 100000 93688 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 98000 99600 98056 100000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 86912 99600 86968 100000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 75824 99600 75880 100000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 64736 99600 64792 100000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 53648 99600 53704 100000 6 io_in[19]
port 11 nsew signal input
rlabel metal3 s 99600 8456 100000 8512 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 42560 99600 42616 100000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 31472 99600 31528 100000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 20384 99600 20440 100000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 9296 99600 9352 100000 6 io_in[23]
port 16 nsew signal input
rlabel metal3 s 0 98168 400 98224 6 io_in[24]
port 17 nsew signal input
rlabel metal3 s 0 91112 400 91168 6 io_in[25]
port 18 nsew signal input
rlabel metal3 s 0 84056 400 84112 6 io_in[26]
port 19 nsew signal input
rlabel metal3 s 0 77000 400 77056 6 io_in[27]
port 20 nsew signal input
rlabel metal3 s 0 69944 400 70000 6 io_in[28]
port 21 nsew signal input
rlabel metal3 s 0 62888 400 62944 6 io_in[29]
port 22 nsew signal input
rlabel metal3 s 99600 15008 100000 15064 6 io_in[2]
port 23 nsew signal input
rlabel metal3 s 0 55832 400 55888 6 io_in[30]
port 24 nsew signal input
rlabel metal3 s 0 48776 400 48832 6 io_in[31]
port 25 nsew signal input
rlabel metal3 s 0 41720 400 41776 6 io_in[32]
port 26 nsew signal input
rlabel metal3 s 0 34664 400 34720 6 io_in[33]
port 27 nsew signal input
rlabel metal3 s 0 27608 400 27664 6 io_in[34]
port 28 nsew signal input
rlabel metal3 s 0 20552 400 20608 6 io_in[35]
port 29 nsew signal input
rlabel metal3 s 0 13496 400 13552 6 io_in[36]
port 30 nsew signal input
rlabel metal3 s 0 6440 400 6496 6 io_in[37]
port 31 nsew signal input
rlabel metal3 s 99600 21560 100000 21616 6 io_in[3]
port 32 nsew signal input
rlabel metal3 s 99600 28112 100000 28168 6 io_in[4]
port 33 nsew signal input
rlabel metal3 s 99600 34664 100000 34720 6 io_in[5]
port 34 nsew signal input
rlabel metal3 s 99600 41216 100000 41272 6 io_in[6]
port 35 nsew signal input
rlabel metal3 s 99600 47768 100000 47824 6 io_in[7]
port 36 nsew signal input
rlabel metal3 s 99600 54320 100000 54376 6 io_in[8]
port 37 nsew signal input
rlabel metal3 s 99600 60872 100000 60928 6 io_in[9]
port 38 nsew signal input
rlabel metal3 s 99600 6272 100000 6328 6 io_oeb[0]
port 39 nsew signal output
rlabel metal3 s 99600 71792 100000 71848 6 io_oeb[10]
port 40 nsew signal output
rlabel metal3 s 99600 78344 100000 78400 6 io_oeb[11]
port 41 nsew signal output
rlabel metal3 s 99600 84896 100000 84952 6 io_oeb[12]
port 42 nsew signal output
rlabel metal3 s 99600 91448 100000 91504 6 io_oeb[13]
port 43 nsew signal output
rlabel metal3 s 99600 98000 100000 98056 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 90608 99600 90664 100000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 79520 99600 79576 100000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 68432 99600 68488 100000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 57344 99600 57400 100000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 46256 99600 46312 100000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal3 s 99600 12824 100000 12880 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 35168 99600 35224 100000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 24080 99600 24136 100000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 12992 99600 13048 100000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 1904 99600 1960 100000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal3 s 0 93464 400 93520 6 io_oeb[24]
port 55 nsew signal output
rlabel metal3 s 0 86408 400 86464 6 io_oeb[25]
port 56 nsew signal output
rlabel metal3 s 0 79352 400 79408 6 io_oeb[26]
port 57 nsew signal output
rlabel metal3 s 0 72296 400 72352 6 io_oeb[27]
port 58 nsew signal output
rlabel metal3 s 0 65240 400 65296 6 io_oeb[28]
port 59 nsew signal output
rlabel metal3 s 0 58184 400 58240 6 io_oeb[29]
port 60 nsew signal output
rlabel metal3 s 99600 19376 100000 19432 6 io_oeb[2]
port 61 nsew signal output
rlabel metal3 s 0 51128 400 51184 6 io_oeb[30]
port 62 nsew signal output
rlabel metal3 s 0 44072 400 44128 6 io_oeb[31]
port 63 nsew signal output
rlabel metal3 s 0 37016 400 37072 6 io_oeb[32]
port 64 nsew signal output
rlabel metal3 s 0 29960 400 30016 6 io_oeb[33]
port 65 nsew signal output
rlabel metal3 s 0 22904 400 22960 6 io_oeb[34]
port 66 nsew signal output
rlabel metal3 s 0 15848 400 15904 6 io_oeb[35]
port 67 nsew signal output
rlabel metal3 s 0 8792 400 8848 6 io_oeb[36]
port 68 nsew signal output
rlabel metal3 s 0 1736 400 1792 6 io_oeb[37]
port 69 nsew signal output
rlabel metal3 s 99600 25928 100000 25984 6 io_oeb[3]
port 70 nsew signal output
rlabel metal3 s 99600 32480 100000 32536 6 io_oeb[4]
port 71 nsew signal output
rlabel metal3 s 99600 39032 100000 39088 6 io_oeb[5]
port 72 nsew signal output
rlabel metal3 s 99600 45584 100000 45640 6 io_oeb[6]
port 73 nsew signal output
rlabel metal3 s 99600 52136 100000 52192 6 io_oeb[7]
port 74 nsew signal output
rlabel metal3 s 99600 58688 100000 58744 6 io_oeb[8]
port 75 nsew signal output
rlabel metal3 s 99600 65240 100000 65296 6 io_oeb[9]
port 76 nsew signal output
rlabel metal3 s 99600 4088 100000 4144 6 io_out[0]
port 77 nsew signal output
rlabel metal3 s 99600 69608 100000 69664 6 io_out[10]
port 78 nsew signal output
rlabel metal3 s 99600 76160 100000 76216 6 io_out[11]
port 79 nsew signal output
rlabel metal3 s 99600 82712 100000 82768 6 io_out[12]
port 80 nsew signal output
rlabel metal3 s 99600 89264 100000 89320 6 io_out[13]
port 81 nsew signal output
rlabel metal3 s 99600 95816 100000 95872 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 94304 99600 94360 100000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 83216 99600 83272 100000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 72128 99600 72184 100000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 61040 99600 61096 100000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 49952 99600 50008 100000 6 io_out[19]
port 87 nsew signal output
rlabel metal3 s 99600 10640 100000 10696 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 38864 99600 38920 100000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 27776 99600 27832 100000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 16688 99600 16744 100000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 5600 99600 5656 100000 6 io_out[23]
port 92 nsew signal output
rlabel metal3 s 0 95816 400 95872 6 io_out[24]
port 93 nsew signal output
rlabel metal3 s 0 88760 400 88816 6 io_out[25]
port 94 nsew signal output
rlabel metal3 s 0 81704 400 81760 6 io_out[26]
port 95 nsew signal output
rlabel metal3 s 0 74648 400 74704 6 io_out[27]
port 96 nsew signal output
rlabel metal3 s 0 67592 400 67648 6 io_out[28]
port 97 nsew signal output
rlabel metal3 s 0 60536 400 60592 6 io_out[29]
port 98 nsew signal output
rlabel metal3 s 99600 17192 100000 17248 6 io_out[2]
port 99 nsew signal output
rlabel metal3 s 0 53480 400 53536 6 io_out[30]
port 100 nsew signal output
rlabel metal3 s 0 46424 400 46480 6 io_out[31]
port 101 nsew signal output
rlabel metal3 s 0 39368 400 39424 6 io_out[32]
port 102 nsew signal output
rlabel metal3 s 0 32312 400 32368 6 io_out[33]
port 103 nsew signal output
rlabel metal3 s 0 25256 400 25312 6 io_out[34]
port 104 nsew signal output
rlabel metal3 s 0 18200 400 18256 6 io_out[35]
port 105 nsew signal output
rlabel metal3 s 0 11144 400 11200 6 io_out[36]
port 106 nsew signal output
rlabel metal3 s 0 4088 400 4144 6 io_out[37]
port 107 nsew signal output
rlabel metal3 s 99600 23744 100000 23800 6 io_out[3]
port 108 nsew signal output
rlabel metal3 s 99600 30296 100000 30352 6 io_out[4]
port 109 nsew signal output
rlabel metal3 s 99600 36848 100000 36904 6 io_out[5]
port 110 nsew signal output
rlabel metal3 s 99600 43400 100000 43456 6 io_out[6]
port 111 nsew signal output
rlabel metal3 s 99600 49952 100000 50008 6 io_out[7]
port 112 nsew signal output
rlabel metal3 s 99600 56504 100000 56560 6 io_out[8]
port 113 nsew signal output
rlabel metal3 s 99600 63056 100000 63112 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 91392 0 91448 400 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 91672 0 91728 400 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 91952 0 92008 400 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 37632 0 37688 400 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 46032 0 46088 400 6 la_data_in[10]
port 119 nsew signal input
rlabel metal2 s 46872 0 46928 400 6 la_data_in[11]
port 120 nsew signal input
rlabel metal2 s 47712 0 47768 400 6 la_data_in[12]
port 121 nsew signal input
rlabel metal2 s 48552 0 48608 400 6 la_data_in[13]
port 122 nsew signal input
rlabel metal2 s 49392 0 49448 400 6 la_data_in[14]
port 123 nsew signal input
rlabel metal2 s 50232 0 50288 400 6 la_data_in[15]
port 124 nsew signal input
rlabel metal2 s 51072 0 51128 400 6 la_data_in[16]
port 125 nsew signal input
rlabel metal2 s 51912 0 51968 400 6 la_data_in[17]
port 126 nsew signal input
rlabel metal2 s 52752 0 52808 400 6 la_data_in[18]
port 127 nsew signal input
rlabel metal2 s 53592 0 53648 400 6 la_data_in[19]
port 128 nsew signal input
rlabel metal2 s 38472 0 38528 400 6 la_data_in[1]
port 129 nsew signal input
rlabel metal2 s 54432 0 54488 400 6 la_data_in[20]
port 130 nsew signal input
rlabel metal2 s 55272 0 55328 400 6 la_data_in[21]
port 131 nsew signal input
rlabel metal2 s 56112 0 56168 400 6 la_data_in[22]
port 132 nsew signal input
rlabel metal2 s 56952 0 57008 400 6 la_data_in[23]
port 133 nsew signal input
rlabel metal2 s 57792 0 57848 400 6 la_data_in[24]
port 134 nsew signal input
rlabel metal2 s 58632 0 58688 400 6 la_data_in[25]
port 135 nsew signal input
rlabel metal2 s 59472 0 59528 400 6 la_data_in[26]
port 136 nsew signal input
rlabel metal2 s 60312 0 60368 400 6 la_data_in[27]
port 137 nsew signal input
rlabel metal2 s 61152 0 61208 400 6 la_data_in[28]
port 138 nsew signal input
rlabel metal2 s 61992 0 62048 400 6 la_data_in[29]
port 139 nsew signal input
rlabel metal2 s 39312 0 39368 400 6 la_data_in[2]
port 140 nsew signal input
rlabel metal2 s 62832 0 62888 400 6 la_data_in[30]
port 141 nsew signal input
rlabel metal2 s 63672 0 63728 400 6 la_data_in[31]
port 142 nsew signal input
rlabel metal2 s 64512 0 64568 400 6 la_data_in[32]
port 143 nsew signal input
rlabel metal2 s 65352 0 65408 400 6 la_data_in[33]
port 144 nsew signal input
rlabel metal2 s 66192 0 66248 400 6 la_data_in[34]
port 145 nsew signal input
rlabel metal2 s 67032 0 67088 400 6 la_data_in[35]
port 146 nsew signal input
rlabel metal2 s 67872 0 67928 400 6 la_data_in[36]
port 147 nsew signal input
rlabel metal2 s 68712 0 68768 400 6 la_data_in[37]
port 148 nsew signal input
rlabel metal2 s 69552 0 69608 400 6 la_data_in[38]
port 149 nsew signal input
rlabel metal2 s 70392 0 70448 400 6 la_data_in[39]
port 150 nsew signal input
rlabel metal2 s 40152 0 40208 400 6 la_data_in[3]
port 151 nsew signal input
rlabel metal2 s 71232 0 71288 400 6 la_data_in[40]
port 152 nsew signal input
rlabel metal2 s 72072 0 72128 400 6 la_data_in[41]
port 153 nsew signal input
rlabel metal2 s 72912 0 72968 400 6 la_data_in[42]
port 154 nsew signal input
rlabel metal2 s 73752 0 73808 400 6 la_data_in[43]
port 155 nsew signal input
rlabel metal2 s 74592 0 74648 400 6 la_data_in[44]
port 156 nsew signal input
rlabel metal2 s 75432 0 75488 400 6 la_data_in[45]
port 157 nsew signal input
rlabel metal2 s 76272 0 76328 400 6 la_data_in[46]
port 158 nsew signal input
rlabel metal2 s 77112 0 77168 400 6 la_data_in[47]
port 159 nsew signal input
rlabel metal2 s 77952 0 78008 400 6 la_data_in[48]
port 160 nsew signal input
rlabel metal2 s 78792 0 78848 400 6 la_data_in[49]
port 161 nsew signal input
rlabel metal2 s 40992 0 41048 400 6 la_data_in[4]
port 162 nsew signal input
rlabel metal2 s 79632 0 79688 400 6 la_data_in[50]
port 163 nsew signal input
rlabel metal2 s 80472 0 80528 400 6 la_data_in[51]
port 164 nsew signal input
rlabel metal2 s 81312 0 81368 400 6 la_data_in[52]
port 165 nsew signal input
rlabel metal2 s 82152 0 82208 400 6 la_data_in[53]
port 166 nsew signal input
rlabel metal2 s 82992 0 83048 400 6 la_data_in[54]
port 167 nsew signal input
rlabel metal2 s 83832 0 83888 400 6 la_data_in[55]
port 168 nsew signal input
rlabel metal2 s 84672 0 84728 400 6 la_data_in[56]
port 169 nsew signal input
rlabel metal2 s 85512 0 85568 400 6 la_data_in[57]
port 170 nsew signal input
rlabel metal2 s 86352 0 86408 400 6 la_data_in[58]
port 171 nsew signal input
rlabel metal2 s 87192 0 87248 400 6 la_data_in[59]
port 172 nsew signal input
rlabel metal2 s 41832 0 41888 400 6 la_data_in[5]
port 173 nsew signal input
rlabel metal2 s 88032 0 88088 400 6 la_data_in[60]
port 174 nsew signal input
rlabel metal2 s 88872 0 88928 400 6 la_data_in[61]
port 175 nsew signal input
rlabel metal2 s 89712 0 89768 400 6 la_data_in[62]
port 176 nsew signal input
rlabel metal2 s 90552 0 90608 400 6 la_data_in[63]
port 177 nsew signal input
rlabel metal2 s 42672 0 42728 400 6 la_data_in[6]
port 178 nsew signal input
rlabel metal2 s 43512 0 43568 400 6 la_data_in[7]
port 179 nsew signal input
rlabel metal2 s 44352 0 44408 400 6 la_data_in[8]
port 180 nsew signal input
rlabel metal2 s 45192 0 45248 400 6 la_data_in[9]
port 181 nsew signal input
rlabel metal2 s 37912 0 37968 400 6 la_data_out[0]
port 182 nsew signal output
rlabel metal2 s 46312 0 46368 400 6 la_data_out[10]
port 183 nsew signal output
rlabel metal2 s 47152 0 47208 400 6 la_data_out[11]
port 184 nsew signal output
rlabel metal2 s 47992 0 48048 400 6 la_data_out[12]
port 185 nsew signal output
rlabel metal2 s 48832 0 48888 400 6 la_data_out[13]
port 186 nsew signal output
rlabel metal2 s 49672 0 49728 400 6 la_data_out[14]
port 187 nsew signal output
rlabel metal2 s 50512 0 50568 400 6 la_data_out[15]
port 188 nsew signal output
rlabel metal2 s 51352 0 51408 400 6 la_data_out[16]
port 189 nsew signal output
rlabel metal2 s 52192 0 52248 400 6 la_data_out[17]
port 190 nsew signal output
rlabel metal2 s 53032 0 53088 400 6 la_data_out[18]
port 191 nsew signal output
rlabel metal2 s 53872 0 53928 400 6 la_data_out[19]
port 192 nsew signal output
rlabel metal2 s 38752 0 38808 400 6 la_data_out[1]
port 193 nsew signal output
rlabel metal2 s 54712 0 54768 400 6 la_data_out[20]
port 194 nsew signal output
rlabel metal2 s 55552 0 55608 400 6 la_data_out[21]
port 195 nsew signal output
rlabel metal2 s 56392 0 56448 400 6 la_data_out[22]
port 196 nsew signal output
rlabel metal2 s 57232 0 57288 400 6 la_data_out[23]
port 197 nsew signal output
rlabel metal2 s 58072 0 58128 400 6 la_data_out[24]
port 198 nsew signal output
rlabel metal2 s 58912 0 58968 400 6 la_data_out[25]
port 199 nsew signal output
rlabel metal2 s 59752 0 59808 400 6 la_data_out[26]
port 200 nsew signal output
rlabel metal2 s 60592 0 60648 400 6 la_data_out[27]
port 201 nsew signal output
rlabel metal2 s 61432 0 61488 400 6 la_data_out[28]
port 202 nsew signal output
rlabel metal2 s 62272 0 62328 400 6 la_data_out[29]
port 203 nsew signal output
rlabel metal2 s 39592 0 39648 400 6 la_data_out[2]
port 204 nsew signal output
rlabel metal2 s 63112 0 63168 400 6 la_data_out[30]
port 205 nsew signal output
rlabel metal2 s 63952 0 64008 400 6 la_data_out[31]
port 206 nsew signal output
rlabel metal2 s 64792 0 64848 400 6 la_data_out[32]
port 207 nsew signal output
rlabel metal2 s 65632 0 65688 400 6 la_data_out[33]
port 208 nsew signal output
rlabel metal2 s 66472 0 66528 400 6 la_data_out[34]
port 209 nsew signal output
rlabel metal2 s 67312 0 67368 400 6 la_data_out[35]
port 210 nsew signal output
rlabel metal2 s 68152 0 68208 400 6 la_data_out[36]
port 211 nsew signal output
rlabel metal2 s 68992 0 69048 400 6 la_data_out[37]
port 212 nsew signal output
rlabel metal2 s 69832 0 69888 400 6 la_data_out[38]
port 213 nsew signal output
rlabel metal2 s 70672 0 70728 400 6 la_data_out[39]
port 214 nsew signal output
rlabel metal2 s 40432 0 40488 400 6 la_data_out[3]
port 215 nsew signal output
rlabel metal2 s 71512 0 71568 400 6 la_data_out[40]
port 216 nsew signal output
rlabel metal2 s 72352 0 72408 400 6 la_data_out[41]
port 217 nsew signal output
rlabel metal2 s 73192 0 73248 400 6 la_data_out[42]
port 218 nsew signal output
rlabel metal2 s 74032 0 74088 400 6 la_data_out[43]
port 219 nsew signal output
rlabel metal2 s 74872 0 74928 400 6 la_data_out[44]
port 220 nsew signal output
rlabel metal2 s 75712 0 75768 400 6 la_data_out[45]
port 221 nsew signal output
rlabel metal2 s 76552 0 76608 400 6 la_data_out[46]
port 222 nsew signal output
rlabel metal2 s 77392 0 77448 400 6 la_data_out[47]
port 223 nsew signal output
rlabel metal2 s 78232 0 78288 400 6 la_data_out[48]
port 224 nsew signal output
rlabel metal2 s 79072 0 79128 400 6 la_data_out[49]
port 225 nsew signal output
rlabel metal2 s 41272 0 41328 400 6 la_data_out[4]
port 226 nsew signal output
rlabel metal2 s 79912 0 79968 400 6 la_data_out[50]
port 227 nsew signal output
rlabel metal2 s 80752 0 80808 400 6 la_data_out[51]
port 228 nsew signal output
rlabel metal2 s 81592 0 81648 400 6 la_data_out[52]
port 229 nsew signal output
rlabel metal2 s 82432 0 82488 400 6 la_data_out[53]
port 230 nsew signal output
rlabel metal2 s 83272 0 83328 400 6 la_data_out[54]
port 231 nsew signal output
rlabel metal2 s 84112 0 84168 400 6 la_data_out[55]
port 232 nsew signal output
rlabel metal2 s 84952 0 85008 400 6 la_data_out[56]
port 233 nsew signal output
rlabel metal2 s 85792 0 85848 400 6 la_data_out[57]
port 234 nsew signal output
rlabel metal2 s 86632 0 86688 400 6 la_data_out[58]
port 235 nsew signal output
rlabel metal2 s 87472 0 87528 400 6 la_data_out[59]
port 236 nsew signal output
rlabel metal2 s 42112 0 42168 400 6 la_data_out[5]
port 237 nsew signal output
rlabel metal2 s 88312 0 88368 400 6 la_data_out[60]
port 238 nsew signal output
rlabel metal2 s 89152 0 89208 400 6 la_data_out[61]
port 239 nsew signal output
rlabel metal2 s 89992 0 90048 400 6 la_data_out[62]
port 240 nsew signal output
rlabel metal2 s 90832 0 90888 400 6 la_data_out[63]
port 241 nsew signal output
rlabel metal2 s 42952 0 43008 400 6 la_data_out[6]
port 242 nsew signal output
rlabel metal2 s 43792 0 43848 400 6 la_data_out[7]
port 243 nsew signal output
rlabel metal2 s 44632 0 44688 400 6 la_data_out[8]
port 244 nsew signal output
rlabel metal2 s 45472 0 45528 400 6 la_data_out[9]
port 245 nsew signal output
rlabel metal2 s 38192 0 38248 400 6 la_oenb[0]
port 246 nsew signal input
rlabel metal2 s 46592 0 46648 400 6 la_oenb[10]
port 247 nsew signal input
rlabel metal2 s 47432 0 47488 400 6 la_oenb[11]
port 248 nsew signal input
rlabel metal2 s 48272 0 48328 400 6 la_oenb[12]
port 249 nsew signal input
rlabel metal2 s 49112 0 49168 400 6 la_oenb[13]
port 250 nsew signal input
rlabel metal2 s 49952 0 50008 400 6 la_oenb[14]
port 251 nsew signal input
rlabel metal2 s 50792 0 50848 400 6 la_oenb[15]
port 252 nsew signal input
rlabel metal2 s 51632 0 51688 400 6 la_oenb[16]
port 253 nsew signal input
rlabel metal2 s 52472 0 52528 400 6 la_oenb[17]
port 254 nsew signal input
rlabel metal2 s 53312 0 53368 400 6 la_oenb[18]
port 255 nsew signal input
rlabel metal2 s 54152 0 54208 400 6 la_oenb[19]
port 256 nsew signal input
rlabel metal2 s 39032 0 39088 400 6 la_oenb[1]
port 257 nsew signal input
rlabel metal2 s 54992 0 55048 400 6 la_oenb[20]
port 258 nsew signal input
rlabel metal2 s 55832 0 55888 400 6 la_oenb[21]
port 259 nsew signal input
rlabel metal2 s 56672 0 56728 400 6 la_oenb[22]
port 260 nsew signal input
rlabel metal2 s 57512 0 57568 400 6 la_oenb[23]
port 261 nsew signal input
rlabel metal2 s 58352 0 58408 400 6 la_oenb[24]
port 262 nsew signal input
rlabel metal2 s 59192 0 59248 400 6 la_oenb[25]
port 263 nsew signal input
rlabel metal2 s 60032 0 60088 400 6 la_oenb[26]
port 264 nsew signal input
rlabel metal2 s 60872 0 60928 400 6 la_oenb[27]
port 265 nsew signal input
rlabel metal2 s 61712 0 61768 400 6 la_oenb[28]
port 266 nsew signal input
rlabel metal2 s 62552 0 62608 400 6 la_oenb[29]
port 267 nsew signal input
rlabel metal2 s 39872 0 39928 400 6 la_oenb[2]
port 268 nsew signal input
rlabel metal2 s 63392 0 63448 400 6 la_oenb[30]
port 269 nsew signal input
rlabel metal2 s 64232 0 64288 400 6 la_oenb[31]
port 270 nsew signal input
rlabel metal2 s 65072 0 65128 400 6 la_oenb[32]
port 271 nsew signal input
rlabel metal2 s 65912 0 65968 400 6 la_oenb[33]
port 272 nsew signal input
rlabel metal2 s 66752 0 66808 400 6 la_oenb[34]
port 273 nsew signal input
rlabel metal2 s 67592 0 67648 400 6 la_oenb[35]
port 274 nsew signal input
rlabel metal2 s 68432 0 68488 400 6 la_oenb[36]
port 275 nsew signal input
rlabel metal2 s 69272 0 69328 400 6 la_oenb[37]
port 276 nsew signal input
rlabel metal2 s 70112 0 70168 400 6 la_oenb[38]
port 277 nsew signal input
rlabel metal2 s 70952 0 71008 400 6 la_oenb[39]
port 278 nsew signal input
rlabel metal2 s 40712 0 40768 400 6 la_oenb[3]
port 279 nsew signal input
rlabel metal2 s 71792 0 71848 400 6 la_oenb[40]
port 280 nsew signal input
rlabel metal2 s 72632 0 72688 400 6 la_oenb[41]
port 281 nsew signal input
rlabel metal2 s 73472 0 73528 400 6 la_oenb[42]
port 282 nsew signal input
rlabel metal2 s 74312 0 74368 400 6 la_oenb[43]
port 283 nsew signal input
rlabel metal2 s 75152 0 75208 400 6 la_oenb[44]
port 284 nsew signal input
rlabel metal2 s 75992 0 76048 400 6 la_oenb[45]
port 285 nsew signal input
rlabel metal2 s 76832 0 76888 400 6 la_oenb[46]
port 286 nsew signal input
rlabel metal2 s 77672 0 77728 400 6 la_oenb[47]
port 287 nsew signal input
rlabel metal2 s 78512 0 78568 400 6 la_oenb[48]
port 288 nsew signal input
rlabel metal2 s 79352 0 79408 400 6 la_oenb[49]
port 289 nsew signal input
rlabel metal2 s 41552 0 41608 400 6 la_oenb[4]
port 290 nsew signal input
rlabel metal2 s 80192 0 80248 400 6 la_oenb[50]
port 291 nsew signal input
rlabel metal2 s 81032 0 81088 400 6 la_oenb[51]
port 292 nsew signal input
rlabel metal2 s 81872 0 81928 400 6 la_oenb[52]
port 293 nsew signal input
rlabel metal2 s 82712 0 82768 400 6 la_oenb[53]
port 294 nsew signal input
rlabel metal2 s 83552 0 83608 400 6 la_oenb[54]
port 295 nsew signal input
rlabel metal2 s 84392 0 84448 400 6 la_oenb[55]
port 296 nsew signal input
rlabel metal2 s 85232 0 85288 400 6 la_oenb[56]
port 297 nsew signal input
rlabel metal2 s 86072 0 86128 400 6 la_oenb[57]
port 298 nsew signal input
rlabel metal2 s 86912 0 86968 400 6 la_oenb[58]
port 299 nsew signal input
rlabel metal2 s 87752 0 87808 400 6 la_oenb[59]
port 300 nsew signal input
rlabel metal2 s 42392 0 42448 400 6 la_oenb[5]
port 301 nsew signal input
rlabel metal2 s 88592 0 88648 400 6 la_oenb[60]
port 302 nsew signal input
rlabel metal2 s 89432 0 89488 400 6 la_oenb[61]
port 303 nsew signal input
rlabel metal2 s 90272 0 90328 400 6 la_oenb[62]
port 304 nsew signal input
rlabel metal2 s 91112 0 91168 400 6 la_oenb[63]
port 305 nsew signal input
rlabel metal2 s 43232 0 43288 400 6 la_oenb[6]
port 306 nsew signal input
rlabel metal2 s 44072 0 44128 400 6 la_oenb[7]
port 307 nsew signal input
rlabel metal2 s 44912 0 44968 400 6 la_oenb[8]
port 308 nsew signal input
rlabel metal2 s 45752 0 45808 400 6 la_oenb[9]
port 309 nsew signal input
rlabel metal4 s 2224 1538 2384 98422 6 vdd
port 310 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 98422 6 vdd
port 310 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 98422 6 vdd
port 310 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 98422 6 vdd
port 310 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 98422 6 vdd
port 310 nsew power bidirectional
rlabel metal4 s 79024 1538 79184 98422 6 vdd
port 310 nsew power bidirectional
rlabel metal4 s 94384 1538 94544 98422 6 vdd
port 310 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 98422 6 vss
port 311 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 98422 6 vss
port 311 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 98422 6 vss
port 311 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 98422 6 vss
port 311 nsew ground bidirectional
rlabel metal4 s 71344 1538 71504 98422 6 vss
port 311 nsew ground bidirectional
rlabel metal4 s 86704 1538 86864 98422 6 vss
port 311 nsew ground bidirectional
rlabel metal2 s 7952 0 8008 400 6 wb_clk_i
port 312 nsew signal input
rlabel metal2 s 8232 0 8288 400 6 wb_rst_i
port 313 nsew signal input
rlabel metal2 s 8512 0 8568 400 6 wbs_ack_o
port 314 nsew signal output
rlabel metal2 s 9632 0 9688 400 6 wbs_adr_i[0]
port 315 nsew signal input
rlabel metal2 s 19152 0 19208 400 6 wbs_adr_i[10]
port 316 nsew signal input
rlabel metal2 s 19992 0 20048 400 6 wbs_adr_i[11]
port 317 nsew signal input
rlabel metal2 s 20832 0 20888 400 6 wbs_adr_i[12]
port 318 nsew signal input
rlabel metal2 s 21672 0 21728 400 6 wbs_adr_i[13]
port 319 nsew signal input
rlabel metal2 s 22512 0 22568 400 6 wbs_adr_i[14]
port 320 nsew signal input
rlabel metal2 s 23352 0 23408 400 6 wbs_adr_i[15]
port 321 nsew signal input
rlabel metal2 s 24192 0 24248 400 6 wbs_adr_i[16]
port 322 nsew signal input
rlabel metal2 s 25032 0 25088 400 6 wbs_adr_i[17]
port 323 nsew signal input
rlabel metal2 s 25872 0 25928 400 6 wbs_adr_i[18]
port 324 nsew signal input
rlabel metal2 s 26712 0 26768 400 6 wbs_adr_i[19]
port 325 nsew signal input
rlabel metal2 s 10752 0 10808 400 6 wbs_adr_i[1]
port 326 nsew signal input
rlabel metal2 s 27552 0 27608 400 6 wbs_adr_i[20]
port 327 nsew signal input
rlabel metal2 s 28392 0 28448 400 6 wbs_adr_i[21]
port 328 nsew signal input
rlabel metal2 s 29232 0 29288 400 6 wbs_adr_i[22]
port 329 nsew signal input
rlabel metal2 s 30072 0 30128 400 6 wbs_adr_i[23]
port 330 nsew signal input
rlabel metal2 s 30912 0 30968 400 6 wbs_adr_i[24]
port 331 nsew signal input
rlabel metal2 s 31752 0 31808 400 6 wbs_adr_i[25]
port 332 nsew signal input
rlabel metal2 s 32592 0 32648 400 6 wbs_adr_i[26]
port 333 nsew signal input
rlabel metal2 s 33432 0 33488 400 6 wbs_adr_i[27]
port 334 nsew signal input
rlabel metal2 s 34272 0 34328 400 6 wbs_adr_i[28]
port 335 nsew signal input
rlabel metal2 s 35112 0 35168 400 6 wbs_adr_i[29]
port 336 nsew signal input
rlabel metal2 s 11872 0 11928 400 6 wbs_adr_i[2]
port 337 nsew signal input
rlabel metal2 s 35952 0 36008 400 6 wbs_adr_i[30]
port 338 nsew signal input
rlabel metal2 s 36792 0 36848 400 6 wbs_adr_i[31]
port 339 nsew signal input
rlabel metal2 s 12992 0 13048 400 6 wbs_adr_i[3]
port 340 nsew signal input
rlabel metal2 s 14112 0 14168 400 6 wbs_adr_i[4]
port 341 nsew signal input
rlabel metal2 s 14952 0 15008 400 6 wbs_adr_i[5]
port 342 nsew signal input
rlabel metal2 s 15792 0 15848 400 6 wbs_adr_i[6]
port 343 nsew signal input
rlabel metal2 s 16632 0 16688 400 6 wbs_adr_i[7]
port 344 nsew signal input
rlabel metal2 s 17472 0 17528 400 6 wbs_adr_i[8]
port 345 nsew signal input
rlabel metal2 s 18312 0 18368 400 6 wbs_adr_i[9]
port 346 nsew signal input
rlabel metal2 s 8792 0 8848 400 6 wbs_cyc_i
port 347 nsew signal input
rlabel metal2 s 9912 0 9968 400 6 wbs_dat_i[0]
port 348 nsew signal input
rlabel metal2 s 19432 0 19488 400 6 wbs_dat_i[10]
port 349 nsew signal input
rlabel metal2 s 20272 0 20328 400 6 wbs_dat_i[11]
port 350 nsew signal input
rlabel metal2 s 21112 0 21168 400 6 wbs_dat_i[12]
port 351 nsew signal input
rlabel metal2 s 21952 0 22008 400 6 wbs_dat_i[13]
port 352 nsew signal input
rlabel metal2 s 22792 0 22848 400 6 wbs_dat_i[14]
port 353 nsew signal input
rlabel metal2 s 23632 0 23688 400 6 wbs_dat_i[15]
port 354 nsew signal input
rlabel metal2 s 24472 0 24528 400 6 wbs_dat_i[16]
port 355 nsew signal input
rlabel metal2 s 25312 0 25368 400 6 wbs_dat_i[17]
port 356 nsew signal input
rlabel metal2 s 26152 0 26208 400 6 wbs_dat_i[18]
port 357 nsew signal input
rlabel metal2 s 26992 0 27048 400 6 wbs_dat_i[19]
port 358 nsew signal input
rlabel metal2 s 11032 0 11088 400 6 wbs_dat_i[1]
port 359 nsew signal input
rlabel metal2 s 27832 0 27888 400 6 wbs_dat_i[20]
port 360 nsew signal input
rlabel metal2 s 28672 0 28728 400 6 wbs_dat_i[21]
port 361 nsew signal input
rlabel metal2 s 29512 0 29568 400 6 wbs_dat_i[22]
port 362 nsew signal input
rlabel metal2 s 30352 0 30408 400 6 wbs_dat_i[23]
port 363 nsew signal input
rlabel metal2 s 31192 0 31248 400 6 wbs_dat_i[24]
port 364 nsew signal input
rlabel metal2 s 32032 0 32088 400 6 wbs_dat_i[25]
port 365 nsew signal input
rlabel metal2 s 32872 0 32928 400 6 wbs_dat_i[26]
port 366 nsew signal input
rlabel metal2 s 33712 0 33768 400 6 wbs_dat_i[27]
port 367 nsew signal input
rlabel metal2 s 34552 0 34608 400 6 wbs_dat_i[28]
port 368 nsew signal input
rlabel metal2 s 35392 0 35448 400 6 wbs_dat_i[29]
port 369 nsew signal input
rlabel metal2 s 12152 0 12208 400 6 wbs_dat_i[2]
port 370 nsew signal input
rlabel metal2 s 36232 0 36288 400 6 wbs_dat_i[30]
port 371 nsew signal input
rlabel metal2 s 37072 0 37128 400 6 wbs_dat_i[31]
port 372 nsew signal input
rlabel metal2 s 13272 0 13328 400 6 wbs_dat_i[3]
port 373 nsew signal input
rlabel metal2 s 14392 0 14448 400 6 wbs_dat_i[4]
port 374 nsew signal input
rlabel metal2 s 15232 0 15288 400 6 wbs_dat_i[5]
port 375 nsew signal input
rlabel metal2 s 16072 0 16128 400 6 wbs_dat_i[6]
port 376 nsew signal input
rlabel metal2 s 16912 0 16968 400 6 wbs_dat_i[7]
port 377 nsew signal input
rlabel metal2 s 17752 0 17808 400 6 wbs_dat_i[8]
port 378 nsew signal input
rlabel metal2 s 18592 0 18648 400 6 wbs_dat_i[9]
port 379 nsew signal input
rlabel metal2 s 10192 0 10248 400 6 wbs_dat_o[0]
port 380 nsew signal output
rlabel metal2 s 19712 0 19768 400 6 wbs_dat_o[10]
port 381 nsew signal output
rlabel metal2 s 20552 0 20608 400 6 wbs_dat_o[11]
port 382 nsew signal output
rlabel metal2 s 21392 0 21448 400 6 wbs_dat_o[12]
port 383 nsew signal output
rlabel metal2 s 22232 0 22288 400 6 wbs_dat_o[13]
port 384 nsew signal output
rlabel metal2 s 23072 0 23128 400 6 wbs_dat_o[14]
port 385 nsew signal output
rlabel metal2 s 23912 0 23968 400 6 wbs_dat_o[15]
port 386 nsew signal output
rlabel metal2 s 24752 0 24808 400 6 wbs_dat_o[16]
port 387 nsew signal output
rlabel metal2 s 25592 0 25648 400 6 wbs_dat_o[17]
port 388 nsew signal output
rlabel metal2 s 26432 0 26488 400 6 wbs_dat_o[18]
port 389 nsew signal output
rlabel metal2 s 27272 0 27328 400 6 wbs_dat_o[19]
port 390 nsew signal output
rlabel metal2 s 11312 0 11368 400 6 wbs_dat_o[1]
port 391 nsew signal output
rlabel metal2 s 28112 0 28168 400 6 wbs_dat_o[20]
port 392 nsew signal output
rlabel metal2 s 28952 0 29008 400 6 wbs_dat_o[21]
port 393 nsew signal output
rlabel metal2 s 29792 0 29848 400 6 wbs_dat_o[22]
port 394 nsew signal output
rlabel metal2 s 30632 0 30688 400 6 wbs_dat_o[23]
port 395 nsew signal output
rlabel metal2 s 31472 0 31528 400 6 wbs_dat_o[24]
port 396 nsew signal output
rlabel metal2 s 32312 0 32368 400 6 wbs_dat_o[25]
port 397 nsew signal output
rlabel metal2 s 33152 0 33208 400 6 wbs_dat_o[26]
port 398 nsew signal output
rlabel metal2 s 33992 0 34048 400 6 wbs_dat_o[27]
port 399 nsew signal output
rlabel metal2 s 34832 0 34888 400 6 wbs_dat_o[28]
port 400 nsew signal output
rlabel metal2 s 35672 0 35728 400 6 wbs_dat_o[29]
port 401 nsew signal output
rlabel metal2 s 12432 0 12488 400 6 wbs_dat_o[2]
port 402 nsew signal output
rlabel metal2 s 36512 0 36568 400 6 wbs_dat_o[30]
port 403 nsew signal output
rlabel metal2 s 37352 0 37408 400 6 wbs_dat_o[31]
port 404 nsew signal output
rlabel metal2 s 13552 0 13608 400 6 wbs_dat_o[3]
port 405 nsew signal output
rlabel metal2 s 14672 0 14728 400 6 wbs_dat_o[4]
port 406 nsew signal output
rlabel metal2 s 15512 0 15568 400 6 wbs_dat_o[5]
port 407 nsew signal output
rlabel metal2 s 16352 0 16408 400 6 wbs_dat_o[6]
port 408 nsew signal output
rlabel metal2 s 17192 0 17248 400 6 wbs_dat_o[7]
port 409 nsew signal output
rlabel metal2 s 18032 0 18088 400 6 wbs_dat_o[8]
port 410 nsew signal output
rlabel metal2 s 18872 0 18928 400 6 wbs_dat_o[9]
port 411 nsew signal output
rlabel metal2 s 10472 0 10528 400 6 wbs_sel_i[0]
port 412 nsew signal input
rlabel metal2 s 11592 0 11648 400 6 wbs_sel_i[1]
port 413 nsew signal input
rlabel metal2 s 12712 0 12768 400 6 wbs_sel_i[2]
port 414 nsew signal input
rlabel metal2 s 13832 0 13888 400 6 wbs_sel_i[3]
port 415 nsew signal input
rlabel metal2 s 9072 0 9128 400 6 wbs_stb_i
port 416 nsew signal input
rlabel metal2 s 9352 0 9408 400 6 wbs_we_i
port 417 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 100000 100000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 7581470
string GDS_FILE /mnt/c/Users/rmprice/Documents/Github/Trollo/openlane/user_proj_example/runs/22_12_05_11_40/results/signoff/user_proj_example.magic.gds
string GDS_START 336942
<< end >>

