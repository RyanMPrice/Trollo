* NGSPICE file created from BinMultiplier.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai33_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai33_1 A1 A2 A3 B1 B2 B3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_2 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyc_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyc_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyb_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyb_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyd_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyd_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

.subckt BinMultiplier Y[0] Y[10] Y[11] Y[12] Y[13] Y[14] Y[15] Y[16] Y[17] Y[18] Y[19]
+ Y[1] Y[20] Y[21] Y[22] Y[23] Y[24] Y[25] Y[26] Y[27] Y[28] Y[29] Y[2] Y[30] Y[31]
+ Y[3] Y[4] Y[5] Y[6] Y[7] Y[8] Y[9] clk dba[0] dba[10] dba[11] dba[12] dba[13] dba[14]
+ dba[15] dba[1] dba[2] dba[3] dba[4] dba[5] dba[6] dba[7] dba[8] dba[9] dbb[0] dbb[10]
+ dbb[11] dbb[12] dbb[13] dbb[14] dbb[15] dbb[1] dbb[2] dbb[3] dbb[4] dbb[5] dbb[6]
+ dbb[7] dbb[8] dbb[9] done enable rst vdd vss yA[0] yA[10] yA[11] yA[12] yA[13] yA[14]
+ yA[15] yA[1] yA[2] yA[3] yA[4] yA[5] yA[6] yA[7] yA[8] yA[9] yB[0] yB[10] yB[11]
+ yB[12] yB[13] yB[14] yB[15] yB[1] yB[2] yB[3] yB[4] yB[5] yB[6] yB[7] yB[8] yB[9]
XTAP_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2106_ _1099_ _1153_ _1154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_27_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2037_ _1045_ _1078_ _1079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_10_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2182__A2 _1070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output37_I net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1445__A1 _0193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1748__A2 _0787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2173__A2 _1226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1684__A1 _1040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1389__I net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2724_ _0366_ _0410_ _0431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2655_ _0318_ _0342_ _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1606_ _1375_ _0526_ _0648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2586_ _0278_ _0283_ _0284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1537_ _0560_ _0578_ _0579_ _0580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1468_ _0428_ _0461_ _0492_ _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_1399_ _1116_ _1138_ _1149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1675__A1 _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2467__A3 _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2155__A2 _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1666__A1 net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1418__A1 _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2440_ net18 net3 _0126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2146__A2 _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2371_ _0043_ _0051_ _0052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_37_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2082__A1 _1050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2385__A2 _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2707_ _0360_ _0381_ _0412_ _0413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2638_ _0334_ _0338_ _0339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2569_ _0241_ _0264_ _0265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1896__A1 _0864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2300__A2 net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1940_ _0364_ _0661_ _0977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2064__A1 net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1871_ _0908_ _0909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2367__A2 _1380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2423_ _0598_ _1009_ _1351_ _0108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2354_ _1350_ _1351_ _0034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1878__A1 net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2285_ _1201_ _1344_ _1345_ _1346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_40_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1802__A1 _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1869__A1 _1127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1869__B2 net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2046__A1 _1192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2070_ _0214_ _0813_ _1114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1923_ _0884_ _0897_ _0960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1397__I net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1854_ net5 _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1785_ _0810_ _0823_ _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__2760__A2 _1384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2406_ _0086_ _0089_ _0090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2337_ _0013_ _0015_ _0016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2268_ _1324_ _1327_ _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_38_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2199_ _1164_ _1173_ _1162_ _1254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_25_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2028__A1 net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2579__A2 _1383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2751__A2 _0300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1711__B1 _0692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1490__A2 _0214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1570_ _0528_ _0611_ _0612_ _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_6_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2122_ _0798_ _0801_ _1170_ _1165_ _1172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_19_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2053_ _1031_ _1095_ _1096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__2258__A1 _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1906_ _0874_ _0881_ _0942_ _0943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1855__I _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1837_ _0095_ _0661_ _0875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1768_ _0745_ _0754_ _0807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1699_ _0689_ _0696_ _0739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1590__I net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2497__A1 net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2421__A1 _0049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput42 net42 Y[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput53 net53 Y[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput64 net64 Y[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput75 net75 yA[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput86 net86 yB[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__2488__A1 _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput97 net97 yB[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2660__A1 _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2740_ _0430_ _0431_ _0445_ _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_8_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2671_ _0814_ _1383_ _1384_ _0747_ _0374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1622_ _0659_ _0663_ _0664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1553_ _0593_ _0594_ _0595_ _0596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1484_ _0524_ _0527_ _0528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2105_ _1120_ _1152_ _1153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2036_ _1047_ _1077_ _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_35_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1914__B1 _0692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1693__A2 _0671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1445__A2 _0247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1684__A2 _0724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2723_ _0400_ _0429_ _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2149__B1 net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2654_ _0320_ _0341_ _0356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1605_ net8 _0584_ _0647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2585_ _0280_ _0281_ _0282_ _0283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_1536_ _0562_ _0577_ _0579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1467_ _1051_ _0482_ _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1398_ _1127_ _1138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__1675__A2 _0568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2467__A4 _0107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2321__B1 _1384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2019_ _0982_ _0986_ _1059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2624__A1 _0274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1666__A2 _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1418__A2 _1116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2615__A1 _0305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2091__A2 net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2370_ net15 net20 _0051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1657__A2 _0665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2706_ _0362_ _0379_ _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2637_ _0335_ _0337_ _0338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__1593__A1 _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2568_ _0246_ _0264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2499_ _0567_ net23 _0190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1519_ _0538_ _0542_ _0561_ _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input29_I dbb[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output97_I net97 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2064__A2 net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1870_ _1127_ net1 _0814_ _0906_ _0908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__1683__I _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2422_ _0046_ _0055_ _0105_ _0107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_36_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2353_ _1350_ _1351_ _0033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1878__A2 _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2284_ _1270_ _1343_ _1345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1802__A2 _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1999_ _0916_ _1035_ _1036_ _0953_ _1037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_4_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1869__A2 _0814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2046__A2 _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1678__I _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2037__A2 _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1922_ _0941_ _0958_ _0959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_30_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1853_ _1160_ net3 _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1548__A1 _0565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1784_ _0812_ _0822_ _0823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2405_ _0087_ _0088_ _0089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2336_ _1318_ _1328_ _0014_ _0015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2267_ _1325_ _1326_ _1253_ _1327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_37_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2198_ _1176_ _1252_ _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_25_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2028__A2 net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2751__A3 _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1711__A1 _1018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1711__B2 net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2121_ _0857_ _0928_ _1170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2052_ _1028_ _1033_ _1095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_34_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1769__A1 _0758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1905_ _0877_ _0880_ _0942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1836_ _0833_ _0871_ _0873_ _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1767_ _0739_ _0804_ _0805_ _0806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1698_ _0738_ net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1941__A1 net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2497__A2 net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2319_ _1066_ _1383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_38_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input11_I dba[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2185__A1 _1065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput43 net43 Y[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__1932__A1 net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput54 net54 Y[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput65 net65 Y[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput76 net76 yA[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput87 net87 yB[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__2488__A2 _0746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput98 net98 yB[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2670_ _0330_ _0372_ _0373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1621_ _0657_ _0660_ _0662_ _0663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_1552_ _1288_ _0471_ _0595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1483_ net1 _0526_ _0527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input3_I dba[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2479__A2 net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2104_ _1122_ _1151_ _1152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2035_ _1058_ _1076_ _1077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_23_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2799_ _0495_ _0505_ _0506_ _0509_ _0510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
X_1819_ _0802_ _0857_ _0858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2167__A1 _1048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1914__A1 _0214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1914__B2 _1375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2646__B _0294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2722_ _0409_ _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2653_ _0354_ _0351_ _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_8_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2149__A1 _1386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2149__B2 _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1604_ _1018_ _0554_ _0646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2584_ _0782_ _0906_ _0282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1535_ _0562_ _0577_ _0578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1466_ _0471_ _0482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1397_ net8 _1127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__2321__A1 _0106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2321__B2 _1299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2018_ _1049_ _1057_ _1058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_35_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output42_I net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2312__A1 _1366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2615__A2 _0306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2551__A1 _0243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2705_ _0366_ _0410_ _0411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2636_ _0321_ _0336_ _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2567_ _0243_ _0263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2542__A1 _0233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2498_ _0187_ _0188_ _0189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1518_ _0533_ _0537_ _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1449_ _0268_ _0290_ _0301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_28_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1805__B1 _0782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2533__A1 _0168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2421_ _0049_ _0054_ _0105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2352_ _0029_ _0030_ _0032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2283_ _1270_ _1343_ _1344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_29_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1998_ _0950_ _0954_ _1036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__2763__A1 _1383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2619_ _0271_ _0284_ _0319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1921_ _0943_ _0957_ _0958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1852_ _0783_ _0888_ _0889_ _0846_ _0890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_30_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1548__A2 _0570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1783_ _0815_ _0821_ _0822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2404_ _1333_ _0012_ _1314_ _1317_ _0088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2335_ _1314_ _1317_ _0014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1720__A2 _0759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2266_ _1173_ _1326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_38_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2197_ _1177_ _1179_ _1251_ _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_25_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1475__A1 _0518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2727__A1 _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2120_ _0998_ _1165_ _1168_ _1169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_13_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2051_ _1024_ _1044_ _1092_ _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_35_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1769__A2 _0787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1904_ _0939_ _0940_ _0941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1835_ _0767_ _0872_ _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1766_ _0741_ _0789_ _0805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1697_ _0683_ _0737_ _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__1941__A2 _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2318_ _0095_ _1237_ _1382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2249_ _1294_ _1306_ _1307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__1457__A1 net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1932__A2 _0584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput55 net55 Y[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput44 net44 Y[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput66 net66 done vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput88 net88 yB[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput77 net77 yA[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_17_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1620__A1 _1040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1620_ _1040_ _0661_ _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1923__A2 _0897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1551_ _1375_ _0375_ _0594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1482_ _0525_ _0526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1687__A1 _0717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2103_ _1134_ _1150_ _1151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_11_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2034_ _1060_ _1075_ _1076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_35_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2100__A2 _1146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1818_ _0803_ _0856_ _0857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2798_ _0467_ _0475_ _0493_ _0507_ _0508_ _0509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_1749_ _0755_ _0788_ _0789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_2_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1850__A1 _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1841__A1 _0526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2721_ _0388_ _0414_ _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2149__A2 _1199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2652_ _0296_ _0299_ _0347_ _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_1603_ _0642_ _0643_ _0644_ _0594_ _0645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_2583_ _0724_ _1199_ _0281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1534_ _0571_ _0576_ _0577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1465_ net12 _0471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1396_ _1105_ _1116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__2321__A2 _1383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2085__A1 _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2017_ _1053_ _1056_ _1057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_35_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1832__A1 _0837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2560__A2 _0255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output35_I net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2615__A3 _0308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2000__A1 net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2067__A1 net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1814__A1 _0837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2704_ _0400_ _0409_ _0410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2635_ _0782_ _0944_ _0336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2566_ _0219_ _0250_ _0262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2497_ net15 net22 _0188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1517_ _0552_ _0558_ _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1448_ _1310_ _0031_ _0279_ _0290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_4_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1805__A1 _1105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1805__B2 _1051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1400__I net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2230__A1 _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2533__A2 _0173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2297__A1 _1346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2420_ _0032_ _0035_ _0104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2351_ _0482_ _0598_ _0944_ net23 _0030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_2282_ _1275_ _1343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_33_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1997_ net12 _0691_ _1035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2763__A2 _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2618_ _0317_ _0318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2549_ _0603_ net23 _0244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2451__A1 net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1920_ _0949_ _0956_ _0957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1851_ _1094_ _0782_ _0848_ _1040_ _0889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1782_ _0817_ _0820_ _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_6_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2403_ _1333_ _0012_ _0087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2334_ _1333_ _0012_ _0013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2265_ _1157_ _1161_ _1325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_38_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2196_ _1189_ _1250_ _1251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_38_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1944__B1 _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1475__A2 _0519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2424__A1 _0107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2727__A2 _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2050_ _1027_ _1043_ _1092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_35_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1903_ _0910_ _0918_ _0940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1834_ net13 _0554_ _0872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1765_ _0741_ _0789_ _0804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1696_ _0733_ _0736_ _0737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2317_ _1367_ _1379_ _1380_ _1381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_2248_ _1297_ _1305_ _1306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_26_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2179_ _0554_ _0723_ _1233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1457__A2 _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput34 net34 Y[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput56 net56 Y[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput45 net45 Y[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput67 net67 yA[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA_output65_I net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput89 net89 yB[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput78 net78 yA[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1620__A2 _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1550_ _0214_ _0095_ _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1481_ net29 _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2102_ _1136_ _1148_ _1150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2033_ _1064_ _1074_ _1075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_35_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1817_ _0806_ _0855_ _0856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2797_ _1384_ _1087_ _0508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1748_ _0758_ _0787_ _0788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1679_ _1105_ _0603_ _0719_ _1051_ _0720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2627__A1 _0272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1403__I _1181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1850__A2 _0847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2094__A2 net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1841__A2 _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2720_ _0426_ net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2651_ _0351_ _0352_ net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_8_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1602_ _0593_ _0595_ _0644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2582_ _0848_ _0814_ _0280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1533_ _0572_ _0575_ _0576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1464_ _1171_ _1375_ _0461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1395_ _1094_ _1105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__2609__A1 _0305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2319__I _1066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2016_ _1048_ _1054_ _1055_ _1056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__2085__A2 _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1520__A1 _1094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2000__A2 _0746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2067__A2 _0691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1578__A1 _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2703_ _0365_ _0408_ _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2634_ _0724_ _1009_ _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2565_ _0222_ _0249_ _0261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1516_ _0552_ _0558_ _0559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1750__A1 _0739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2496_ net16 net21 _0187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1447_ _1342_ _0020_ _0279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_36_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1805__A2 _0724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2230__A2 _0747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2221__A2 _1270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2350_ _0598_ _0944_ _1009_ _0482_ _0029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2281_ _1278_ _1309_ _1340_ _1341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_37_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1996_ _1028_ _1033_ _1034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2617_ _0316_ _0287_ _0719_ _1087_ _0317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2548_ _0126_ _0233_ _0242_ _0177_ _0243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1723__A1 _0106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2479_ net30 net7 _0168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input27_I dbb[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2451__A2 net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2203__A2 _1250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1850_ _1084_ _0847_ _0888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1781_ _0749_ _0818_ _0819_ _0820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_30_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1953__A1 _0974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2402_ _0082_ _1324_ _0013_ _0086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2333_ _1334_ _1336_ _0011_ _0012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_34_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2264_ _1176_ _1320_ _1322_ _1323_ _1157_ _1161_ _1324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai33_1
XFILLER_37_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2195_ _1191_ _1249_ _1250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_37_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1979_ _0945_ _0948_ _1015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_4_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1944__A1 _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1944__B2 net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1902_ _0914_ _0917_ _0939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2179__A1 _0554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1833_ _0828_ _0834_ _0871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1764_ _0790_ _0792_ _0803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__1926__A1 net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1695_ _0734_ _0735_ _0736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2351__A1 _0482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2316_ _0584_ _0781_ _1380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2247_ _1301_ _1304_ _1305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_38_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2103__A1 _1134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2178_ _1140_ _1147_ _1231_ _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_26_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1917__A1 _0471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2590__A1 _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput57 net57 Y[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput46 net46 Y[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput35 net35 Y[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput79 net79 yA[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput68 net68 yA[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA_output58_I net58 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2645__A2 _0346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1908__A1 net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2581__A1 _0274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1480_ _0085_ _0523_ _0407_ _0386_ _0524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2101_ _1140_ _1147_ _1148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2032_ _1068_ _1072_ _1074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_35_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1816_ _0807_ _0809_ _0854_ _0855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_2796_ _1383_ _1199_ _0491_ _0507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_7_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1747_ _0771_ _0773_ _0786_ _0787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_1678_ _0661_ _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__2324__A1 _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2315__A1 _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2650_ _0313_ _0315_ _0350_ _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_9_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1601_ _0095_ _0471_ _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2554__A1 _0222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2581_ _0274_ _0277_ _0278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1532_ _0573_ _0574_ _0575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_4_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1463_ _0010_ _0428_ _0439_ _0204_ _0450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA_input1_I dba[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1394_ _1084_ _1094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_27_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2609__A2 _0306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2015_ _0525_ _0661_ _1055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2242__B1 _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2779_ _1384_ _1087_ _0433_ _0489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__2545__A1 _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1520__A2 net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2784__A1 _0446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2536__A1 _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1578__A2 _0617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2702_ _0402_ _0406_ _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2633_ _0328_ _0333_ _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2564_ _0253_ _0259_ _0252_ _0260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1515_ _0555_ _0557_ _0558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2495_ _0067_ _0176_ _0127_ _0124_ _0186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_4_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1446_ _0160_ _0258_ _0268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_28_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1569__A2 _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output40_I net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2280_ _1280_ _1308_ _1340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_1_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2748__A1 _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1995_ _1031_ _1032_ _1033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2616_ _0188_ _0316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1971__A2 _0992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2547_ _0176_ _0178_ _0242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2478_ _0123_ _0129_ _0166_ _0167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1723__A2 _0568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1429_ _1138_ _1299_ _0085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1487__A1 _1094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1478__A1 _0518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1780_ _1375_ _0632_ _0819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2401_ _1173_ _0083_ _0084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2332_ _1339_ _0009_ _0011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_27_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2263_ _1089_ _1156_ _1252_ _1175_ _1323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2194_ _1215_ _1248_ _1249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__1469__A1 _0450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1978_ _0946_ _0947_ _1014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1944__A2 _0847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1632__A1 _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1699__A1 _0689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1623__A1 _0656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1901_ _0899_ _0921_ _0937_ _0938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1832_ _0837_ _0868_ _0869_ _0870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2179__A2 _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1763_ _0798_ _0801_ _0802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1694_ _0674_ _0672_ _0735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1926__A2 _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2315_ _0632_ _0723_ _1379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2351__A2 _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2246_ _1298_ _1302_ _1303_ _1304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_2177_ _1143_ _1146_ _1231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1862__A1 _1181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1917__A2 _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2590__A2 _1009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput47 net47 Y[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput36 net36 Y[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput58 net58 Y[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput69 net69 yA[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1853__A1 _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1605__A1 net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2030__A1 net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1908__A2 _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2100_ _1143_ _1146_ _1147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2031_ _1065_ _1069_ _1071_ _1072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__2097__A1 net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2795_ _0484_ _0500_ _0498_ _0501_ _0506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1815_ _0824_ _0827_ _0853_ _0854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__2021__A1 net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1746_ _0776_ _0785_ _0786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1677_ _1094_ _0661_ _0718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2324__A2 _1066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2229_ _1139_ _1283_ _1284_ _1233_ _1285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_26_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2315__A2 _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2079__A1 _1048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2251__A1 _1280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1600_ _1299_ _0225_ _0642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2580_ _0272_ _0275_ _0276_ _0277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_1531_ _1299_ _0225_ _0106_ _1386_ _0574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1462_ _1116_ _1386_ _0225_ _1062_ _0439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2306__A2 _1367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1393_ net24 _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__2609__A3 _0308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2014_ net14 _0583_ _1054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2616__I _0188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2242__A1 net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2242__B2 _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2778_ _0467_ _0475_ _0488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1729_ _0766_ _0768_ _0769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2545__A2 _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1430__I net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2536__A2 _1066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2472__A1 _0136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2224__A1 _1230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1578__A3 _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2701_ _0403_ _0405_ _0406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_9_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2632_ _0329_ _0331_ _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2563_ _0156_ _0198_ _0259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1514_ _0527_ _0556_ _0557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2494_ _0183_ _0184_ _0185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1445_ _0193_ _0247_ _0258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_4_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2454__A1 _0136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2445__A1 net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1994_ net10 _0813_ _0905_ _1018_ _1032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2615_ _0305_ _0306_ _0308_ _0314_ _0315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_2546_ _0138_ _0240_ _0189_ _0190_ _0241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_2477_ _0119_ _0122_ _0166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1428_ _1277_ _0042_ _0074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_18_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1487__A2 _0471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2400_ _1325_ _1253_ _0082_ _0013_ _0083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_2331_ _1341_ _0008_ _0009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2262_ _1177_ _1319_ _1322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_38_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2193_ _1217_ _1247_ _1248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__2666__A1 _0747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1469__A2 _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2418__A1 _0041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1977_ _1011_ _1012_ _1013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2529_ _0220_ _0221_ _0222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input32_I dbb[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1632__A2 _0617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1900_ _0870_ _0898_ _0937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1831_ _0839_ _0852_ _0869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1762_ _0799_ _0800_ _0801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1693_ _0668_ _0671_ _0734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2314_ _1297_ _1305_ _1377_ _1378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2351__A3 _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2245_ net27 _0984_ _1303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2176_ _1220_ _1229_ _1230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_26_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1862__A2 _0814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2590__A3 _0188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput48 net48 Y[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput37 net37 Y[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput59 net59 Y[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1550__A1 _0214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1853__A2 net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1605__A2 _0584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2030__A2 _1070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2030_ net17 _1070_ _1071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2097__A2 net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2794_ _0477_ _0478_ _0497_ _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1814_ _0837_ _0839_ _0852_ _0853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__2021__A2 net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1745_ _0779_ _0784_ _0785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1676_ _0704_ _0715_ _0716_ _0717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__1780__A1 _1375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2228_ _1221_ _1234_ _1284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2159_ _1206_ _1210_ _1211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_26_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2812__I net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output63_I net63 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1523__A1 _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1530_ _1375_ _1299_ _0225_ _0106_ _0573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_1461_ _1105_ _0214_ _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1392_ _1029_ _1062_ _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2013_ _0886_ _1050_ _1052_ _0977_ _1053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_35_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2242__A2 _1066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2777_ _0477_ _0478_ _0487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1728_ _0759_ _0767_ _0768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1659_ _0651_ _0698_ _0699_ _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1505__A1 _0519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2807__I net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2481__A2 _0168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1992__A1 net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2700_ _0372_ _0404_ _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_9_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1983__A1 _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2631_ _0326_ _0330_ _0331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2562_ _0257_ net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1735__A1 _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1513_ net8 _0554_ _0556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2493_ _0137_ _0140_ _0184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_4_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1444_ _0171_ _0204_ _0236_ _0247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_36_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1974__A1 _1192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2829_ net48 net95 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_2_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1726__A1 net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1441__I net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2390__A1 _0041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2445__A2 net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1993_ _0947_ _1030_ _1031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_33_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2614_ _0302_ _0314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1708__A1 net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2545_ _0719_ _0944_ _0240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2476_ _0131_ _0143_ _0164_ _0165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1427_ _0053_ net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2820__I net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2363__A1 _1287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2330_ _1359_ _0007_ _0008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2261_ _1177_ _1319_ _1320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_38_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2192_ _1230_ _1245_ _1247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2666__A2 _1384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1976_ _0941_ _0958_ _1012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1929__A1 net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2528_ _0181_ _0194_ _0221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2459_ _0103_ _0146_ _0147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_input25_I dbb[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2815__I net64 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1830_ _0839_ _0852_ _0868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_30_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1761_ _0793_ _0794_ _0795_ _0800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2584__A1 _0782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1692_ _0684_ _0732_ _0733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_7_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2313_ _1301_ _1304_ _1377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2351__A4 net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2244_ net28 _0892_ _1302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2175_ _1223_ _1228_ _1229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_38_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1959_ _0802_ _0857_ _0928_ _0996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__2575__A1 _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput49 net49 Y[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput38 net38 Y[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__1550__A2 _0095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1838__B1 _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2566__A1 _0219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2318__A1 _0095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2793_ _0504_ net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1813_ _0842_ _0851_ _0852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_7_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1744_ _0777_ _0780_ _0783_ _0784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__2309__A1 _1362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1675_ _1288_ _0568_ _0716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1780__A2 _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1532__A2 _0574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2227_ _0526_ _0847_ _1283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2158_ _1207_ _1209_ _1210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2089_ _1068_ _1072_ _1135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2796__A1 _1383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1523__A2 _0471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output56_I net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1619__I net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2539__A1 _0747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1460_ _0386_ _0407_ _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_4_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1391_ _1051_ _1062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2012_ _0966_ _0978_ _1052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_23_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2776_ _0486_ net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1727_ net12 _0525_ _0767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1658_ _0653_ _0665_ _0699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1589_ _0582_ _0588_ _0630_ _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2823__I net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2218__B1 _0906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1992__A2 net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1432__A1 _1181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1983__A2 _0990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2630_ _0747_ _1383_ _0330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2561_ _0209_ _0256_ _0257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2492_ _0132_ _0138_ _0183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1735__A2 _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1512_ _1138_ _0526_ _0554_ _1181_ _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_4_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1443_ _1051_ _0225_ _0236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1974__A2 _1009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2828_ net47 net94 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2759_ _0440_ _0467_ _0468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1726__A2 _0584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2818__I net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1662__A1 _0586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1414__A1 _1181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1653__A1 _1138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1992_ net10 net21 _1030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2613_ _0312_ _0300_ _0313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2544_ _0224_ _0238_ _0239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__1708__A2 _0747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2381__A2 _0984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2475_ _0115_ _0130_ _0164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1426_ _1277_ _0042_ _0053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_28_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2436__A3 _0121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1644__A1 _0638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2363__A2 _0043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2260_ _1179_ _1251_ _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_34_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2191_ _1232_ _1244_ _1245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__1874__A1 net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1975_ _0943_ _0957_ _1011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1929__A2 _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2527_ _0167_ _0180_ _0220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2354__A2 _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2458_ _0110_ _0145_ _0146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__2106__A2 _1153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1409_ _1214_ _1246_ _1256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2389_ _0056_ _0058_ _0070_ _0071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA_input18_I dbb[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2290__A1 _0471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2831__I net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1856__A1 net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1760_ _0793_ _0794_ _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_30_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2584__A2 _0906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1691_ _0686_ _0731_ _0732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2312_ _1366_ _1374_ _1376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_2_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2243_ _1145_ _1298_ _1300_ _1240_ _1301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_25_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1847__A1 _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2174_ _1224_ _1227_ _1228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_15_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1958_ _0930_ _0994_ _0995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2575__A2 _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1889_ _0807_ _0925_ _0926_ _0927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xoutput39 net39 Y[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1838__A1 _0095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1838__B2 _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2826__I net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2015__A1 _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2318__A2 _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2792_ _0498_ _0502_ _0504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1812_ _0845_ _0850_ _0851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_30_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1743_ _1040_ _0782_ _0783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1674_ _0482_ _0375_ _0715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2309__A2 _1371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2226_ _1131_ _1281_ _1227_ _1224_ _1282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_38_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2157_ _1205_ _1208_ _1209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_26_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2088_ _1125_ _1133_ _1134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_41_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2245__A1 net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2796__A2 _1199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2548__A2 _0233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output49_I net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2484__A1 _0168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2539__A2 _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1390_ _1040_ _1051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2011_ net27 net3 _1050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2475__A1 _0115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2227__A1 _0526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2775_ _0465_ _0481_ _0485_ _0486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__1738__B1 _0724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1726_ net10 _0584_ _0766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1657_ _0653_ _0665_ _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1588_ _0527_ _0556_ _0589_ _0630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XTAP_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2209_ _1215_ _1248_ _1263_ _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_26_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2218__A1 _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2218__B2 _0482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1455__I net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2286__I _1282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1432__A2 _0106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2560_ _0210_ _0255_ _0256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1511_ _0553_ _0554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2491_ _0167_ _0180_ _0181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_4_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1442_ _0214_ _0225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_4_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1984__B _1020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2827_ net46 net93 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2758_ _0466_ _0444_ _0467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1709_ net9 _0691_ _0749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2689_ _0392_ _0393_ _0394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2439__A1 net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2834__I net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1662__A2 _0701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1414__A2 _1299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1653__A2 _1181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1991_ _1127_ _0944_ _1028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2602__A1 _0260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1956__A3 _0992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2612_ _0260_ _0312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2543_ _0232_ _0237_ _0238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2474_ _0030_ _0162_ _0163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1425_ _1310_ _0031_ _0042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2669__A1 _0814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2829__I net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1399__A1 _1116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2739__I _0446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2190_ _1235_ _1243_ _1244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_27_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1874__A2 _0691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1626__A2 _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1974_ _1192_ _1009_ _1010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2526_ _0185_ _0192_ _0218_ _0219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2457_ _0113_ _0144_ _0145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_29_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1408_ _1116_ _1138_ net34 _1246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2388_ _0065_ _0069_ _0070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_29_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2290__A2 _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output79_I net79 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1856__A2 _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1690_ _0697_ _0730_ _0731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_7_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2311_ _1369_ _1373_ _1374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2242_ net26 _1066_ _1237_ _1160_ _1300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_38_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1847__A2 _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2173_ _1218_ _1226_ _1227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_18_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2024__A2 net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1957_ _0933_ _0993_ _0994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1888_ _0809_ _0854_ _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2509_ _0101_ _0147_ _0200_ _0201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1535__A1 _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input30_I dbb[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1838__A2 _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2015__A2 _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1526__A1 _1040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1462__B1 _0225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1811_ _0843_ _0846_ _0849_ _0850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_31_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2791_ _0484_ _0500_ _0501_ _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_7_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1742_ _0781_ _0782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_7_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1673_ _0656_ _0664_ _0713_ _0714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1517__A1 _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2225_ _0661_ net32 _1281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2156_ net12 net20 _1208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2087_ _1129_ _1132_ _1133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__2245__A2 _0984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1508__A1 _1138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2837__I net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1741__I net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1747__A1 _0771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2172__A1 _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2010_ _0879_ _1048_ _0971_ _0969_ _1049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__1651__I _0691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2227__A2 _0847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2774_ _0483_ _0484_ _0485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1738__B2 _1062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1738__A1 _1105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1725_ _0655_ _0763_ _0764_ _0715_ _0765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_1656_ _0689_ _0696_ _0697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1587_ _0629_ net64 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2163__A1 _1136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1910__A1 net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2208_ _1217_ _1247_ _1263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2139_ _1187_ _1188_ _1189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2218__A2 _0813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output61_I net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2567__I _0243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2457__A2 _0144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2490_ _0175_ _0179_ _0180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1510_ net30 _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1441_ net11 _0214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_4_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2826_ net44 net92 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2757_ _0442_ _0466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2384__A1 _0724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1708_ net1 _0747_ _0748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2688_ _0294_ _0347_ _0393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1639_ _0680_ net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2687__A2 _0346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2439__A2 net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1466__I _0471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1990_ _1025_ _0973_ _1026_ _1027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_13_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2602__A2 _0300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2611_ _0310_ net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2366__A1 _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2542_ _0233_ _0234_ _0235_ _0237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__2118__A1 _1004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2473_ _0135_ _0142_ _0161_ _0162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2669__A2 _1384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1424_ _1342_ _0020_ _0031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_36_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2809_ net56 net75 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2357__A1 _0028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1399__A2 _1138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2348__A1 _1369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1973_ net23 _1009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2525_ _0186_ _0217_ _0218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2456_ _0131_ _0143_ _0144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1407_ _1225_ net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2387_ _0066_ _0068_ _0069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_28_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2578__A1 _0747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2310_ _1370_ _1372_ _1373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__1544__A2 _0586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2241_ net26 _1070_ _1298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2172_ _0602_ net32 _1226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1956_ _0936_ _0938_ _0992_ _0993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_1887_ _0809_ _0854_ _0925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2508_ _0103_ _0146_ _0200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2439_ net32 net4 _0125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input23_I dbb[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1526__A2 _0568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1462__B2 _1062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1462__A1 _1116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1810_ net17 _0848_ _0849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2790_ _0465_ _0481_ _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_7_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1741_ net3 _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_7_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1672_ _0659_ _0663_ _0713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2224_ _1230_ _1245_ _1279_ _1280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2155_ _0214_ _0905_ _1207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2086_ _1123_ _1130_ _1131_ _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__1453__A1 _0193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1559__I net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1939_ _0887_ _0896_ _0975_ _0976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1508__A2 _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2484__A3 _0173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2172__A2 net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2773_ _0455_ _0463_ _0484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1738__A2 _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1724_ _0704_ _0716_ _0764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_7_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1655_ _0690_ _0693_ _0695_ _0696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1586_ _0623_ _0628_ _0629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1910__A2 net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2207_ _1202_ _1261_ _1262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__1674__A1 _0482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2138_ _1183_ _1186_ _1188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2069_ _0954_ _1111_ _1112_ _1038_ _1113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_26_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2606__C _0304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output54_I net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1440_ _1029_ _1171_ _0204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1656__A1 _0689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1408__A1 _1116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2081__A1 net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2825_ net43 net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2756_ _0452_ _0449_ _0465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_8_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2384__A2 _0692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1707_ _0746_ _0747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2687_ _0391_ _0346_ _0392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1638_ _0676_ _0679_ _0680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1569_ _0530_ _0543_ _0612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2617__B _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1482__I _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1653__A4 _0692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2063__A1 _1127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1810__A1 net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2610_ _0302_ _0309_ _0310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2366__A2 _0847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2541_ _0782_ _0813_ _0235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2472_ _0136_ _0159_ _0161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1423_ _1353_ _1364_ _0010_ _0020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__1877__A1 _1018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2054__A1 _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1801__A1 _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2808_ net45 net74 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2739_ _0446_ _0447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_3_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1556__B1 _0568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2284__A1 _1270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1972_ _0936_ _1006_ _1007_ _1008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1387__I net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2524_ _0191_ _0217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2455_ _0135_ _0142_ _0143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2386_ _0047_ _0067_ _0068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1406_ _1062_ _1192_ _1225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_24_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2027__A1 _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2578__A2 _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2240_ _1283_ _1295_ _1296_ _1297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_2_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2171_ _0567_ _0691_ _1224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_18_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2009__A1 _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1955_ _0959_ _0991_ _0992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1886_ _0923_ _0924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2507_ _0156_ _0198_ _0199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2438_ _0723_ _0746_ _0124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2496__A1 net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2369_ _0567_ _0905_ _0050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input16_I dba[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2184__B1 _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2487__A1 net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2239__A1 _0554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1462__A2 _1386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1740_ _1171_ _0719_ _0780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1671_ _0703_ _0711_ _0712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_input8_I dba[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2223_ _1232_ _1244_ _1279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2154_ _1035_ _1205_ _1117_ _1114_ _1206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_2085_ _0602_ _0583_ _1131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_19_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1453__A2 _0247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1938_ _0890_ _0895_ _0975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1869_ _1127_ _0814_ _0906_ net1 _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_29_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2772_ _0427_ _0454_ _0483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__1395__I _1094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1723_ _0106_ _0568_ _0763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1654_ _0694_ _0695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1585_ _0624_ _0627_ _0628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__2699__A1 _0906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2206_ _1259_ _1260_ _1261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1674__A2 _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2137_ _1183_ _1186_ _1187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2068_ _1035_ _1039_ _1112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_41_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output47_I net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2378__B1 _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1408__A2 _1138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2081__A2 net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2824_ net42 net90 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2755_ _0464_ net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1706_ net19 _0746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2686_ _0344_ _0391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1592__A1 _1192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1637_ _0677_ _0678_ _0679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1568_ _0530_ _0543_ _0611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1499_ _0538_ _0542_ _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2617__C _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1583__A1 _0518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2063__A2 net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1810__A2 _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2540_ _0724_ _0905_ _0234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1574__A1 _0610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2471_ _0141_ _0159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1422_ _1062_ _1386_ _0010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1877__A2 _0747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1801__A2 _0568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2807_ net34 net67 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2738_ _0430_ _0431_ _0445_ _0446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2669_ _0814_ _1384_ _0372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1556__B2 _1062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1556__A1 _1116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1971_ _0938_ _0992_ _1007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__1795__A1 _0535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2523_ _0213_ _0215_ _0216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2454_ _0136_ _0141_ _0142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2385_ net32 _0781_ _0067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1405_ _1073_ _1149_ _1203_ _1214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_29_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput1 dba[0] net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_37_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2027__A2 _1065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1529__A1 _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2170_ _1050_ _1221_ _1222_ _1137_ _1223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_19_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2009__A2 _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1398__I _1127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1954_ _0962_ _0990_ _0991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__1768__A1 _0745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1885_ _0864_ _0867_ _0922_ _0923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__2193__A1 _1217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2506_ _0158_ _0197_ _0198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__1940__A1 _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2437_ _0119_ _0122_ _0123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2368_ _1296_ _0047_ _0048_ _1379_ _0049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__2496__A2 net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2299_ _1292_ _1307_ _1360_ _1361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_37_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2184__B2 _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2184__A1 _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output77_I net77 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2487__A2 net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2239__A2 _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2411__A2 _0091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1670_ _0706_ _0710_ _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_3_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2222_ _1265_ _1268_ _1276_ _1278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_38_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2153_ net13 _0746_ _1205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2084_ net14 net32 _1130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1438__B1 _1386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1937_ _0965_ _0973_ _0974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1868_ _0905_ _0906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__2166__A1 _1123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1799_ _0779_ _0784_ _0838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_1_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1913__A1 net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1591__I _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2469__A2 _0144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2771_ _0480_ _0481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_31_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1722_ _0760_ _0761_ _0762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1653_ _1138_ _1181_ _0633_ _0692_ _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_1584_ _0625_ _0626_ _0627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2699__A2 _1383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2205_ _1195_ _1213_ _1260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2136_ _1184_ _1185_ _1186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2067_ net13 _0691_ _1111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2311__A1 _1369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2378__A1 _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2378__B2 _0095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1408__A3 net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2823_ net41 net83 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2754_ _0455_ _0463_ _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2369__A1 _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1705_ _0742_ _0711_ _0744_ _0745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2685_ _0388_ _0389_ _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1636_ _0623_ _0628_ _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1567_ _1192_ _0526_ _0524_ _0610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2541__A1 _0782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1498_ _0540_ _0541_ _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_39_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2119_ _1005_ _1001_ _1166_ _1167_ _1168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_27_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2532__A1 _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2470_ _0110_ _0145_ _0157_ _0158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1421_ _1375_ _1386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__2025__I _0984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2806_ net33 clk net66 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2737_ _0442_ _0444_ _0445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2668_ _0893_ _0906_ _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1619_ net16 _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2599_ _0216_ _0251_ _0298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2806__CLK clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1774__I net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1556__A2 _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1492__A1 _1040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1970_ _0938_ _0992_ _1006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__1795__A2 _0526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2522_ _0163_ _0196_ _0215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2453_ _0137_ _0140_ _0141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2384_ _0724_ _0692_ _0066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1404_ _1171_ _1192_ _1203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
Xinput2 dba[10] net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1483__A1 net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2432__B1 _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2735__A1 _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2671__B1 _1384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2726__A1 _1383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1529__A2 _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1953_ _0974_ _0989_ _0990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_21_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1884_ _0899_ _0921_ _0922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2505_ _0163_ _0196_ _0197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__1940__A2 _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2436_ _0116_ _0120_ _0121_ _0122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_2367_ _1367_ _1380_ _0048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_29_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2298_ _1294_ _1306_ _1360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2184__A2 _1066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1695__A1 _0734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2221_ _1201_ _1270_ _1275_ _1276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_38_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2152_ _1200_ _1202_ _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_38_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2083_ _0978_ _1126_ _1128_ _1061_ _1129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_19_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1438__A1 _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1438__B2 _1062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1936_ _0968_ _0972_ _0973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1867_ net21 _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1798_ _0829_ _0836_ _0837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__1913__A2 _0691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2419_ _0038_ _0072_ _0102_ _0103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_input21_I dbb[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1677__A1 _1094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1429__A1 _1138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1601__A1 _0095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1668__A1 _1018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2093__A1 _1126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1840__A1 net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2770_ _0477_ _0479_ _0480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_12_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1721_ _0708_ _0709_ _0761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_7_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1652_ _1181_ _0692_ _0693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1583_ _0518_ _0517_ _0547_ _0618_ _0626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XTAP_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2204_ _1198_ _1212_ _1259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2135_ _1107_ _1109_ _1185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2066_ _1107_ _1109_ _1110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_26_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2084__A1 net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1867__I net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1919_ _0952_ _0955_ _0956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__1898__A1 _0904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2378__A2 _1066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1889__A1 _0807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1813__A1 _0842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2822_ net40 net73 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2753_ _0315_ _0457_ _0459_ _0462_ _0463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__2369__A2 _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1704_ _0706_ _0743_ _0744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2684_ _0356_ _0357_ _0387_ _0389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_1635_ _0621_ _0622_ _0677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1566_ _0559_ _0580_ _0608_ _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XTAP_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2541__A2 _0813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1497_ _1127_ _0375_ _0541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2118_ _1004_ _1082_ _1167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2049_ _1019_ _1080_ _1090_ _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_35_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1804__A1 _1094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2532__A2 _1070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output52_I net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2296__A1 _1349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1420_ net10 _1375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_36_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2805_ _0513_ _0514_ net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2736_ _0402_ _0406_ _0443_ _0444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2667_ _0276_ _0369_ _0331_ _0329_ _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__1565__A3 _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1618_ _1160_ _0567_ _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2598_ _0216_ _0251_ _0297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1549_ _0571_ _0576_ _0591_ _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_39_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2278__A1 _1268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2450__A1 _0568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2202__A1 _1191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1492__A2 _0535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2521_ _0212_ _0195_ _0213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2452_ _0132_ _0138_ _0140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_39_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2383_ _0061_ _0064_ _0065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1403_ _1181_ _1192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput3 dba[11] net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2680__A1 _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1483__A2 _0526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2432__A1 _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2432__B2 _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2719_ _0421_ _0425_ _0426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_3_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1538__A3 _0574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2735__A2 _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2499__A1 _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2671__A1 _0814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2671__B2 _0747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2423__A1 _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2726__A2 _1199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2662__A1 _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1952_ _0976_ _0988_ _0989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_14_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1883_ _0901_ _0920_ _0921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2504_ _0165_ _0195_ _0196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2435_ _0553_ _0984_ _0121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2366_ _0583_ _0847_ _0047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2350__B1 _1009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2297_ _1346_ _1358_ _1359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_2_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1392__A1 _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2644__A1 _0266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2220_ _1271_ _1274_ _1275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2151_ _1108_ _1201_ _1202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2082_ _1050_ _1063_ _1128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_19_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1438__A2 _1116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2635__A1 _0782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1935_ _0969_ _0971_ _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_21_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1866_ _0902_ _0836_ _0903_ _0904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1797_ _0832_ _0835_ _0836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2418_ _0041_ _0071_ _0102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2349_ _1366_ _1374_ _0027_ _0028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1677__A2 _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input14_I dba[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2626__A1 _0692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1429__A2 _1299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1601__A2 _0471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output82_I net82 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1668__A2 _0584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2093__A2 _1137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1840__A2 _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1720_ _0648_ _0759_ _0760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_7_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1651_ _0691_ _0692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__1973__I net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1582_ _0610_ _0613_ _0614_ _0625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XTAP_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input6_I dba[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2203_ _1189_ _1250_ _1257_ _1258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2134_ _1030_ _1108_ _1184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_39_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2065_ _1030_ _1108_ _1109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__2608__B2 _0255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2084__A2 net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1918_ _0950_ _0953_ _0954_ _0955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_1849_ _0875_ _0885_ _0886_ _0887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_27_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2075__A2 _1106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2821_ net39 net72 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2752_ _0354_ _0460_ _0456_ _0462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_31_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1703_ _0710_ _0743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_8_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2683_ _0356_ _0357_ _0387_ _0388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1634_ _0672_ _0675_ _0676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1565_ _0590_ _0592_ _0607_ _0608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1496_ _0523_ _0539_ _0540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2117_ _1004_ _1082_ _1166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2048_ _1021_ _1079_ _1090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1804__A2 _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1740__A1 _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output45_I net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2804_ _1062_ _1138_ _1192_ _1116_ _0514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2735_ _0848_ _1087_ _0408_ _0443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2666_ _0747_ _1384_ _0369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1617_ _0569_ _0657_ _0658_ _0601_ _0659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_2597_ _0294_ _0295_ _0296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1548_ _0565_ _0570_ _0591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1479_ _1018_ _0106_ _0523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1401__I _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1789__A1 _0471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2450__A2 net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2520_ _0165_ _0212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_5_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2451_ net15 net21 _0138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1402_ net1 _1181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2382_ _0059_ _0062_ _0063_ _0064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
Xinput4 dba[12] net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_37_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2432__A2 _1066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2718_ _0423_ _0424_ _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1943__A1 _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2649_ _0313_ _0315_ _0350_ _0351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_10_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2499__A2 net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2671__A2 _1383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2423__A2 _1009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2187__A1 net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2662__A2 _1009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1951_ _0979_ _0987_ _0988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_41_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1882_ _0904_ _0919_ _0920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2503_ _0181_ _0194_ _0195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_6_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1925__A1 _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2434_ net31 _0892_ _0120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2365_ _0044_ _0045_ _0046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2350__B2 _0482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2350__A1 _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2296_ _1349_ _1357_ _1358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_37_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2102__A1 _1136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2169__A1 _1126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1916__A1 net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1392__A2 _1062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2580__A1 _0272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2150_ _1386_ net23 _1201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2081_ net27 net4 _1126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_19_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2635__A2 _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1934_ _0963_ _0970_ _0971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_14_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1865_ _0832_ _0835_ _0903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1796_ _0828_ _0833_ _0834_ _0835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__2571__A1 _0224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2417_ _0026_ _0037_ _0100_ _0101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2323__A1 _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2348_ _1369_ _1373_ _0027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2279_ _1265_ _1337_ _1338_ _1339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_37_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2626__A2 _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1650_ net18 _0691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_8_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1581_ _0519_ _0517_ _0548_ _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_3_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2202_ _1191_ _1249_ _1257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2133_ _1102_ _1180_ _1182_ _1183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_14_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2064_ net9 net22 _1108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_19_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1917_ _0471_ _0632_ _0954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1848_ _1288_ _0723_ _0886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1595__A2 _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2544__A1 _0224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1779_ net8 _0746_ _0818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_1_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2480__B1 _1070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2535__A1 net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2820_ net38 net71 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2751_ _0312_ _0300_ _0349_ _0460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_12_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1702_ _0703_ _0742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2682_ _0382_ _0385_ _0387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1633_ _0673_ _0620_ _0674_ _0675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1564_ _0596_ _0606_ _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1495_ _1375_ _1299_ _0539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2116_ _0995_ _1083_ _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_27_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2047_ _1086_ _1088_ _1089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1568__A2 _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1740__A2 _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output38_I net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1495__A1 _1375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2803_ _1246_ _0513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2734_ _0440_ _0441_ _0442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2665_ _0363_ _0367_ _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1616_ _1040_ _0603_ _0568_ _1105_ _0658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2596_ _0261_ _0262_ _0293_ _0295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__1970__A2 _0992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1547_ _0557_ _0589_ _0590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1478_ _0518_ _0517_ _0522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_39_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1789__A2 _0554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2450_ _0568_ net22 _0137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1401_ _1160_ _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2381_ net29 _0984_ _0063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput5 dba[13] net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2717_ _0393_ _0390_ _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2196__A2 _1250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1943__A2 _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2648_ _0349_ _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2579_ _0692_ _1383_ _0276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_19_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1412__I net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2423__A3 _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1631__A1 _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2187__A2 _0984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2111__A2 _1081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1870__A1 _1127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1950_ _0982_ _0986_ _0987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_14_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1881_ _0910_ _0918_ _0919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2502_ _0185_ _0192_ _0194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2433_ _0002_ _0116_ _0118_ _0062_ _0119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__1689__A1 _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2364_ _1370_ _1372_ _0045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2350__A2 _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2295_ _1354_ _1356_ _1357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_37_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1861__A1 _0870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1613__A1 _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1916__A2 _0746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1604__A1 _1018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2080_ _0970_ _1123_ _1124_ _1054_ _1125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_16_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2096__A1 _0985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2096__B2 _1069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2148__I _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1933_ _0525_ _0602_ _0970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput30 dbb[7] net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_1864_ _0829_ _0902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1795_ _0535_ _0526_ _0834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2416_ _0028_ _0036_ _0100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2323__A2 _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2347_ _1354_ _1356_ _0026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__1531__B1 _0106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2278_ _1268_ _1276_ _1338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1834__A1 net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2011__A1 net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output68_I net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1580_ _0621_ _0622_ _0623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2305__A2 _1296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2201_ _1255_ net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2132_ _1106_ _1119_ _1182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_19_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2063_ _1127_ net23 _1107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1816__A1 _0807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2241__A1 net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1916_ net10 _0746_ _0953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1847_ _0364_ _0603_ _0885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1778_ _0816_ _0817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_1_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1807__A1 _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2480__A1 _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1420__I net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2535__A2 _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2750_ _0420_ _0458_ _0459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2774__A2 _0484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1701_ _0697_ _0730_ _0740_ _0741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_8_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2681_ _0383_ _0384_ _0385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1632_ _0609_ _0617_ _0674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_8_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1563_ _0600_ _0605_ _0606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_3_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1494_ _0533_ _0537_ _0538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2115_ _1162_ _1163_ _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2046_ _1192_ _1087_ _1017_ _1088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_10_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2214__A1 _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1495__A2 _1299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2444__A1 _0115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2802_ _0511_ net63 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2733_ _0435_ _0438_ _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2664_ _0366_ _0367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1615_ _1084_ _0602_ _0657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2595_ _0261_ _0262_ _0293_ _0294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1546_ _0582_ _0588_ _0589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1477_ _0521_ net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2029_ net7 _1070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__2435__A1 _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output50_I net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_26_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1400_ net25 _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2380_ _0553_ _0892_ _0062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput6 dba[14] net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1640__A2 _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2716_ _0354_ _0351_ _0422_ _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2647_ _0347_ _0348_ _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2578_ _0747_ _0893_ _0275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1529_ _1029_ _0375_ _0572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_19_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1631__A2 _0617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1870__A2 net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1880_ _0914_ _0917_ _0918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2501_ _0186_ _0191_ _0192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2432_ _0525_ _1066_ _1237_ _0364_ _0118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_37_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1689__A2 _0729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2363_ _1287_ _0043_ _0044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_2_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2294_ _1272_ _1355_ _1356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_37_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2638__A1 _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1861__A2 _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1613__A2 net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2629__A1 _0813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1604__A2 _0554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2203__B _1257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1932_ net13 _0584_ _0969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1863_ _0817_ _0820_ _0900_ _0901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput31 dbb[8] net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput20 dbb[12] net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1794_ net11 _0584_ _0833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2415_ _0023_ _0075_ _0099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2346_ _1359_ _0007_ _0024_ _0025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1531__A1 _1299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1531__B2 _1386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2277_ _1268_ _1276_ _1337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2087__A2 _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1834__A2 _0554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2011__A2 net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2078__A2 net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2200_ _1253_ _1254_ _1255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1513__A1 net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2131_ _1106_ _1119_ _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2062_ _1103_ _1057_ _1104_ _1106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1915_ _0819_ _0950_ _0951_ _0915_ _0952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__2241__A2 _1070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1846_ _0842_ _0851_ _0883_ _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1777_ _0690_ _0749_ _0751_ _0748_ _0816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_2329_ _1361_ _0006_ _0007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA_input12_I dba[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1807__A2 _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2480__A2 _0984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2232__A2 _1287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1991__A1 _1127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1743__A1 _1040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output80_I net80 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2680_ _0323_ _0340_ _0384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1700_ _0700_ _0729_ _0740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1631_ _0609_ _0617_ _0673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_4_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1734__A1 _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1562_ _0597_ _0601_ _0604_ _0605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XTAP_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1493_ _0531_ _0534_ _0536_ _0537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XTAP_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input4_I dba[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2114_ _1157_ _1161_ _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2045_ _1009_ _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_35_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2214__A2 _0814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1829_ _0824_ _0865_ _0866_ _0867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_38_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2150__A1 _1386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1431__I _0095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2801_ _0624_ _0627_ _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_32_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2732_ _0435_ _0438_ _0440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_8_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2663_ _0336_ _0365_ _0366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1614_ _0643_ _0654_ _0655_ _0656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_2594_ _0266_ _0292_ _0293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1545_ _0585_ _0587_ _0588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__2380__A1 _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1476_ _0517_ _0520_ _0521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_39_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2132__A1 _1106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2028_ net25 net5 _1069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2435__A2 _0984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1946__A1 _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2810__I net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2371__A1 _0043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output43_I net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2362__A1 net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput7 dba[15] net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_1
XFILLER_37_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2715_ _0395_ _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2646_ _0296_ _0299_ _0294_ _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2577_ _0173_ _0272_ _0273_ _0229_ _0274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_1528_ _0565_ _0570_ _0571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1459_ _0139_ _0397_ _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_19_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2408__A2 _0091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1616__B1 _0568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2344__A1 _1346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1870__A3 _0814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2500_ _0189_ _0190_ _0191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__2583__A1 _0724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2431_ net29 net7 _0116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2362_ net16 net19 _0043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2293_ _1271_ _1274_ _1355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_37_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2629_ _0813_ _0893_ _0329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2629__A2 _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2801__A2 _0627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2565__A1 _0222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2317__A1 _1367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1931_ _0841_ _0966_ _0967_ _0885_ _0968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_14_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1862_ _1181_ _0814_ _0821_ _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_30_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput10 dba[3] net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput21 dbb[13] net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput32 dbb[9] net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1793_ _0716_ _0830_ _0831_ _0774_ _0832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__2308__A1 net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2414_ _0025_ _0073_ _0098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1524__I net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2345_ _1361_ _0006_ _0024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1531__A2 _0225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2276_ _1262_ _1312_ _1335_ _1336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_37_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2795__A1 _0484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2538__A1 _0228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1513__A2 _0554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2130_ _1097_ _1154_ _1178_ _1179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_2061_ _1053_ _1056_ _1104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1914_ _0214_ _0633_ _0692_ _1375_ _0951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_30_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1845_ _0845_ _0850_ _0883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1776_ _1181_ _0814_ _0815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2328_ _1376_ _1378_ _0005_ _0006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_25_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2259_ _1314_ _1317_ _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_13_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2813__I net62 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1440__A1 _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1991__A2 _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1743__A2 _0782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1630_ _0668_ _0671_ _0672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1561_ _1051_ _0603_ _0604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1734__A2 _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1492_ _1040_ _0535_ _0536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_12_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2113_ _1157_ _1161_ _1162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_35_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2044_ _1014_ _1015_ _1013_ _1086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1422__A1 _1062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1828_ _0827_ _0853_ _0866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1759_ _0683_ _0737_ _0793_ _0798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_2_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2808__I net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2150__A2 net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1652__A1 _1181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2800_ _0510_ net58 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2731_ _0436_ _0437_ _0438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1404__A1 _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1955__A2 _0991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2662_ _0848_ _1009_ _0365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1613_ _1288_ net13 _0655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2593_ _0269_ _0291_ _0292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_5_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1544_ _0556_ _0586_ _0587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__2380__A2 _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1475_ _0518_ _0519_ _0520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2027_ _0894_ _1065_ _1067_ _0983_ _1068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_24_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1643__A1 _1192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1946__A2 net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_2_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1707__I _0746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1442__I _0214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1882__A1 _0904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output36_I net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput8 dba[1] net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__1873__A1 _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1625__A1 _0638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2183__I _1070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2714_ _0419_ _0420_ _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2050__A1 _1027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2645_ _0344_ _0346_ _0347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__2353__A2 _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2576_ _0226_ _0230_ _0273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1527_ _0563_ _0566_ _0569_ _0570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_1458_ _1029_ _1299_ _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_19_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1389_ net17 _1040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_28_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1616__B2 _1105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1616__A1 _1040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2821__I net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2041__A1 _1004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1870__A4 _0906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2804__B1 _1192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2280__A1 _1280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2583__A2 _1199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2430_ _0065_ _0069_ _0114_ _0115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2361_ _1376_ _0039_ _0040_ _0041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2292_ _1350_ _1351_ _1352_ _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_2_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1846__A1 _0842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2023__A1 _1050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2628_ _0230_ _0326_ _0327_ _0275_ _0328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_2559_ _0252_ _0254_ _0255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__1837__A1 _0095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2816__I net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2014__A1 net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1828__A1 _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1930_ _0875_ _0886_ _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_30_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1861_ _0870_ _0898_ _0899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
Xinput11 dba[4] net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput22 dbb[14] net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2005__A1 _1027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput33 enable net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_1792_ _0763_ _0775_ _0831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_42_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2413_ _0019_ _0076_ _0097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2344_ _1346_ _0021_ _0022_ _0023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_29_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2275_ _1264_ _1311_ _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2244__A1 net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2547__A2 _0178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2483__A1 _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2235__A1 _1282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1994__B1 _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2710__A2 _0388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2060_ _1049_ _1103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2474__A1 _0030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1913_ net11 _0691_ _0950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1844_ _0874_ _0881_ _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1775_ _0813_ _0814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2327_ _1381_ _0004_ _0005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_38_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2258_ _1093_ _1096_ _1315_ _1316_ _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_38_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2189_ _1239_ _1242_ _1243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_25_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2217__A1 _0482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1440__A2 _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2208__A1 _1217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1560_ _0602_ _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_3_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1491_ net13 _0535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2112_ _1158_ _1082_ _1159_ _1161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_2043_ _1085_ net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1422__A2 _1386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1827_ _0827_ _0853_ _0865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1758_ _0797_ net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1689_ _0700_ _0729_ _0730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_1_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2438__A1 _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2824__I net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1652__A2 _0692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1404__A2 _1192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2730_ _0403_ _0405_ _0437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2661_ _0848_ _1199_ _1009_ _0782_ _0363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_8_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1612_ _0214_ _0375_ _0654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2592_ _0285_ _0289_ _0291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_5_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1543_ net9 _0525_ _0586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1474_ _0074_ _0301_ _0519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2668__A1 _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2026_ _1084_ _0892_ _1066_ net17 _1067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_23_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2819__I net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput9 dba[2] net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_36_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2713_ _0392_ _0390_ _0417_ _0420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__1808__I net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2644_ _0266_ _0292_ _0345_ _0346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2575_ _0632_ _1237_ _0272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1526_ _1040_ _0568_ _0569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1561__A1 _1051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1457_ net1 _0375_ _0386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1388_ _1018_ _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_28_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2009_ _0602_ _0553_ _1048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1616__A2 _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1552__A1 _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2804__B2 _1116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2804__A1 _1062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1791__A1 _0106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2360_ _1378_ _0005_ _0040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1543__A1 net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2291_ _0225_ net23 _1352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_2_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2023__A2 _1061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2627_ _0272_ _0276_ _0327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2558_ _0156_ _0198_ _0253_ _0254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2489_ _0176_ _0177_ _0178_ _0179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_1509_ _0523_ _0539_ _0551_ _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input28_I dbb[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1837__A2 _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2832__I net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2014__A2 _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2317__A3 _1380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1828__A2 _0853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1860_ _0882_ _0884_ _0897_ _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
Xinput12 dba[5] net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1791_ _0106_ _0603_ _0830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput23 dbb[15] net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_6_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2412_ _0093_ _0094_ _0096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1516__A1 _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2343_ _1349_ _1357_ _0022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2274_ _1202_ _1261_ _1334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2244__A2 _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1989_ _0968_ _0972_ _1026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2180__A1 _0526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2827__I net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2483__A2 net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1994__A1 net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1994__B2 _1018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1746__A1 _0776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2171__A1 _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1912_ _0945_ _0948_ _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_30_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1843_ _0877_ _0880_ _0881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_7_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1737__A1 _1094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1774_ net20 _0813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_7_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2326_ _0000_ _0003_ _0004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2257_ _1179_ _1251_ _1316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2188_ _1236_ _1240_ _1241_ _1242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__2217__A2 _0535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1728__A1 _0759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2153__A1 net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output59_I net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1900__A1 _0870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1719__A1 net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1490_ _1171_ _0214_ _0534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2144__A1 _1110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_12_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2111_ _1008_ _1081_ _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2042_ _1003_ _1083_ _1085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_22_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1826_ _0862_ _0863_ _0864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1757_ _0793_ _0794_ _0796_ _0797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_1688_ _0712_ _0714_ _0728_ _0729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_2309_ _1362_ _1371_ _1372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__2438__A2 _0746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input10_I dba[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1456__I _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2601__A2 _0299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2660_ _0334_ _0338_ _0361_ _0362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1611_ _0596_ _0606_ _0652_ _0653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_5_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2591_ _0287_ _0288_ _0289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_4_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1542_ net1 _0584_ _0585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1473_ _0268_ _0290_ _0518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2117__A1 _1004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input2_I dba[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2668__A2 _0906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2025_ _0984_ _1066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_35_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1643__A3 _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2789_ _0465_ _0481_ _0499_ _0500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1809_ _0847_ _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__2835__I net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2056__B _1098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2712_ _0392_ _0390_ _0417_ _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_13_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2643_ _0269_ _0291_ _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2574_ _0232_ _0237_ _0270_ _0271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1525_ _0567_ _0568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__1561__A2 _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1456_ _0364_ _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_19_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1387_ net9 _1018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_35_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2008_ _0974_ _0989_ _1046_ _1047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_35_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2026__B1 _1066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2577__B2 _0229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2577__A1 _0173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1552__A2 _0471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output41_I net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2804__A2 _1138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1791__A2 _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1543__A2 _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2290_ _0471_ _0944_ _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_2_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2626_ _0692_ _1237_ _0326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2557_ _0158_ _0197_ _0253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2488_ _0781_ _0746_ _0178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1508_ _1138_ _0375_ _0540_ _0551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1439_ _1073_ _0171_ _0182_ _1364_ _0193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_28_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1461__A1 _1105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput13 dba[6] net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1790_ _0707_ _0828_ _0768_ _0766_ _0829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
Xinput24 dbb[1] net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_2411_ _0081_ _0091_ _0094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2342_ _1358_ _0021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_28_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2273_ _1187_ _1330_ _1332_ _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_25_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1452__A1 _0193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1988_ _0965_ _1025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_20_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2609_ _0305_ _0306_ _0308_ _0309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2180__A2 _0782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1443__A1 _1051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1994__A2 _0813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2171__A2 _0691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1911_ _0946_ _0947_ _0948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_30_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1434__A1 _1127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1842_ _0872_ _0878_ _0879_ _0880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_30_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1737__A2 _0724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1773_ _0762_ _0770_ _0811_ _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_6_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2325_ _1382_ _0001_ _0002_ _0003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_38_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2256_ _1179_ _1251_ _1315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_27_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2187_ net26 _0984_ _1241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1673__A1 _0656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2217__A3 _0813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2153__A2 _0746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2838__I net58 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1742__I _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1900__A2 _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1719__A2 _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2110_ _1004_ _1158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2041_ _1004_ _1005_ _1082_ _1083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_35_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1825_ _0810_ _0823_ _0863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1756_ _0683_ _0737_ _0795_ _0796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1687_ _0717_ _0727_ _0728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2308_ net15 net19 _1371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2239_ _0554_ _0781_ _1296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2071__A1 net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1885__A1 _0864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1610_ _0600_ _0605_ _0652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2590_ _0719_ _1009_ _0188_ _0288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1541_ _0583_ _0584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1472_ _0150_ _0516_ _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_5_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2024_ net24 net6 _1065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1800__A1 _0776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1808_ net4 _0847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2788_ _0483_ _0499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1739_ _0662_ _0777_ _0778_ _0722_ _0779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_39_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2283__A1 _1270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2035__A1 _1058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2711_ _0414_ _0416_ _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2642_ _0318_ _0342_ _0344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2573_ _0228_ _0231_ _0270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1524_ net14 _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1455_ net28 _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_42_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2007_ _0976_ _0988_ _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2026__A1 _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2026__B2 net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2577__A2 _0272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output34_I net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2017__A1 _1053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2008__A1 _0974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2625_ _0278_ _0283_ _0324_ _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2556_ _0211_ _0216_ _0251_ _0252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_1507_ _0550_ net62 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2487_ net2 net20 _0177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1438_ _1029_ _1116_ _1386_ _1062_ _0182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2495__A1 _0067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2486__A1 net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2238__A1 _0584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1461__A2 _0214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput14 dba[7] net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput25 dbb[2] net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2410_ _0077_ _0080_ _0093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2341_ _0017_ _0018_ _0019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2272_ _1258_ _1313_ _1332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2477__A1 _0119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1390__I _1040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1452__A2 _0247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1987_ _0949_ _0956_ _1023_ _1024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2608_ _0205_ _0303_ _0307_ _0255_ _0308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_2539_ _0747_ _0848_ _0233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input33_I enable vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1443__A2 _0225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2640__A1 _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1910_ net9 net20 _0947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1434__A2 _0106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1841_ _0526_ _0567_ _0879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1772_ _0765_ _0769_ _0811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_6_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2698__A1 _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2324_ _0364_ _1066_ _0002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2255_ _1187_ _1258_ _1313_ _1314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_38_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2186_ net27 _0892_ _1240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2217__A4 _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2040_ _1008_ _1081_ _1082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_35_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2080__A2 _1123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1824_ _0812_ _0822_ _0862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1755_ _0735_ _0733_ _0795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1686_ _0721_ _0726_ _0727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_38_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2307_ _0567_ _0813_ _1370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2238_ _0584_ _0723_ _1295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2169_ _1126_ _1139_ _1222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_26_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1949__A3 _0985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2071__A2 _0746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1582__A1 _0610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output64_I net64 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1540_ net31 _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_5_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1471_ _0353_ _0515_ _0516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_5_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2023_ _1050_ _1061_ _1063_ _1064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_35_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1807_ _1160_ _0723_ _0846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2787_ _0487_ _0497_ _0498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_2_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1738_ _1105_ _0719_ _0724_ _1062_ _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1669_ _0708_ _0709_ _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_26_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2292__A2 _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_20_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2710_ _0415_ _0388_ _0416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1794__A1 net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2641_ _0320_ _0341_ _0342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2572_ _0239_ _0248_ _0267_ _0269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1523_ _1160_ _0471_ _0566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1454_ _0160_ _0332_ _0343_ _0353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_4_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2006_ _1024_ _1044_ _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_35_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2274__A2 _1261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2026__A2 _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1776__A1 _1181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1528__A1 _0565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1700__A1 _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1388__I _1018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1767__A1 _0739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2624_ _0274_ _0277_ _0324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2192__A1 _1230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2555_ _0219_ _0250_ _0251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1506_ _0548_ _0549_ _0550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2486_ net18 net4 _0176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1437_ _1116_ _1386_ _0171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2486__A2 net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2238__A2 _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1997__A1 net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput15 dba[8] net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput26 dbb[3] net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_6_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2340_ _1339_ _0009_ _0018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2271_ _1258_ _1313_ _1330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1921__A1 _0943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2477__A2 _0122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1986_ _0952_ _1022_ _1023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2165__A1 _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2607_ _0210_ _0208_ _0307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2538_ _0228_ _0231_ _0232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2469_ _0113_ _0144_ _0157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA_input26_I dbb[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2156__A1 net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1491__I net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1840_ net12 _0583_ _0878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1771_ _0694_ _0753_ _0810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_10_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2323_ _0525_ _0893_ _0001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2698__A2 _1199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2254_ _1262_ _1312_ _1313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_38_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2185_ _1065_ _1236_ _1238_ _1144_ _1239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_38_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1969_ _0933_ _0993_ _1005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__2386__A1 _0047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2138__A1 _1183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2613__A2 _0300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2377__A1 net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2110__I _1004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2301__A1 _1226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1823_ _0806_ _0855_ _0861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2368__A1 _1296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1396__I _1105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1754_ _0734_ _0733_ _0794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1685_ _0718_ _0722_ _0725_ _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_2306_ _1234_ _1367_ _1368_ _1295_ _1369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__2540__A1 _0724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2237_ _1235_ _1243_ _1293_ _1294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2168_ _0364_ _0847_ _1221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2099_ _1141_ _1144_ _1145_ _1146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output57_I net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1470_ _0418_ _0512_ _0515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_10_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2022_ net26 _0847_ _1063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2589__A1 _0178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1806_ _0725_ _0843_ _0844_ _0780_ _0845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_2786_ _0495_ _0496_ _0497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__1854__I net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1737_ _1094_ _0724_ _0777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1668_ _1018_ _0584_ _0709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1599_ _0639_ _0640_ _0641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_38_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1794__A2 _0584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2640_ _0323_ _0340_ _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2571_ _0224_ _0238_ _0267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1522_ _0492_ _0563_ _0564_ _0534_ _0565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_1453_ _0193_ _0247_ _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2005_ _1027_ _1043_ _1044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_35_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2838_ net58 net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2769_ _0447_ _0478_ _0479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1776__A2 _0814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1528__A2 _0570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2725__A1 _0906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1700__A2 _0729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1464__A1 _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2661__B1 _1009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2623_ _0235_ _0321_ _0322_ _0281_ _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_2554_ _0222_ _0249_ _0250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1505_ _0519_ _0517_ _0549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2485_ _0170_ _0174_ _0175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1436_ _0128_ _0150_ _0160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1997__A2 _0691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput16 dba[9] net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput27 dbb[4] net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_6_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2270_ _1329_ net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_18_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1437__A1 _1116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1985_ _0955_ _1022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_9_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2606_ _1169_ _1172_ _0083_ _0304_ _0306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__2165__A2 _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2537_ _0226_ _0229_ _0230_ _0231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_2468_ _0104_ _0109_ _0155_ _0156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1419_ _1138_ _1171_ _1364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2399_ _1314_ _1317_ _0082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_input19_I dbb[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1600__A1 _1299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2156__A2 net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1667__A1 _0701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1419__A1 _1138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2092__A1 net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1947__I net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1770_ _0755_ _0788_ _0808_ _0809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_7_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1682__I net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2322_ _1241_ _1382_ _1385_ _1302_ _0000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_2253_ _1264_ _1311_ _1312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_26_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2184_ _1160_ _1066_ _1237_ _1084_ _1238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_25_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2083__B2 _1061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2386__A2 _0067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1968_ _0908_ _0935_ _1004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1899_ _0908_ _0935_ _0936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1649__A1 _1127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2074__A1 _1110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2377__A2 _1070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2129__A2 _1153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2301__A2 _1362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1822_ _0802_ _0857_ _0859_ _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2368__A2 _0047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1753_ _0790_ _0792_ _0793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1684_ _1040_ _0724_ _0725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2305_ _1283_ _1296_ _1368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__2540__A2 _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2236_ _1239_ _1242_ _1293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2167_ _1048_ _1218_ _1219_ _1130_ _1220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_2098_ net25 net6 _1145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2021_ net28 net2 _1061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2785_ _0446_ _0476_ _0494_ _0496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1805_ _1105_ _0724_ _0782_ _1051_ _0844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1736_ _0763_ _0774_ _0775_ _0776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__2210__A1 _1206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1667_ _0701_ _0707_ _0708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1598_ _0585_ _0587_ _0640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2513__A2 _0091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2277__A1 _1268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2219_ _1272_ _1273_ _1274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_26_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2440__A1 net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2570_ _0263_ _0245_ _0265_ _0266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1521_ _1105_ _0482_ _0535_ _1051_ _0564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1452_ _0193_ _0247_ _0332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_36_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2004_ _1034_ _1042_ _1043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_36_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2837_ net57 net88 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2768_ _0451_ _0449_ _0478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1719_ net11 _0553_ _0759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2699_ _0906_ _1383_ _0404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_27_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1775__I _0813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2725__A2 _1384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1464__A2 _1375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2661__B2 _0782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2661__A1 _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2622_ _0280_ _0282_ _0322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2553_ _0239_ _0248_ _0249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1504_ _0522_ _0547_ _0548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_5_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2484_ _0168_ _0172_ _0173_ _0174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_1435_ _1310_ _0139_ _0150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_24_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput17 dbb[0] net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput28 dbb[5] net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_2_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2634__A1 _0724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1437__A2 _1386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1984_ _0959_ _0991_ _1020_ _1021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2605_ _0086_ _0089_ _0304_ _0305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2536_ _0632_ _1066_ _0230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2467_ _0598_ _1087_ _1351_ _0107_ _0155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_1418_ _1029_ _1116_ _1353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2322__B1 _1385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2398_ _0077_ _0080_ _0081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_28_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1600__A2 _0225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1419__A2 _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2092__A2 _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2321_ _0106_ _1383_ _1384_ _1299_ _1385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2252_ _1278_ _1309_ _1311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2183_ _1070_ _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_19_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1658__A2 _0665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2083__A2 _1126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1967_ _1001_ _1002_ _1003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1898_ _0904_ _0919_ _0934_ _0935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2519_ _0030_ _0162_ _0211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input31_I dbb[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1821_ _0803_ _0856_ _0859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1752_ _0684_ _0732_ _0791_ _0792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1576__A1 _0610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1683_ _0723_ _0724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2304_ _0554_ _0847_ _1367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2235_ _1282_ _1291_ _1292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2166_ _1123_ _1131_ _1219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_38_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2029__I net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2097_ net26 net5 _1144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1868__I _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2056__A2 _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1567__A1 _1192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1558__A1 _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2020_ _0979_ _0987_ _1059_ _1060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_35_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2784_ _0446_ _0476_ _0494_ _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_1804_ _1094_ _0781_ _0843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1735_ _1288_ _0603_ _0775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1666_ net11 _0525_ _0707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1597_ _0556_ _0586_ _0639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_39_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2218_ _0598_ _0813_ _0906_ _0482_ _1273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2149_ _1386_ _1199_ net23 _1029_ _1200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1788__A1 _0771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output62_I net62 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1779__A1 net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2440__A2 net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1520_ _1094_ net13 _0563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1451_ _0311_ net60 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_4_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2003_ _1037_ _1041_ _1042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_23_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2431__A2 net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2836_ net55 net87 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2767_ _0476_ _0477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2195__A1 _1191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1718_ _0712_ _0756_ _0757_ _0758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2698_ _0893_ _1199_ _0403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1649_ _1127_ _0633_ _0690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2498__A2 _0188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_27_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2186__A1 net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1933__A1 _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2661__A2 _1199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2621_ _0848_ _0906_ _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2552_ _0241_ _0246_ _0248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1503_ _0544_ _0546_ _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_5_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2483_ _0583_ net6 _0173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1434_ _1127_ _0106_ _0139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2652__A2 _0299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2819_ net37 net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2168__A1 _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1679__B1 _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1851__B1 _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput18 dbb[10] net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_10_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput29 dbb[6] net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_6_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2159__A1 _1206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2095__B1 _1070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2634__A2 _1009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1983_ _0962_ _0990_ _1020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2604_ _0081_ _0153_ _0303_ _0304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_2535_ net18 _0892_ _0229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2320__I _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2466_ _0154_ net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1417_ _1321_ _1203_ _1331_ _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2397_ _1334_ _0078_ _0079_ _0080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_28_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2320_ _1237_ _1384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_2_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2251_ _1280_ _1308_ _1309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__2304__A1 _0554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2182_ net25 _1070_ _1236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_18_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1966_ _0995_ _0999_ _1002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2791__A1 _0484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1897_ _0901_ _0920_ _0934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__1594__A2 _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2518_ _0199_ _0201_ _0210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2449_ _1380_ _0125_ _0068_ _0066_ _0136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA_input24_I dbb[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1585__A2 _0627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2534__A1 _0121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1820_ _0858_ net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1751_ _0686_ _0731_ _0791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1682_ net2 _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_7_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2303_ _1363_ _1365_ _1366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_31_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2234_ _1285_ _1290_ _1291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2165_ _0583_ _0661_ _1218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2096_ _0985_ _1141_ _1142_ _1069_ _1143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_21_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2045__I _1009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1949_ _0980_ _0983_ _0985_ _0986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__1567__A2 _0526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1558__A2 _0535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2783_ _0488_ _0493_ _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1803_ _0830_ _0840_ _0841_ _0842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_1734_ _0375_ _0598_ _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1665_ _0595_ _0704_ _0705_ _0654_ _0706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_1596_ _0590_ _0636_ _0637_ _0638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_39_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2217_ _0482_ _0535_ _0813_ _0905_ _1272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_39_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2148_ _0944_ _1199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__1485__A1 _0450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2079_ _1048_ _1055_ _1124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_14_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output55_I net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1779__A2 _0746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1450_ _0074_ _0301_ _0311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_4_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2002_ _1035_ _1038_ _1039_ _1041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__1467__A1 _1051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2835_ net54 net86 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2766_ _0468_ _0475_ _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1717_ _0714_ _0728_ _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2697_ _0373_ _0401_ _0402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_6_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1648_ _0641_ _0650_ _0688_ _0689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1579_ _0518_ _0517_ _0547_ _0619_ _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XTAP_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1458__A1 _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1402__I net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_10_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2186__A2 _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1933__A2 _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2489__A3 _0178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2620_ _0285_ _0289_ _0319_ _0320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2177__A2 _1146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2551_ _0243_ _0245_ _0246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1502_ _0150_ _0516_ _0545_ _0546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2482_ net32 net5 _0172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1924__A2 _0897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1433_ _0085_ _0117_ _0128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1688__A1 _0712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1860__A1 _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1612__A1 _0214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2818_ net36 net69 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2749_ _0419_ _0424_ _0458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2168__A2 _0847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1679__B2 _1051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1679__A1 _1105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1851__A1 _1094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1851__B2 _1040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput19 dbb[11] net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_10_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2095__B2 net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2095__A1 _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1982_ _1010_ _1017_ _1019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2603_ _0203_ _0256_ _0303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2534_ _0121_ _0226_ _0227_ _0172_ _0228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_5_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2465_ _0096_ _0153_ _0154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2396_ _1336_ _0011_ _0079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1416_ _1073_ _1149_ _1331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_3_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2086__A1 _1123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1521__B1 _0535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2077__A1 _1058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1824__A1 _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2001__A1 net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2250_ _1292_ _1307_ _1308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2304__A2 _0847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2181_ _1221_ _1233_ _1234_ _1235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__1512__B1 _0554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1965_ _0930_ _0994_ _1001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1896_ _0864_ _0931_ _0932_ _0933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2517_ _0203_ _0206_ _0208_ _0209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2448_ _0133_ _0134_ _0135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2379_ _1303_ _0059_ _0060_ _0001_ _0061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_29_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input17_I dbb[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2231__A1 _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2534__A2 _0226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1750_ _0739_ _0741_ _0789_ _0790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_1681_ _1171_ _0602_ _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2302_ _1286_ _1289_ _1365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_input9_I dba[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2233_ _1286_ _1289_ _1290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2289__A1 _0535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2164_ _1134_ _1150_ _1216_ _1217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_38_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1500__A3 _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2095_ _1084_ _0984_ _1070_ net17 _1142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_19_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1948_ net17 _0984_ _0985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1879_ _0912_ _0915_ _0916_ _0917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2204__A1 _1198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2782_ _0489_ _0491_ _0493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1802_ _1288_ _0719_ _0841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1733_ _0717_ _0727_ _0772_ _0773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1664_ _0643_ _0655_ _0705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1595_ _0592_ _0607_ _0637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2216_ _0225_ _1199_ _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2147_ _1196_ _1133_ _1197_ _1198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1485__A2 _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2078_ net30 net16 _1123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output48_I net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2001_ net13 _0632_ _1039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1467__A2 _0482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2416__A1 _0028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2834_ net53 net85 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2765_ _0472_ _0474_ _0475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_8_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1716_ _0714_ _0728_ _0756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2696_ _0371_ _0376_ _0401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1647_ _0645_ _0687_ _0688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1578_ _0609_ _0617_ _0620_ _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XTAP_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1458__A2 _1299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1630__A2 _0671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2550_ _0240_ _0244_ _0245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1501_ _0353_ _0515_ _0545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2481_ _0063_ _0168_ _0169_ _0120_ _0170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_1432_ _1181_ _0106_ _0117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1612__A2 _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2817_ net35 net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2748_ _0349_ _0456_ _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2679_ _0325_ _0339_ _0383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1679__A2 _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1413__I _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2628__A1 _0230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1851__A2 _0782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2095__A2 _0984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1981_ _1013_ _1016_ _1017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_9_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2602_ _0260_ _0300_ _0302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2533_ _0168_ _0173_ _0227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2464_ _0097_ _0152_ _0153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2395_ _1336_ _0011_ _0078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1415_ _1073_ _1149_ _1321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1530__A1 _1375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2010__A2 _1048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1521__A1 _1105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1521__B2 _1051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2001__A2 _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2180_ _0526_ _0782_ _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1512__A1 _1138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1512__B2 _1181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1815__A2 _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1964_ _1000_ net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1579__A1 _0518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1895_ _0867_ _0922_ _0932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__2612__I _0260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2516_ _0098_ _0099_ _0148_ _0202_ _0208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2447_ _0050_ _0052_ _0134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2378_ _0364_ _1066_ _1237_ _0095_ _0060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_17_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2231__A2 _0691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output78_I net78 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2222__A2 _1268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1680_ _0604_ _0718_ _0720_ _0660_ _0721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_2301_ _1226_ _1362_ _1363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1733__A1 _0717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2232_ _1281_ _1287_ _1289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__2289__A2 _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2163_ _1136_ _1148_ _1216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2094_ net24 net7 _1141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1511__I _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1947_ net6 _0984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1878_ net11 _0632_ _0916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1488__B1 _0482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1421__I _1375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1963__A1 _0995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1715__A1 _0745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2140__A1 _1122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1801_ _0364_ _0568_ _0840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2781_ _0440_ _0475_ _0490_ _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_7_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1732_ _0721_ _0726_ _0772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1954__A1 _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1663_ _0095_ _0535_ _0704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1594_ _0592_ _0607_ _0636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2215_ _1115_ _1269_ _1209_ _1207_ _1270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XANTENNA__2131__A1 _1106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2146_ _1129_ _1132_ _1197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2077_ _1058_ _1076_ _1121_ _1122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2434__A2 _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2370__A1 net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2122__A1 _0798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2000_ net11 _0746_ _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2833_ net52 net84 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2764_ _0469_ _0473_ _0474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1715_ _0745_ _0754_ _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2695_ _0398_ _0399_ _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1646_ _0649_ _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1577_ _0618_ _0619_ _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2104__A1 _1122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2129_ _1099_ _1153_ _1178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2343__A1 _1349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output60_I net60 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2646__A2 _0299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1909__A1 net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2582__A1 _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1500_ _0528_ _0530_ _0543_ _0544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_2480_ _0553_ _0984_ _1070_ net29 _0169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_5_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1431_ _0095_ _0106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xoutput90 net90 yB[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_24_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1860__A3 _0897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2816_ net65 net82 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2747_ _0422_ _0417_ _0456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__2573__A1 _0228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2678_ _0360_ _0381_ _0382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1629_ _0559_ _0669_ _0670_ _0671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2316__A1 _0584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_33_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1980_ _1014_ _1015_ _1016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_20_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2601_ _0296_ _0299_ _0300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2532_ _0583_ _1070_ _0226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2555__A1 _0219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2307__A1 _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2463_ _0149_ _0151_ _0152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2394_ _0019_ _0076_ _0077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1414_ _1181_ _1299_ _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1530__A2 _1299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1597__A2 _0586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1521__A2 _0482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2785__A1 _0446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2537__A1 _0226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1512__A2 _0526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1815__A3 _0853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1963_ _0995_ _0999_ _1000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_14_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1894_ _0867_ _0922_ _0931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__2240__A3 _1296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2515_ _0207_ net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2446_ _1371_ _0132_ _0133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2377_ net28 _1070_ _0059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2519__A1 _0030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2300_ net16 net18 _1362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2231_ _0602_ _0691_ _1287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2162_ _1195_ _1213_ _1215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__1497__A1 _1127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2093_ _1126_ _1137_ _1139_ _1140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1946_ _1160_ net4 _0983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1877_ _1018_ _0747_ _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2429_ _0061_ _0064_ _0114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input22_I dbb[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1488__A1 _1105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1488__B2 _1051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1660__A1 net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1479__A1 _1018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1800_ _0776_ _0785_ _0838_ _0839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2780_ _0472_ _0474_ _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1731_ _0762_ _0770_ _0771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__1954__A2 _0990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1662_ _0586_ _0701_ _0702_ _0647_ _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_1593_ _0631_ _0634_ _0635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2214_ _0598_ _0814_ _1269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2145_ _1125_ _1196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2076_ _1060_ _1075_ _1121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_19_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1929_ net27 _0723_ _0966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2370__A2 net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2122__A2 _0801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2832_ net51 net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2763_ _1383_ _1087_ _0473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1714_ _0694_ _0753_ _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2694_ _0368_ _0378_ _0399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1645_ _0635_ _0667_ _0685_ _0686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1576_ _0610_ _0613_ _0614_ _0619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__2352__A2 _0030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2128_ _1093_ _1096_ _1177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_42_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2059_ _1034_ _1042_ _1101_ _1102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_26_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1615__A1 _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2811__I net60 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output53_I net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1606__A1 _1375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2031__A1 _1065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1909__A2 _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2582__A2 _0814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1430_ net27 _0095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xoutput91 net91 yB[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput80 net80 yA[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__2098__A1 net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2815_ net64 net81 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2746_ _0427_ _0454_ _0455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2022__A1 net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2677_ _0380_ _0381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1628_ _0580_ _0608_ _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1559_ net15 _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2316__A2 _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1827__A1 _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2600_ _0211_ _0297_ _0298_ _0299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2531_ _0175_ _0179_ _0223_ _0224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2307__A2 _0813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2462_ _0098_ _0099_ _0148_ _0151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_2393_ _0023_ _0075_ _0076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1413_ _1288_ _1299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_3_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1530__A3 _0225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2729_ _0372_ _0404_ _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_3_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2482__A1 net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2537__A2 _0229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1962_ _0996_ _0998_ _0999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__2225__A1 _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1893_ _0924_ _0927_ _0930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2514_ _0203_ _0206_ _0207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2445_ net16 net20 _0132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1525__I _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2376_ _1381_ _0004_ _0057_ _0058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_24_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2216__A1 _0225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2230_ _0567_ _0747_ _1286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2161_ _1198_ _1212_ _1213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__1497__A2 _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2092_ net28 _0781_ _1139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2446__A1 _1371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1945_ _0849_ _0980_ _0981_ _0891_ _0982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_9_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1876_ _0911_ _0912_ _0913_ _0818_ _0914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_2428_ _0056_ _0111_ _0112_ _0113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2359_ _1378_ _0005_ _0039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1488__A2 _0225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2685__A1 _0388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2437__A1 _0119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input15_I dba[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2814__I net63 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1660__A2 _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1479__A2 _0106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1730_ _0765_ _0769_ _0770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1661_ _0646_ _0648_ _0702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_7_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1592_ _1192_ _0633_ _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2213_ _1266_ _1229_ _1267_ _1268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input7_I dba[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2144_ _1110_ _1193_ _1194_ _1195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_26_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2075_ _1102_ _1106_ _1119_ _1120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_19_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1928_ _0834_ _0963_ _0964_ _0878_ _0965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_30_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1859_ _0887_ _0896_ _0897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_30_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2809__I net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1633__A2 _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2831_ net50 net97 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2762_ _0404_ _0469_ _0434_ _0470_ _0472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_8_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1713_ _0748_ _0752_ _0753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2693_ _0370_ _0377_ _0398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_6_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1644_ _0638_ _0666_ _0685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1575_ _0544_ _0546_ _0618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2127_ _1089_ _1156_ _1175_ _1176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2058_ _1037_ _1100_ _1101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1615__A2 _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2040__A2 _1081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1551__A1 _1375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output46_I net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1606__A2 _0526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2031__A2 _1069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput70 net70 yA[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput92 net92 yB[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__1542__A1 net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput81 net81 yA[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__2098__A2 net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2814_ net63 net80 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2745_ _0449_ _0453_ _0454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2022__A2 _0847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2676_ _0362_ _0379_ _0380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1627_ _0580_ _0608_ _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1558_ _1171_ _0535_ _0601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1489_ _0236_ _0531_ _0532_ _0461_ _0533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2822__I net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2013__A2 _1050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1827__A2 _0853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2530_ _0170_ _0174_ _0223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1763__A1 _0798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2461_ _0098_ _0099_ _0148_ _0149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_5_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1412_ net26 _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2392_ _0025_ _0073_ _0075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_3_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1530__A4 _0106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2728_ _0432_ _0433_ _0434_ _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__1754__A1 _0734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2659_ _0328_ _0333_ _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2817__I net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2482__A2 net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2537__A3 _0230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2170__B2 _1137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2170__A1 _1050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1961_ _0861_ _0859_ _0930_ _0997_ _0998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__2225__A2 net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1892_ _0929_ net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2513_ _0081_ _0091_ _0153_ _0205_ _0206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_2444_ _0115_ _0130_ _0131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2375_ _0000_ _0003_ _0057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2161__A1 _1198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1541__I _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2216__A2 _1199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1975__A1 _0943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1727__A1 net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2207__A2 _1261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1966__A1 _0995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1718__A1 _0712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2160_ _1204_ _1211_ _1212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2091_ net29 net2 _1137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_19_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1944_ _1084_ _0847_ _0893_ net17 _0981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_21_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1875_ _1386_ _0633_ _0692_ _1018_ _0913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1709__A1 net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2427_ _0058_ _0070_ _0112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2358_ _0026_ _0037_ _0038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_29_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2289_ _0535_ _0905_ _1350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2437__A2 _0122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1948__A1 net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2830__I net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2373__A1 _0049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output76_I net76 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1660_ net10 _0553_ _0701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1591_ _0632_ _0633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2116__A1 _0995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2212_ _1223_ _1228_ _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2143_ _1113_ _1118_ _1194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1875__B1 _0692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2074_ _1110_ _1113_ _1118_ _1119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_22_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1927_ _0872_ _0879_ _0964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1858_ _0890_ _0895_ _0896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1789_ _0471_ _0554_ _0828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2825__I net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2594__A1 _0266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2830_ net49 net96 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1624__A3 _0665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2761_ _0432_ _0433_ _0470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_12_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2692_ _0396_ net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1712_ _0750_ _0751_ _0752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_6_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1643_ _1192_ _0633_ _0631_ _0684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_6_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1574_ _0610_ _0615_ _0616_ _0617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2126_ _1091_ _1155_ _1175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XPHY_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_19_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2057_ _1041_ _1100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_35_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2576__A1 _0226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1551__A2 _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output39_I net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput60 net60 Y[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput71 net71 yA[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput93 net93 yB[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__1542__A2 _0584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput82 net82 yA[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_23_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2813_ net62 net79 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1809__I _0847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2744_ _0451_ _0452_ _0453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2675_ _0368_ _0378_ _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1626_ _0635_ _0667_ _0668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1557_ _0536_ _0597_ _0599_ _0566_ _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1488_ _1105_ _0225_ _0482_ _1051_ _0532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2109_ _1089_ _1156_ _1157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_14_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2797__A1 _1384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2549__A1 _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2721__A1 _0388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1763__A2 _0801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2460_ _0101_ _0147_ _0148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1411_ _1214_ _1246_ _1277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2391_ _0038_ _0072_ _0073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_36_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2779__A1 _1384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2727_ _0893_ _1087_ _0434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2658_ _0358_ _0359_ _0360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2589_ _0178_ _0280_ _0286_ _0234_ _0287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_1609_ _0641_ _0650_ _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_27_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2833__I net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1681__A1 _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1960_ _0924_ _0927_ _0997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1891_ _0860_ _0928_ _0929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__1984__A2 _0991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2512_ _0097_ _0093_ _0152_ _0205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_5_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2443_ _0123_ _0129_ _0130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2374_ _0046_ _0055_ _0056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_29_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1727__A2 _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2828__I net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1663__A1 _0095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1907__I net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2090_ _1064_ _1074_ _1135_ _1136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_19_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1943_ _1084_ _0892_ _0980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1406__A1 _1062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1874_ net10 _0691_ _0912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1709__A2 _0691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2426_ _0058_ _0070_ _0111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2648__I _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2357_ _0028_ _0036_ _0037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_29_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2288_ _1347_ _1291_ _1348_ _1349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_37_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1948__A2 _0984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2070__A1 _0214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2061__A1 _1053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1590_ net32 _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2211_ _1220_ _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_38_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2142_ _1113_ _1118_ _1193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1875__A1 _1386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1875__B2 _1018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2073_ _1114_ _1117_ _1118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1926_ net14 _0553_ _0963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1857_ _0888_ _0891_ _0894_ _0895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_1_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1788_ _0771_ _0825_ _0826_ _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_1_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2409_ _0092_ net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input20_I dbb[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1618__A1 _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2291__A1 _0225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2760_ _1199_ _1384_ _0469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2691_ _0355_ _0395_ _0396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1711_ _1018_ _0633_ _0692_ net8 _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1642_ _0681_ _0676_ _0682_ _0678_ _0683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_8_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1573_ _0613_ _0614_ _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1848__A1 _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2125_ _1174_ net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2056_ _1045_ _1078_ _1098_ _1099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_26_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2576__A2 _0230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1909_ net8 _0905_ _0946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_1_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2836__I net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2016__A1 _1048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput50 net50 Y[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput61 net61 Y[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput72 net72 yA[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput83 net83 yB[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput94 net94 yB[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1650__I net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2812_ net61 net78 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2743_ _0415_ _0414_ _0452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2674_ _0370_ _0377_ _0378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1625_ _0638_ _0666_ _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1556_ _1116_ _0598_ _0568_ _1062_ _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1487_ _1094_ _0471_ _0531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1560__I _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2108_ _1091_ _1155_ _1156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_42_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2039_ _1019_ _1080_ _1081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__2797__A2 _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2605__B _0304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2549__A2 net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output51_I net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2485__A1 _0170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1410_ _1256_ net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2390_ _0041_ _0071_ _0072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_36_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2779__A2 _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2726_ _1383_ _1199_ _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1555__I _0535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2657_ _0335_ _0337_ _0359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1608_ _0645_ _0649_ _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2588_ _0233_ _0235_ _0286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1539_ _0573_ _0581_ _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2467__A1 _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1465__I net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1681__A2 _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1890_ _0861_ _0924_ _0927_ _0928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__2630__A1 _0747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2511_ _0149_ _0202_ _0203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2442_ _0124_ _0127_ _0129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_38_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2373_ _0049_ _0054_ _0055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__2449__A1 _1380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2621__A1 _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2709_ _0382_ _0385_ _0415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__2688__A1 _0294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1663__A2 _0535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1942_ _0966_ _0977_ _0978_ _0979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_14_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1406__A2 _1192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1873_ _1029_ _0633_ _0911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2425_ _0104_ _0109_ _0110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2356_ _0032_ _0035_ _0036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2287_ _1285_ _1290_ _1348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1645__A2 _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2070__A2 _0813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1581__A1 _0519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2210_ _1206_ _1210_ _1211_ _1204_ _1265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2141_ _1120_ _1152_ _1190_ _1191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2072_ _1111_ _1115_ _1117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_19_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1925_ _0882_ _0960_ _0961_ _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1856_ net17 _0893_ _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1787_ _0773_ _0786_ _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2408_ _0081_ _0091_ _0092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2339_ _1341_ _0008_ _0017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input13_I dba[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1618__A2 _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2291__A2 net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1554__A1 _1094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output81_I net81 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2690_ _0390_ _0394_ _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_8_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1710_ _0690_ _0749_ _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1641_ _0677_ _0681_ _0682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1572_ _0613_ _0614_ _0615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input5_I dba[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1848__A2 _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2124_ _1164_ _1173_ _1174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_35_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2055_ _1047_ _1077_ _1098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_19_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1908_ net1 _0944_ _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1839_ _0775_ _0875_ _0876_ _0840_ _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__1784__A1 _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1536__A1 _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput51 net51 Y[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput40 net40 Y[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput73 net73 yA[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput62 net62 Y[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput84 net84 yB[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput95 net95 yB[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_36_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2811_ net60 net77 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2742_ _0411_ _0413_ _0451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2673_ _0371_ _0376_ _0377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1624_ _0651_ _0653_ _0665_ _0666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_1555_ _0535_ _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1486_ _0418_ _0512_ _0529_ _0530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2107_ _1097_ _1154_ _1155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2038_ _1021_ _1079_ _1080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_22_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2182__A1 net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output44_I net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1748__A1 _0758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2725_ _0906_ _1384_ _0432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2656_ _0321_ _0336_ _0358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1607_ _0646_ _0647_ _0648_ _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__2164__A1 _1134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2587_ _0271_ _0284_ _0285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1538_ _0572_ _0573_ _0574_ _0581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1469_ _0450_ _0503_ _0512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__2467__A2 _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2155__A1 _0214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2630__A2 _1383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2510_ _0199_ _0201_ _0202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_5_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2441_ _0125_ _0126_ _0127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_5_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2372_ _0050_ _0052_ _0054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__1391__I _1051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2621__A2 _0906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2385__A1 net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2708_ _0411_ _0413_ _0414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2137__A1 _1183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2639_ _0325_ _0339_ _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_28_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2128__A1 _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2300__A1 net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1941_ net26 _0781_ _0978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1872_ _0907_ _0909_ _0910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2367__A1 _1367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2424_ _0107_ _0108_ _0109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2355_ _0033_ _1352_ _0034_ _0035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2286_ _1282_ _1347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_37_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2530__A1 _0170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1869__B1 _0906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2597__A1 _0294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2349__A1 _1366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2140_ _1122_ _1151_ _1190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2071_ net12 _0746_ _1115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1924_ _0884_ _0897_ _0961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2588__A1 _0233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1855_ _0892_ _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_30_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1786_ _0773_ _0786_ _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2760__A1 _1199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2407_ _0084_ _0090_ _0091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_29_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2338_ _0016_ net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2269_ _1318_ _1328_ _1329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_38_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2579__A1 _0692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1554__A2 _0568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1857__A3 _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1490__A1 _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1640_ _0673_ _0620_ _0672_ _0681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_6_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1571_ _0560_ _0578_ _0614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_6_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2123_ _1169_ _1172_ _1173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_13_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2054_ _1093_ _1096_ _1097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_35_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1907_ net22 _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1838_ _0095_ _0603_ _0719_ _1288_ _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1769_ _0758_ _0787_ _0808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_25_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput52 net52 Y[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput41 net41 Y[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput63 net63 Y[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput74 net74 yA[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput85 net85 yB[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput96 net96 yB[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_36_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2810_ net59 net76 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2741_ _0447_ _0448_ _0449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2672_ _0373_ _0374_ _0376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__1394__I _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1623_ _0656_ _0664_ _0665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1554_ _1094_ _0568_ _0597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1485_ _0450_ _0503_ _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
.ends

