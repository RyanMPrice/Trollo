VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO BinMultiplier
  CLASS BLOCK ;
  FOREIGN BinMultiplier ;
  ORIGIN 0.000 0.000 ;
  SIZE 400.000 BY 200.000 ;
  PIN Y[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 8.400 196.000 8.960 200.000 ;
    END
  END Y[0]
  PIN Y[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 131.600 196.000 132.160 200.000 ;
    END
  END Y[10]
  PIN Y[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 143.920 196.000 144.480 200.000 ;
    END
  END Y[11]
  PIN Y[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 156.240 196.000 156.800 200.000 ;
    END
  END Y[12]
  PIN Y[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 168.560 196.000 169.120 200.000 ;
    END
  END Y[13]
  PIN Y[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 180.880 196.000 181.440 200.000 ;
    END
  END Y[14]
  PIN Y[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 193.200 196.000 193.760 200.000 ;
    END
  END Y[15]
  PIN Y[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 205.520 196.000 206.080 200.000 ;
    END
  END Y[16]
  PIN Y[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 217.840 196.000 218.400 200.000 ;
    END
  END Y[17]
  PIN Y[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 230.160 196.000 230.720 200.000 ;
    END
  END Y[18]
  PIN Y[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 242.480 196.000 243.040 200.000 ;
    END
  END Y[19]
  PIN Y[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 20.720 196.000 21.280 200.000 ;
    END
  END Y[1]
  PIN Y[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 254.800 196.000 255.360 200.000 ;
    END
  END Y[20]
  PIN Y[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 267.120 196.000 267.680 200.000 ;
    END
  END Y[21]
  PIN Y[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 279.440 196.000 280.000 200.000 ;
    END
  END Y[22]
  PIN Y[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 291.760 196.000 292.320 200.000 ;
    END
  END Y[23]
  PIN Y[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 304.080 196.000 304.640 200.000 ;
    END
  END Y[24]
  PIN Y[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 316.400 196.000 316.960 200.000 ;
    END
  END Y[25]
  PIN Y[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 328.720 196.000 329.280 200.000 ;
    END
  END Y[26]
  PIN Y[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 341.040 196.000 341.600 200.000 ;
    END
  END Y[27]
  PIN Y[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 353.360 196.000 353.920 200.000 ;
    END
  END Y[28]
  PIN Y[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 365.680 196.000 366.240 200.000 ;
    END
  END Y[29]
  PIN Y[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 33.040 196.000 33.600 200.000 ;
    END
  END Y[2]
  PIN Y[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 378.000 196.000 378.560 200.000 ;
    END
  END Y[30]
  PIN Y[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 390.320 196.000 390.880 200.000 ;
    END
  END Y[31]
  PIN Y[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 45.360 196.000 45.920 200.000 ;
    END
  END Y[3]
  PIN Y[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 57.680 196.000 58.240 200.000 ;
    END
  END Y[4]
  PIN Y[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 70.000 196.000 70.560 200.000 ;
    END
  END Y[5]
  PIN Y[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 82.320 196.000 82.880 200.000 ;
    END
  END Y[6]
  PIN Y[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 94.640 196.000 95.200 200.000 ;
    END
  END Y[7]
  PIN Y[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 106.960 196.000 107.520 200.000 ;
    END
  END Y[8]
  PIN Y[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 119.280 196.000 119.840 200.000 ;
    END
  END Y[9]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 13.440 0.000 14.000 4.000 ;
    END
  END clk
  PIN dba[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 56.000 0.000 56.560 4.000 ;
    END
  END dba[0]
  PIN dba[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 162.400 0.000 162.960 4.000 ;
    END
  END dba[10]
  PIN dba[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 173.040 0.000 173.600 4.000 ;
    END
  END dba[11]
  PIN dba[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 183.680 0.000 184.240 4.000 ;
    END
  END dba[12]
  PIN dba[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 194.320 0.000 194.880 4.000 ;
    END
  END dba[13]
  PIN dba[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 204.960 0.000 205.520 4.000 ;
    END
  END dba[14]
  PIN dba[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 215.600 0.000 216.160 4.000 ;
    END
  END dba[15]
  PIN dba[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 66.640 0.000 67.200 4.000 ;
    END
  END dba[1]
  PIN dba[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 77.280 0.000 77.840 4.000 ;
    END
  END dba[2]
  PIN dba[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 87.920 0.000 88.480 4.000 ;
    END
  END dba[3]
  PIN dba[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 98.560 0.000 99.120 4.000 ;
    END
  END dba[4]
  PIN dba[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 109.200 0.000 109.760 4.000 ;
    END
  END dba[5]
  PIN dba[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 119.840 0.000 120.400 4.000 ;
    END
  END dba[6]
  PIN dba[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 130.480 0.000 131.040 4.000 ;
    END
  END dba[7]
  PIN dba[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 141.120 0.000 141.680 4.000 ;
    END
  END dba[8]
  PIN dba[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 151.760 0.000 152.320 4.000 ;
    END
  END dba[9]
  PIN dbb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 226.240 0.000 226.800 4.000 ;
    END
  END dbb[0]
  PIN dbb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 332.640 0.000 333.200 4.000 ;
    END
  END dbb[10]
  PIN dbb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 343.280 0.000 343.840 4.000 ;
    END
  END dbb[11]
  PIN dbb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 353.920 0.000 354.480 4.000 ;
    END
  END dbb[12]
  PIN dbb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 364.560 0.000 365.120 4.000 ;
    END
  END dbb[13]
  PIN dbb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 375.200 0.000 375.760 4.000 ;
    END
  END dbb[14]
  PIN dbb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 385.840 0.000 386.400 4.000 ;
    END
  END dbb[15]
  PIN dbb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 236.880 0.000 237.440 4.000 ;
    END
  END dbb[1]
  PIN dbb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 247.520 0.000 248.080 4.000 ;
    END
  END dbb[2]
  PIN dbb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 258.160 0.000 258.720 4.000 ;
    END
  END dbb[3]
  PIN dbb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 268.800 0.000 269.360 4.000 ;
    END
  END dbb[4]
  PIN dbb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 279.440 0.000 280.000 4.000 ;
    END
  END dbb[5]
  PIN dbb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 290.080 0.000 290.640 4.000 ;
    END
  END dbb[6]
  PIN dbb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 300.720 0.000 301.280 4.000 ;
    END
  END dbb[7]
  PIN dbb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 311.360 0.000 311.920 4.000 ;
    END
  END dbb[8]
  PIN dbb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 322.000 0.000 322.560 4.000 ;
    END
  END dbb[9]
  PIN done
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 45.360 0.000 45.920 4.000 ;
    END
  END done
  PIN enable
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 34.720 0.000 35.280 4.000 ;
    END
  END enable
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 24.080 0.000 24.640 4.000 ;
    END
  END rst
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 54.220 15.380 55.820 184.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 150.820 15.380 152.420 184.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 247.420 15.380 249.020 184.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 344.020 15.380 345.620 184.540 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 102.520 15.380 104.120 184.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 199.120 15.380 200.720 184.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 295.720 15.380 297.320 184.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 392.320 15.380 393.920 184.540 ;
    END
  END vss
  PIN yA[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 7.280 400.000 7.840 ;
    END
  END yA[0]
  PIN yA[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 130.480 400.000 131.040 ;
    END
  END yA[10]
  PIN yA[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 142.800 400.000 143.360 ;
    END
  END yA[11]
  PIN yA[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 155.120 400.000 155.680 ;
    END
  END yA[12]
  PIN yA[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 167.440 400.000 168.000 ;
    END
  END yA[13]
  PIN yA[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 179.760 400.000 180.320 ;
    END
  END yA[14]
  PIN yA[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 192.080 400.000 192.640 ;
    END
  END yA[15]
  PIN yA[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 19.600 400.000 20.160 ;
    END
  END yA[1]
  PIN yA[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 31.920 400.000 32.480 ;
    END
  END yA[2]
  PIN yA[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 44.240 400.000 44.800 ;
    END
  END yA[3]
  PIN yA[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 56.560 400.000 57.120 ;
    END
  END yA[4]
  PIN yA[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 68.880 400.000 69.440 ;
    END
  END yA[5]
  PIN yA[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 81.200 400.000 81.760 ;
    END
  END yA[6]
  PIN yA[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 93.520 400.000 94.080 ;
    END
  END yA[7]
  PIN yA[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 105.840 400.000 106.400 ;
    END
  END yA[8]
  PIN yA[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 118.160 400.000 118.720 ;
    END
  END yA[9]
  PIN yB[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 7.280 4.000 7.840 ;
    END
  END yB[0]
  PIN yB[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 130.480 4.000 131.040 ;
    END
  END yB[10]
  PIN yB[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 142.800 4.000 143.360 ;
    END
  END yB[11]
  PIN yB[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 155.120 4.000 155.680 ;
    END
  END yB[12]
  PIN yB[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 167.440 4.000 168.000 ;
    END
  END yB[13]
  PIN yB[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 179.760 4.000 180.320 ;
    END
  END yB[14]
  PIN yB[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 192.080 4.000 192.640 ;
    END
  END yB[15]
  PIN yB[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 19.600 4.000 20.160 ;
    END
  END yB[1]
  PIN yB[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 31.920 4.000 32.480 ;
    END
  END yB[2]
  PIN yB[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 44.240 4.000 44.800 ;
    END
  END yB[3]
  PIN yB[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 56.560 4.000 57.120 ;
    END
  END yB[4]
  PIN yB[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 68.880 4.000 69.440 ;
    END
  END yB[5]
  PIN yB[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 81.200 4.000 81.760 ;
    END
  END yB[6]
  PIN yB[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 93.520 4.000 94.080 ;
    END
  END yB[7]
  PIN yB[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 105.840 4.000 106.400 ;
    END
  END yB[8]
  PIN yB[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 118.160 4.000 118.720 ;
    END
  END yB[9]
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 393.920 184.540 ;
      LAYER Metal2 ;
        RECT 6.860 195.700 8.100 196.420 ;
        RECT 9.260 195.700 20.420 196.420 ;
        RECT 21.580 195.700 32.740 196.420 ;
        RECT 33.900 195.700 45.060 196.420 ;
        RECT 46.220 195.700 57.380 196.420 ;
        RECT 58.540 195.700 69.700 196.420 ;
        RECT 70.860 195.700 82.020 196.420 ;
        RECT 83.180 195.700 94.340 196.420 ;
        RECT 95.500 195.700 106.660 196.420 ;
        RECT 107.820 195.700 118.980 196.420 ;
        RECT 120.140 195.700 131.300 196.420 ;
        RECT 132.460 195.700 143.620 196.420 ;
        RECT 144.780 195.700 155.940 196.420 ;
        RECT 157.100 195.700 168.260 196.420 ;
        RECT 169.420 195.700 180.580 196.420 ;
        RECT 181.740 195.700 192.900 196.420 ;
        RECT 194.060 195.700 205.220 196.420 ;
        RECT 206.380 195.700 217.540 196.420 ;
        RECT 218.700 195.700 229.860 196.420 ;
        RECT 231.020 195.700 242.180 196.420 ;
        RECT 243.340 195.700 254.500 196.420 ;
        RECT 255.660 195.700 266.820 196.420 ;
        RECT 267.980 195.700 279.140 196.420 ;
        RECT 280.300 195.700 291.460 196.420 ;
        RECT 292.620 195.700 303.780 196.420 ;
        RECT 304.940 195.700 316.100 196.420 ;
        RECT 317.260 195.700 328.420 196.420 ;
        RECT 329.580 195.700 340.740 196.420 ;
        RECT 341.900 195.700 353.060 196.420 ;
        RECT 354.220 195.700 365.380 196.420 ;
        RECT 366.540 195.700 377.700 196.420 ;
        RECT 378.860 195.700 390.020 196.420 ;
        RECT 391.180 195.700 395.780 196.420 ;
        RECT 6.860 4.300 395.780 195.700 ;
        RECT 6.860 3.500 13.140 4.300 ;
        RECT 14.300 3.500 23.780 4.300 ;
        RECT 24.940 3.500 34.420 4.300 ;
        RECT 35.580 3.500 45.060 4.300 ;
        RECT 46.220 3.500 55.700 4.300 ;
        RECT 56.860 3.500 66.340 4.300 ;
        RECT 67.500 3.500 76.980 4.300 ;
        RECT 78.140 3.500 87.620 4.300 ;
        RECT 88.780 3.500 98.260 4.300 ;
        RECT 99.420 3.500 108.900 4.300 ;
        RECT 110.060 3.500 119.540 4.300 ;
        RECT 120.700 3.500 130.180 4.300 ;
        RECT 131.340 3.500 140.820 4.300 ;
        RECT 141.980 3.500 151.460 4.300 ;
        RECT 152.620 3.500 162.100 4.300 ;
        RECT 163.260 3.500 172.740 4.300 ;
        RECT 173.900 3.500 183.380 4.300 ;
        RECT 184.540 3.500 194.020 4.300 ;
        RECT 195.180 3.500 204.660 4.300 ;
        RECT 205.820 3.500 215.300 4.300 ;
        RECT 216.460 3.500 225.940 4.300 ;
        RECT 227.100 3.500 236.580 4.300 ;
        RECT 237.740 3.500 247.220 4.300 ;
        RECT 248.380 3.500 257.860 4.300 ;
        RECT 259.020 3.500 268.500 4.300 ;
        RECT 269.660 3.500 279.140 4.300 ;
        RECT 280.300 3.500 289.780 4.300 ;
        RECT 290.940 3.500 300.420 4.300 ;
        RECT 301.580 3.500 311.060 4.300 ;
        RECT 312.220 3.500 321.700 4.300 ;
        RECT 322.860 3.500 332.340 4.300 ;
        RECT 333.500 3.500 342.980 4.300 ;
        RECT 344.140 3.500 353.620 4.300 ;
        RECT 354.780 3.500 364.260 4.300 ;
        RECT 365.420 3.500 374.900 4.300 ;
        RECT 376.060 3.500 385.540 4.300 ;
        RECT 386.700 3.500 395.780 4.300 ;
      LAYER Metal3 ;
        RECT 4.300 191.780 395.700 192.500 ;
        RECT 4.000 180.620 396.000 191.780 ;
        RECT 4.300 179.460 395.700 180.620 ;
        RECT 4.000 168.300 396.000 179.460 ;
        RECT 4.300 167.140 395.700 168.300 ;
        RECT 4.000 155.980 396.000 167.140 ;
        RECT 4.300 154.820 395.700 155.980 ;
        RECT 4.000 143.660 396.000 154.820 ;
        RECT 4.300 142.500 395.700 143.660 ;
        RECT 4.000 131.340 396.000 142.500 ;
        RECT 4.300 130.180 395.700 131.340 ;
        RECT 4.000 119.020 396.000 130.180 ;
        RECT 4.300 117.860 395.700 119.020 ;
        RECT 4.000 106.700 396.000 117.860 ;
        RECT 4.300 105.540 395.700 106.700 ;
        RECT 4.000 94.380 396.000 105.540 ;
        RECT 4.300 93.220 395.700 94.380 ;
        RECT 4.000 82.060 396.000 93.220 ;
        RECT 4.300 80.900 395.700 82.060 ;
        RECT 4.000 69.740 396.000 80.900 ;
        RECT 4.300 68.580 395.700 69.740 ;
        RECT 4.000 57.420 396.000 68.580 ;
        RECT 4.300 56.260 395.700 57.420 ;
        RECT 4.000 45.100 396.000 56.260 ;
        RECT 4.300 43.940 395.700 45.100 ;
        RECT 4.000 32.780 396.000 43.940 ;
        RECT 4.300 31.620 395.700 32.780 ;
        RECT 4.000 20.460 396.000 31.620 ;
        RECT 4.300 19.300 395.700 20.460 ;
        RECT 4.000 8.140 396.000 19.300 ;
        RECT 4.300 6.980 395.700 8.140 ;
        RECT 4.000 4.060 396.000 6.980 ;
      LAYER Metal4 ;
        RECT 75.740 18.570 102.220 175.750 ;
        RECT 104.420 18.570 150.520 175.750 ;
        RECT 152.720 18.570 198.820 175.750 ;
        RECT 201.020 18.570 247.120 175.750 ;
        RECT 249.320 18.570 295.420 175.750 ;
        RECT 297.620 18.570 343.720 175.750 ;
        RECT 345.920 18.570 390.180 175.750 ;
  END
END BinMultiplier
END LIBRARY

