magic
tech gf180mcuC
magscale 1 10
timestamp 1670260751
<< metal1 >>
rect 1344 36874 78624 36908
rect 1344 36822 10874 36874
rect 10926 36822 10978 36874
rect 11030 36822 11082 36874
rect 11134 36822 30194 36874
rect 30246 36822 30298 36874
rect 30350 36822 30402 36874
rect 30454 36822 49514 36874
rect 49566 36822 49618 36874
rect 49670 36822 49722 36874
rect 49774 36822 68834 36874
rect 68886 36822 68938 36874
rect 68990 36822 69042 36874
rect 69094 36822 78624 36874
rect 1344 36788 78624 36822
rect 33518 36594 33570 36606
rect 77982 36594 78034 36606
rect 2034 36542 2046 36594
rect 2098 36542 2110 36594
rect 4162 36542 4174 36594
rect 4226 36542 4238 36594
rect 6962 36542 6974 36594
rect 7026 36542 7038 36594
rect 9762 36542 9774 36594
rect 9826 36542 9838 36594
rect 11778 36542 11790 36594
rect 11842 36542 11854 36594
rect 14354 36542 14366 36594
rect 14418 36542 14430 36594
rect 19282 36542 19294 36594
rect 19346 36542 19358 36594
rect 21634 36542 21646 36594
rect 21698 36542 21710 36594
rect 23874 36542 23886 36594
rect 23938 36542 23950 36594
rect 26674 36542 26686 36594
rect 26738 36542 26750 36594
rect 29362 36542 29374 36594
rect 29426 36542 29438 36594
rect 31266 36542 31278 36594
rect 31330 36542 31342 36594
rect 34066 36542 34078 36594
rect 34130 36542 34142 36594
rect 37202 36542 37214 36594
rect 37266 36542 37278 36594
rect 41458 36542 41470 36594
rect 41522 36542 41534 36594
rect 46386 36542 46398 36594
rect 46450 36542 46462 36594
rect 48962 36542 48974 36594
rect 49026 36542 49038 36594
rect 50978 36542 50990 36594
rect 51042 36542 51054 36594
rect 54338 36542 54350 36594
rect 54402 36542 54414 36594
rect 56802 36542 56814 36594
rect 56866 36542 56878 36594
rect 58818 36542 58830 36594
rect 58882 36542 58894 36594
rect 61730 36542 61742 36594
rect 61794 36542 61806 36594
rect 64642 36542 64654 36594
rect 64706 36542 64718 36594
rect 66434 36542 66446 36594
rect 66498 36542 66510 36594
rect 68562 36542 68574 36594
rect 68626 36542 68638 36594
rect 70690 36542 70702 36594
rect 70754 36542 70766 36594
rect 74050 36542 74062 36594
rect 74114 36542 74126 36594
rect 76962 36542 76974 36594
rect 77026 36542 77038 36594
rect 33518 36530 33570 36542
rect 77982 36530 78034 36542
rect 13694 36482 13746 36494
rect 17726 36482 17778 36494
rect 3154 36430 3166 36482
rect 3218 36430 3230 36482
rect 4946 36430 4958 36482
rect 5010 36430 5022 36482
rect 8082 36430 8094 36482
rect 8146 36430 8158 36482
rect 10658 36430 10670 36482
rect 10722 36430 10734 36482
rect 12562 36430 12574 36482
rect 12626 36430 12638 36482
rect 15474 36430 15486 36482
rect 15538 36430 15550 36482
rect 17490 36430 17502 36482
rect 17554 36430 17566 36482
rect 13694 36418 13746 36430
rect 17726 36418 17778 36430
rect 17950 36482 18002 36494
rect 35646 36482 35698 36494
rect 20402 36430 20414 36482
rect 20466 36430 20478 36482
rect 22754 36430 22766 36482
rect 22818 36430 22830 36482
rect 24546 36430 24558 36482
rect 24610 36430 24622 36482
rect 27794 36430 27806 36482
rect 27858 36430 27870 36482
rect 30482 36430 30494 36482
rect 30546 36430 30558 36482
rect 32386 36430 32398 36482
rect 32450 36430 32462 36482
rect 35186 36430 35198 36482
rect 35250 36430 35262 36482
rect 17950 36418 18002 36430
rect 35646 36418 35698 36430
rect 35870 36482 35922 36494
rect 35870 36418 35922 36430
rect 36206 36482 36258 36494
rect 37426 36430 37438 36482
rect 37490 36430 37502 36482
rect 38658 36430 38670 36482
rect 38722 36430 38734 36482
rect 42578 36430 42590 36482
rect 42642 36430 42654 36482
rect 47506 36430 47518 36482
rect 47570 36430 47582 36482
rect 49858 36430 49870 36482
rect 49922 36430 49934 36482
rect 51874 36430 51886 36482
rect 51938 36430 51950 36482
rect 53666 36430 53678 36482
rect 53730 36430 53742 36482
rect 57698 36430 57710 36482
rect 57762 36430 57774 36482
rect 59826 36430 59838 36482
rect 59890 36430 59902 36482
rect 61282 36430 61294 36482
rect 61346 36430 61358 36482
rect 65762 36430 65774 36482
rect 65826 36430 65838 36482
rect 67554 36430 67566 36482
rect 67618 36430 67630 36482
rect 69458 36430 69470 36482
rect 69522 36430 69534 36482
rect 71362 36430 71374 36482
rect 71426 36430 71438 36482
rect 73378 36430 73390 36482
rect 73442 36430 73454 36482
rect 75394 36430 75406 36482
rect 75458 36430 75470 36482
rect 76290 36430 76302 36482
rect 76354 36430 76366 36482
rect 36206 36418 36258 36430
rect 16718 36370 16770 36382
rect 16718 36306 16770 36318
rect 18062 36370 18114 36382
rect 18062 36306 18114 36318
rect 25790 36370 25842 36382
rect 25790 36306 25842 36318
rect 28590 36370 28642 36382
rect 28590 36306 28642 36318
rect 36094 36370 36146 36382
rect 36094 36306 36146 36318
rect 39454 36370 39506 36382
rect 39454 36306 39506 36318
rect 43822 36370 43874 36382
rect 43822 36306 43874 36318
rect 44158 36370 44210 36382
rect 44158 36306 44210 36318
rect 52782 36370 52834 36382
rect 52782 36306 52834 36318
rect 62862 36370 62914 36382
rect 62862 36306 62914 36318
rect 63198 36370 63250 36382
rect 63198 36306 63250 36318
rect 72494 36370 72546 36382
rect 72494 36306 72546 36318
rect 5630 36258 5682 36270
rect 5630 36194 5682 36206
rect 6078 36258 6130 36270
rect 6078 36194 6130 36206
rect 8542 36258 8594 36270
rect 8542 36194 8594 36206
rect 16382 36258 16434 36270
rect 16382 36194 16434 36206
rect 18734 36258 18786 36270
rect 18734 36194 18786 36206
rect 25230 36258 25282 36270
rect 25230 36194 25282 36206
rect 25902 36258 25954 36270
rect 25902 36194 25954 36206
rect 26126 36258 26178 36270
rect 26126 36194 26178 36206
rect 43038 36258 43090 36270
rect 43038 36194 43090 36206
rect 45054 36258 45106 36270
rect 45054 36194 45106 36206
rect 45278 36258 45330 36270
rect 45278 36194 45330 36206
rect 45390 36258 45442 36270
rect 45390 36194 45442 36206
rect 45502 36258 45554 36270
rect 45502 36194 45554 36206
rect 47966 36258 48018 36270
rect 47966 36194 48018 36206
rect 53118 36258 53170 36270
rect 53118 36194 53170 36206
rect 60510 36258 60562 36270
rect 60510 36194 60562 36206
rect 63870 36258 63922 36270
rect 63870 36194 63922 36206
rect 72830 36258 72882 36270
rect 72830 36194 72882 36206
rect 75182 36258 75234 36270
rect 75182 36194 75234 36206
rect 1344 36090 78784 36124
rect 1344 36038 20534 36090
rect 20586 36038 20638 36090
rect 20690 36038 20742 36090
rect 20794 36038 39854 36090
rect 39906 36038 39958 36090
rect 40010 36038 40062 36090
rect 40114 36038 59174 36090
rect 59226 36038 59278 36090
rect 59330 36038 59382 36090
rect 59434 36038 78494 36090
rect 78546 36038 78598 36090
rect 78650 36038 78702 36090
rect 78754 36038 78784 36090
rect 1344 36004 78784 36038
rect 5294 35922 5346 35934
rect 5294 35858 5346 35870
rect 14366 35922 14418 35934
rect 14366 35858 14418 35870
rect 24894 35922 24946 35934
rect 31166 35922 31218 35934
rect 26786 35870 26798 35922
rect 26850 35870 26862 35922
rect 27458 35870 27470 35922
rect 27522 35870 27534 35922
rect 28466 35870 28478 35922
rect 28530 35870 28542 35922
rect 24894 35858 24946 35870
rect 31166 35858 31218 35870
rect 33966 35922 34018 35934
rect 33966 35858 34018 35870
rect 40574 35922 40626 35934
rect 40574 35858 40626 35870
rect 49758 35922 49810 35934
rect 49758 35858 49810 35870
rect 53342 35922 53394 35934
rect 53342 35858 53394 35870
rect 60062 35922 60114 35934
rect 60062 35858 60114 35870
rect 67454 35922 67506 35934
rect 67454 35858 67506 35870
rect 67902 35922 67954 35934
rect 67902 35858 67954 35870
rect 70478 35922 70530 35934
rect 70478 35858 70530 35870
rect 71710 35922 71762 35934
rect 71710 35858 71762 35870
rect 73278 35922 73330 35934
rect 73278 35858 73330 35870
rect 3614 35810 3666 35822
rect 1922 35758 1934 35810
rect 1986 35758 1998 35810
rect 3614 35746 3666 35758
rect 4510 35810 4562 35822
rect 4510 35746 4562 35758
rect 4846 35810 4898 35822
rect 4846 35746 4898 35758
rect 12014 35810 12066 35822
rect 12014 35746 12066 35758
rect 15038 35810 15090 35822
rect 34862 35810 34914 35822
rect 17826 35758 17838 35810
rect 17890 35758 17902 35810
rect 28578 35758 28590 35810
rect 28642 35758 28654 35810
rect 15038 35746 15090 35758
rect 34862 35746 34914 35758
rect 34974 35810 35026 35822
rect 42702 35810 42754 35822
rect 52110 35810 52162 35822
rect 36530 35758 36542 35810
rect 36594 35758 36606 35810
rect 38994 35758 39006 35810
rect 39058 35758 39070 35810
rect 43922 35758 43934 35810
rect 43986 35758 43998 35810
rect 34974 35746 35026 35758
rect 42702 35746 42754 35758
rect 52110 35746 52162 35758
rect 62974 35810 63026 35822
rect 62974 35746 63026 35758
rect 72270 35810 72322 35822
rect 72270 35746 72322 35758
rect 72606 35810 72658 35822
rect 72606 35746 72658 35758
rect 74398 35810 74450 35822
rect 76066 35758 76078 35810
rect 76130 35758 76142 35810
rect 77858 35758 77870 35810
rect 77922 35758 77934 35810
rect 74398 35746 74450 35758
rect 3950 35698 4002 35710
rect 3042 35646 3054 35698
rect 3106 35646 3118 35698
rect 3950 35634 4002 35646
rect 11006 35698 11058 35710
rect 11006 35634 11058 35646
rect 11454 35698 11506 35710
rect 11454 35634 11506 35646
rect 11902 35698 11954 35710
rect 11902 35634 11954 35646
rect 12238 35698 12290 35710
rect 12238 35634 12290 35646
rect 12686 35698 12738 35710
rect 12686 35634 12738 35646
rect 12910 35698 12962 35710
rect 22430 35698 22482 35710
rect 23998 35698 24050 35710
rect 13570 35646 13582 35698
rect 13634 35646 13646 35698
rect 16370 35646 16382 35698
rect 16434 35646 16446 35698
rect 18834 35646 18846 35698
rect 18898 35646 18910 35698
rect 19730 35646 19742 35698
rect 19794 35646 19806 35698
rect 19954 35646 19966 35698
rect 20018 35646 20030 35698
rect 21970 35646 21982 35698
rect 22034 35646 22046 35698
rect 23314 35646 23326 35698
rect 23378 35646 23390 35698
rect 12910 35634 12962 35646
rect 22430 35634 22482 35646
rect 23998 35634 24050 35646
rect 24558 35698 24610 35710
rect 24558 35634 24610 35646
rect 26462 35698 26514 35710
rect 29374 35698 29426 35710
rect 27346 35646 27358 35698
rect 27410 35646 27422 35698
rect 28466 35646 28478 35698
rect 28530 35646 28542 35698
rect 26462 35634 26514 35646
rect 29374 35634 29426 35646
rect 29598 35698 29650 35710
rect 31054 35698 31106 35710
rect 29810 35646 29822 35698
rect 29874 35646 29886 35698
rect 29598 35634 29650 35646
rect 31054 35634 31106 35646
rect 31390 35698 31442 35710
rect 32734 35698 32786 35710
rect 32386 35646 32398 35698
rect 32450 35646 32462 35698
rect 31390 35634 31442 35646
rect 32734 35634 32786 35646
rect 32846 35698 32898 35710
rect 32846 35634 32898 35646
rect 33630 35698 33682 35710
rect 33630 35634 33682 35646
rect 35086 35698 35138 35710
rect 45614 35698 45666 35710
rect 47854 35698 47906 35710
rect 51998 35698 52050 35710
rect 37650 35646 37662 35698
rect 37714 35646 37726 35698
rect 40114 35646 40126 35698
rect 40178 35646 40190 35698
rect 41794 35646 41806 35698
rect 41858 35646 41870 35698
rect 44930 35646 44942 35698
rect 44994 35646 45006 35698
rect 46050 35646 46062 35698
rect 46114 35646 46126 35698
rect 48066 35646 48078 35698
rect 48130 35646 48142 35698
rect 51426 35646 51438 35698
rect 51490 35646 51502 35698
rect 35086 35634 35138 35646
rect 45614 35634 45666 35646
rect 47854 35634 47906 35646
rect 51998 35634 52050 35646
rect 55358 35698 55410 35710
rect 55358 35634 55410 35646
rect 55918 35698 55970 35710
rect 55918 35634 55970 35646
rect 56030 35698 56082 35710
rect 56030 35634 56082 35646
rect 56142 35698 56194 35710
rect 56142 35634 56194 35646
rect 59166 35698 59218 35710
rect 59166 35634 59218 35646
rect 61406 35698 61458 35710
rect 64206 35698 64258 35710
rect 61842 35646 61854 35698
rect 61906 35646 61918 35698
rect 61406 35634 61458 35646
rect 64206 35634 64258 35646
rect 64430 35698 64482 35710
rect 64430 35634 64482 35646
rect 64766 35698 64818 35710
rect 66558 35698 66610 35710
rect 65650 35646 65662 35698
rect 65714 35646 65726 35698
rect 64766 35634 64818 35646
rect 66558 35634 66610 35646
rect 67118 35698 67170 35710
rect 67118 35634 67170 35646
rect 70814 35698 70866 35710
rect 74162 35646 74174 35698
rect 74226 35646 74238 35698
rect 74946 35646 74958 35698
rect 75010 35646 75022 35698
rect 76738 35646 76750 35698
rect 76802 35646 76814 35698
rect 70814 35634 70866 35646
rect 10446 35586 10498 35598
rect 16718 35586 16770 35598
rect 15138 35534 15150 35586
rect 15202 35534 15214 35586
rect 16034 35534 16046 35586
rect 16098 35534 16110 35586
rect 10446 35522 10498 35534
rect 16718 35522 16770 35534
rect 19518 35586 19570 35598
rect 26238 35586 26290 35598
rect 21522 35534 21534 35586
rect 21586 35534 21598 35586
rect 23090 35534 23102 35586
rect 23154 35534 23166 35586
rect 19518 35522 19570 35534
rect 26238 35522 26290 35534
rect 38110 35586 38162 35598
rect 48750 35586 48802 35598
rect 42018 35534 42030 35586
rect 42082 35534 42094 35586
rect 46498 35534 46510 35586
rect 46562 35534 46574 35586
rect 38110 35522 38162 35534
rect 48750 35522 48802 35534
rect 50542 35586 50594 35598
rect 50542 35522 50594 35534
rect 52558 35586 52610 35598
rect 57486 35586 57538 35598
rect 56578 35534 56590 35586
rect 56642 35534 56654 35586
rect 52558 35522 52610 35534
rect 57486 35522 57538 35534
rect 58046 35586 58098 35598
rect 58046 35522 58098 35534
rect 58942 35586 58994 35598
rect 58942 35522 58994 35534
rect 60510 35586 60562 35598
rect 60510 35522 60562 35534
rect 62302 35586 62354 35598
rect 64542 35586 64594 35598
rect 68350 35586 68402 35598
rect 62850 35534 62862 35586
rect 62914 35534 62926 35586
rect 65762 35534 65774 35586
rect 65826 35534 65838 35586
rect 62302 35522 62354 35534
rect 64542 35522 64594 35534
rect 68350 35522 68402 35534
rect 69022 35586 69074 35598
rect 69022 35522 69074 35534
rect 69694 35586 69746 35598
rect 69694 35522 69746 35534
rect 71262 35586 71314 35598
rect 71262 35522 71314 35534
rect 14814 35474 14866 35486
rect 49534 35474 49586 35486
rect 35522 35422 35534 35474
rect 35586 35422 35598 35474
rect 14814 35410 14866 35422
rect 49534 35410 49586 35422
rect 49870 35474 49922 35486
rect 49870 35410 49922 35422
rect 57710 35474 57762 35486
rect 57710 35410 57762 35422
rect 59390 35474 59442 35486
rect 59390 35410 59442 35422
rect 59614 35474 59666 35486
rect 59614 35410 59666 35422
rect 60622 35474 60674 35486
rect 60622 35410 60674 35422
rect 63198 35474 63250 35486
rect 63198 35410 63250 35422
rect 69582 35474 69634 35486
rect 69582 35410 69634 35422
rect 1344 35306 78624 35340
rect 1344 35254 10874 35306
rect 10926 35254 10978 35306
rect 11030 35254 11082 35306
rect 11134 35254 30194 35306
rect 30246 35254 30298 35306
rect 30350 35254 30402 35306
rect 30454 35254 49514 35306
rect 49566 35254 49618 35306
rect 49670 35254 49722 35306
rect 49774 35254 68834 35306
rect 68886 35254 68938 35306
rect 68990 35254 69042 35306
rect 69094 35254 78624 35306
rect 1344 35220 78624 35254
rect 15038 35138 15090 35150
rect 15038 35074 15090 35086
rect 19742 35138 19794 35150
rect 22654 35138 22706 35150
rect 20066 35086 20078 35138
rect 20130 35086 20142 35138
rect 19742 35074 19794 35086
rect 22654 35074 22706 35086
rect 22990 35138 23042 35150
rect 22990 35074 23042 35086
rect 26014 35138 26066 35150
rect 47182 35138 47234 35150
rect 32050 35086 32062 35138
rect 32114 35086 32126 35138
rect 26014 35074 26066 35086
rect 47182 35074 47234 35086
rect 48190 35138 48242 35150
rect 48190 35074 48242 35086
rect 48302 35138 48354 35150
rect 48302 35074 48354 35086
rect 48526 35138 48578 35150
rect 57362 35086 57374 35138
rect 57426 35135 57438 35138
rect 58146 35135 58158 35138
rect 57426 35089 58158 35135
rect 57426 35086 57438 35089
rect 58146 35086 58158 35089
rect 58210 35086 58222 35138
rect 59154 35086 59166 35138
rect 59218 35086 59230 35138
rect 64978 35086 64990 35138
rect 65042 35086 65054 35138
rect 48526 35074 48578 35086
rect 4398 35026 4450 35038
rect 2146 34974 2158 35026
rect 2210 34974 2222 35026
rect 4398 34962 4450 34974
rect 4846 35026 4898 35038
rect 12014 35026 12066 35038
rect 11666 34974 11678 35026
rect 11730 34974 11742 35026
rect 4846 34962 4898 34974
rect 12014 34962 12066 34974
rect 13918 35026 13970 35038
rect 13918 34962 13970 34974
rect 14142 35026 14194 35038
rect 14142 34962 14194 34974
rect 17278 35026 17330 35038
rect 17278 34962 17330 34974
rect 19518 35026 19570 35038
rect 19518 34962 19570 34974
rect 21870 35026 21922 35038
rect 21870 34962 21922 34974
rect 27470 35026 27522 35038
rect 27470 34962 27522 34974
rect 27918 35026 27970 35038
rect 44718 35026 44770 35038
rect 31378 34974 31390 35026
rect 31442 34974 31454 35026
rect 42578 34974 42590 35026
rect 42642 34974 42654 35026
rect 27918 34962 27970 34974
rect 44718 34962 44770 34974
rect 46174 35026 46226 35038
rect 57038 35026 57090 35038
rect 55682 34974 55694 35026
rect 55746 34974 55758 35026
rect 46174 34962 46226 34974
rect 57038 34962 57090 34974
rect 58158 35026 58210 35038
rect 66222 35026 66274 35038
rect 74062 35026 74114 35038
rect 62738 34974 62750 35026
rect 62802 34974 62814 35026
rect 69458 34974 69470 35026
rect 69522 34974 69534 35026
rect 76066 34974 76078 35026
rect 76130 34974 76142 35026
rect 58158 34962 58210 34974
rect 66222 34962 66274 34974
rect 74062 34962 74114 34974
rect 3950 34914 4002 34926
rect 14366 34914 14418 34926
rect 3042 34862 3054 34914
rect 3106 34862 3118 34914
rect 11330 34862 11342 34914
rect 11394 34862 11406 34914
rect 12674 34862 12686 34914
rect 12738 34862 12750 34914
rect 3950 34850 4002 34862
rect 14366 34850 14418 34862
rect 14590 34914 14642 34926
rect 14590 34850 14642 34862
rect 16382 34914 16434 34926
rect 18958 34914 19010 34926
rect 16818 34862 16830 34914
rect 16882 34862 16894 34914
rect 16382 34850 16434 34862
rect 18958 34850 19010 34862
rect 20526 34914 20578 34926
rect 20526 34850 20578 34862
rect 23550 34914 23602 34926
rect 23550 34850 23602 34862
rect 23886 34914 23938 34926
rect 23886 34850 23938 34862
rect 25342 34914 25394 34926
rect 25342 34850 25394 34862
rect 26574 34914 26626 34926
rect 28814 34914 28866 34926
rect 34750 34914 34802 34926
rect 35646 34914 35698 34926
rect 26786 34862 26798 34914
rect 26850 34862 26862 34914
rect 31266 34862 31278 34914
rect 31330 34862 31342 34914
rect 35186 34862 35198 34914
rect 35250 34862 35262 34914
rect 26574 34850 26626 34862
rect 28814 34850 28866 34862
rect 34750 34850 34802 34862
rect 35646 34850 35698 34862
rect 36542 34914 36594 34926
rect 40350 34914 40402 34926
rect 39778 34862 39790 34914
rect 39842 34862 39854 34914
rect 36542 34850 36594 34862
rect 40350 34850 40402 34862
rect 40462 34914 40514 34926
rect 40462 34850 40514 34862
rect 41358 34914 41410 34926
rect 49982 34914 50034 34926
rect 44034 34862 44046 34914
rect 44098 34862 44110 34914
rect 47170 34862 47182 34914
rect 47234 34862 47246 34914
rect 41358 34850 41410 34862
rect 49982 34850 50034 34862
rect 50878 34914 50930 34926
rect 56030 34914 56082 34926
rect 55234 34862 55246 34914
rect 55298 34862 55310 34914
rect 50878 34850 50930 34862
rect 56030 34850 56082 34862
rect 56590 34914 56642 34926
rect 56590 34850 56642 34862
rect 57262 34914 57314 34926
rect 57262 34850 57314 34862
rect 59054 34914 59106 34926
rect 65550 34914 65602 34926
rect 59714 34862 59726 34914
rect 59778 34862 59790 34914
rect 62514 34862 62526 34914
rect 62578 34862 62590 34914
rect 64978 34862 64990 34914
rect 65042 34862 65054 34914
rect 65314 34862 65326 34914
rect 65378 34862 65390 34914
rect 59054 34850 59106 34862
rect 65550 34850 65602 34862
rect 65998 34914 66050 34926
rect 65998 34850 66050 34862
rect 66670 34914 66722 34926
rect 66670 34850 66722 34862
rect 73278 34914 73330 34926
rect 74946 34862 74958 34914
rect 75010 34862 75022 34914
rect 73278 34850 73330 34862
rect 12910 34802 12962 34814
rect 12910 34738 12962 34750
rect 15822 34802 15874 34814
rect 15822 34738 15874 34750
rect 18622 34802 18674 34814
rect 18622 34738 18674 34750
rect 22430 34802 22482 34814
rect 22430 34738 22482 34750
rect 23662 34802 23714 34814
rect 23662 34738 23714 34750
rect 28478 34802 28530 34814
rect 28478 34738 28530 34750
rect 30494 34802 30546 34814
rect 30494 34738 30546 34750
rect 36206 34802 36258 34814
rect 36206 34738 36258 34750
rect 36654 34802 36706 34814
rect 36654 34738 36706 34750
rect 36766 34802 36818 34814
rect 36766 34738 36818 34750
rect 37550 34802 37602 34814
rect 46622 34802 46674 34814
rect 42802 34750 42814 34802
rect 42866 34750 42878 34802
rect 37550 34738 37602 34750
rect 46622 34738 46674 34750
rect 47518 34802 47570 34814
rect 47518 34738 47570 34750
rect 48638 34802 48690 34814
rect 48638 34738 48690 34750
rect 49758 34802 49810 34814
rect 49758 34738 49810 34750
rect 51774 34802 51826 34814
rect 51774 34738 51826 34750
rect 52110 34802 52162 34814
rect 52110 34738 52162 34750
rect 56814 34802 56866 34814
rect 56814 34738 56866 34750
rect 63198 34802 63250 34814
rect 63198 34738 63250 34750
rect 63982 34802 64034 34814
rect 63982 34738 64034 34750
rect 66446 34802 66498 34814
rect 72158 34802 72210 34814
rect 69682 34750 69694 34802
rect 69746 34750 69758 34802
rect 71362 34750 71374 34802
rect 71426 34750 71438 34802
rect 66446 34738 66498 34750
rect 72158 34738 72210 34750
rect 72270 34802 72322 34814
rect 72270 34738 72322 34750
rect 72494 34802 72546 34814
rect 72494 34738 72546 34750
rect 77310 34802 77362 34814
rect 77310 34738 77362 34750
rect 78094 34802 78146 34814
rect 78094 34738 78146 34750
rect 3614 34690 3666 34702
rect 3614 34626 3666 34638
rect 18174 34690 18226 34702
rect 18174 34626 18226 34638
rect 25006 34690 25058 34702
rect 25006 34626 25058 34638
rect 25678 34690 25730 34702
rect 25678 34626 25730 34638
rect 25902 34690 25954 34702
rect 25902 34626 25954 34638
rect 29598 34690 29650 34702
rect 29598 34626 29650 34638
rect 30270 34690 30322 34702
rect 30270 34626 30322 34638
rect 30382 34690 30434 34702
rect 30382 34626 30434 34638
rect 32622 34690 32674 34702
rect 32622 34626 32674 34638
rect 37662 34690 37714 34702
rect 37662 34626 37714 34638
rect 37774 34690 37826 34702
rect 37774 34626 37826 34638
rect 41470 34690 41522 34702
rect 41470 34626 41522 34638
rect 41694 34690 41746 34702
rect 41694 34626 41746 34638
rect 45390 34690 45442 34702
rect 45390 34626 45442 34638
rect 49198 34690 49250 34702
rect 51214 34690 51266 34702
rect 50306 34638 50318 34690
rect 50370 34638 50382 34690
rect 49198 34626 49250 34638
rect 51214 34626 51266 34638
rect 57598 34690 57650 34702
rect 57598 34626 57650 34638
rect 61294 34690 61346 34702
rect 61294 34626 61346 34638
rect 64094 34690 64146 34702
rect 64094 34626 64146 34638
rect 64766 34690 64818 34702
rect 64766 34626 64818 34638
rect 67118 34690 67170 34702
rect 73614 34690 73666 34702
rect 71250 34638 71262 34690
rect 71314 34638 71326 34690
rect 67118 34626 67170 34638
rect 73614 34626 73666 34638
rect 77646 34690 77698 34702
rect 77646 34626 77698 34638
rect 1344 34522 78784 34556
rect 1344 34470 20534 34522
rect 20586 34470 20638 34522
rect 20690 34470 20742 34522
rect 20794 34470 39854 34522
rect 39906 34470 39958 34522
rect 40010 34470 40062 34522
rect 40114 34470 59174 34522
rect 59226 34470 59278 34522
rect 59330 34470 59382 34522
rect 59434 34470 78494 34522
rect 78546 34470 78598 34522
rect 78650 34470 78702 34522
rect 78754 34470 78784 34522
rect 1344 34436 78784 34470
rect 12350 34354 12402 34366
rect 12350 34290 12402 34302
rect 15598 34354 15650 34366
rect 15598 34290 15650 34302
rect 16494 34354 16546 34366
rect 16494 34290 16546 34302
rect 17838 34354 17890 34366
rect 17838 34290 17890 34302
rect 18622 34354 18674 34366
rect 18622 34290 18674 34302
rect 18846 34354 18898 34366
rect 18846 34290 18898 34302
rect 26238 34354 26290 34366
rect 26238 34290 26290 34302
rect 27470 34354 27522 34366
rect 27470 34290 27522 34302
rect 30718 34354 30770 34366
rect 30718 34290 30770 34302
rect 31502 34354 31554 34366
rect 31502 34290 31554 34302
rect 33854 34354 33906 34366
rect 33854 34290 33906 34302
rect 37438 34354 37490 34366
rect 37438 34290 37490 34302
rect 39790 34354 39842 34366
rect 39790 34290 39842 34302
rect 40462 34354 40514 34366
rect 40462 34290 40514 34302
rect 40686 34354 40738 34366
rect 40686 34290 40738 34302
rect 42478 34354 42530 34366
rect 58270 34354 58322 34366
rect 43474 34302 43486 34354
rect 43538 34302 43550 34354
rect 42478 34290 42530 34302
rect 58270 34290 58322 34302
rect 59726 34354 59778 34366
rect 59726 34290 59778 34302
rect 62750 34354 62802 34366
rect 62750 34290 62802 34302
rect 65774 34354 65826 34366
rect 65774 34290 65826 34302
rect 70142 34354 70194 34366
rect 70142 34290 70194 34302
rect 72382 34354 72434 34366
rect 72382 34290 72434 34302
rect 73614 34354 73666 34366
rect 73614 34290 73666 34302
rect 8990 34242 9042 34254
rect 8990 34178 9042 34190
rect 13470 34242 13522 34254
rect 13470 34178 13522 34190
rect 13806 34242 13858 34254
rect 13806 34178 13858 34190
rect 14590 34242 14642 34254
rect 14590 34178 14642 34190
rect 16942 34242 16994 34254
rect 16942 34178 16994 34190
rect 17726 34242 17778 34254
rect 17726 34178 17778 34190
rect 17950 34242 18002 34254
rect 17950 34178 18002 34190
rect 21982 34242 22034 34254
rect 21982 34178 22034 34190
rect 24894 34242 24946 34254
rect 24894 34178 24946 34190
rect 26014 34242 26066 34254
rect 26014 34178 26066 34190
rect 27134 34242 27186 34254
rect 27134 34178 27186 34190
rect 27246 34242 27298 34254
rect 27246 34178 27298 34190
rect 31278 34242 31330 34254
rect 39454 34242 39506 34254
rect 35746 34190 35758 34242
rect 35810 34190 35822 34242
rect 31278 34178 31330 34190
rect 39454 34178 39506 34190
rect 40350 34242 40402 34254
rect 40350 34178 40402 34190
rect 43934 34242 43986 34254
rect 43934 34178 43986 34190
rect 51550 34242 51602 34254
rect 51550 34178 51602 34190
rect 51774 34242 51826 34254
rect 51774 34178 51826 34190
rect 52446 34242 52498 34254
rect 52446 34178 52498 34190
rect 52558 34242 52610 34254
rect 52558 34178 52610 34190
rect 53902 34242 53954 34254
rect 53902 34178 53954 34190
rect 55134 34242 55186 34254
rect 55134 34178 55186 34190
rect 59390 34242 59442 34254
rect 59390 34178 59442 34190
rect 59502 34242 59554 34254
rect 59502 34178 59554 34190
rect 60174 34242 60226 34254
rect 60174 34178 60226 34190
rect 62974 34242 63026 34254
rect 62974 34178 63026 34190
rect 65662 34242 65714 34254
rect 65662 34178 65714 34190
rect 71150 34242 71202 34254
rect 71150 34178 71202 34190
rect 74062 34242 74114 34254
rect 74062 34178 74114 34190
rect 74398 34242 74450 34254
rect 74398 34178 74450 34190
rect 76750 34242 76802 34254
rect 76750 34178 76802 34190
rect 77086 34242 77138 34254
rect 77086 34178 77138 34190
rect 77646 34242 77698 34254
rect 77646 34178 77698 34190
rect 13022 34130 13074 34142
rect 3042 34078 3054 34130
rect 3106 34078 3118 34130
rect 7186 34078 7198 34130
rect 7250 34078 7262 34130
rect 8194 34078 8206 34130
rect 8258 34078 8270 34130
rect 13022 34066 13074 34078
rect 13246 34130 13298 34142
rect 13246 34066 13298 34078
rect 13694 34130 13746 34142
rect 13694 34066 13746 34078
rect 18958 34130 19010 34142
rect 23886 34130 23938 34142
rect 20066 34078 20078 34130
rect 20130 34078 20142 34130
rect 21186 34078 21198 34130
rect 21250 34078 21262 34130
rect 23314 34078 23326 34130
rect 23378 34078 23390 34130
rect 18958 34066 19010 34078
rect 23886 34066 23938 34078
rect 26238 34130 26290 34142
rect 26238 34066 26290 34078
rect 26462 34130 26514 34142
rect 26462 34066 26514 34078
rect 32846 34130 32898 34142
rect 32846 34066 32898 34078
rect 33742 34130 33794 34142
rect 33742 34066 33794 34078
rect 33966 34130 34018 34142
rect 35422 34130 35474 34142
rect 43598 34130 43650 34142
rect 51886 34130 51938 34142
rect 34290 34078 34302 34130
rect 34354 34078 34366 34130
rect 43138 34078 43150 34130
rect 43202 34078 43214 34130
rect 50642 34078 50654 34130
rect 50706 34078 50718 34130
rect 33966 34066 34018 34078
rect 35422 34066 35474 34078
rect 43598 34066 43650 34078
rect 51886 34066 51938 34078
rect 52782 34130 52834 34142
rect 52782 34066 52834 34078
rect 53790 34130 53842 34142
rect 53790 34066 53842 34078
rect 57710 34130 57762 34142
rect 57710 34066 57762 34078
rect 57934 34130 57986 34142
rect 57934 34066 57986 34078
rect 58158 34130 58210 34142
rect 58158 34066 58210 34078
rect 58382 34130 58434 34142
rect 58382 34066 58434 34078
rect 60286 34130 60338 34142
rect 60286 34066 60338 34078
rect 60510 34130 60562 34142
rect 60510 34066 60562 34078
rect 60622 34130 60674 34142
rect 60622 34066 60674 34078
rect 63086 34130 63138 34142
rect 70254 34130 70306 34142
rect 77982 34130 78034 34142
rect 65986 34078 65998 34130
rect 66050 34078 66062 34130
rect 70914 34078 70926 34130
rect 70978 34078 70990 34130
rect 74946 34078 74958 34130
rect 75010 34078 75022 34130
rect 63086 34066 63138 34078
rect 70254 34066 70306 34078
rect 77982 34066 78034 34078
rect 9662 34018 9714 34030
rect 15150 34018 15202 34030
rect 24334 34018 24386 34030
rect 1922 33966 1934 34018
rect 1986 33966 1998 34018
rect 6738 33966 6750 34018
rect 6802 33966 6814 34018
rect 14690 33966 14702 34018
rect 14754 33966 14766 34018
rect 20178 33966 20190 34018
rect 20242 33966 20254 34018
rect 22978 33966 22990 34018
rect 23042 33966 23054 34018
rect 9662 33954 9714 33966
rect 15150 33954 15202 33966
rect 24334 33954 24386 33966
rect 35198 34018 35250 34030
rect 51102 34018 51154 34030
rect 37538 33966 37550 34018
rect 37602 33966 37614 34018
rect 42578 33966 42590 34018
rect 42642 33966 42654 34018
rect 50306 33966 50318 34018
rect 50370 33966 50382 34018
rect 35198 33954 35250 33966
rect 51102 33954 51154 33966
rect 53118 34018 53170 34030
rect 57486 34018 57538 34030
rect 55234 33966 55246 34018
rect 55298 33966 55310 34018
rect 53118 33954 53170 33966
rect 57486 33954 57538 33966
rect 71822 34018 71874 34030
rect 76066 33966 76078 34018
rect 76130 33966 76142 34018
rect 71822 33954 71874 33966
rect 14366 33906 14418 33918
rect 14366 33842 14418 33854
rect 31614 33906 31666 33918
rect 31614 33842 31666 33854
rect 37214 33906 37266 33918
rect 37214 33842 37266 33854
rect 42254 33906 42306 33918
rect 42254 33842 42306 33854
rect 43486 33906 43538 33918
rect 43486 33842 43538 33854
rect 53902 33906 53954 33918
rect 53902 33842 53954 33854
rect 54910 33906 54962 33918
rect 54910 33842 54962 33854
rect 70142 33906 70194 33918
rect 70142 33842 70194 33854
rect 1344 33738 78624 33772
rect 1344 33686 10874 33738
rect 10926 33686 10978 33738
rect 11030 33686 11082 33738
rect 11134 33686 30194 33738
rect 30246 33686 30298 33738
rect 30350 33686 30402 33738
rect 30454 33686 49514 33738
rect 49566 33686 49618 33738
rect 49670 33686 49722 33738
rect 49774 33686 68834 33738
rect 68886 33686 68938 33738
rect 68990 33686 69042 33738
rect 69094 33686 78624 33738
rect 1344 33652 78624 33686
rect 13806 33570 13858 33582
rect 13806 33506 13858 33518
rect 23550 33570 23602 33582
rect 42814 33570 42866 33582
rect 23874 33518 23886 33570
rect 23938 33518 23950 33570
rect 30594 33518 30606 33570
rect 30658 33518 30670 33570
rect 23550 33506 23602 33518
rect 42814 33506 42866 33518
rect 61518 33570 61570 33582
rect 61518 33506 61570 33518
rect 63198 33570 63250 33582
rect 63198 33506 63250 33518
rect 65102 33570 65154 33582
rect 65102 33506 65154 33518
rect 72270 33570 72322 33582
rect 73938 33518 73950 33570
rect 74002 33567 74014 33570
rect 74386 33567 74398 33570
rect 74002 33521 74398 33567
rect 74002 33518 74014 33521
rect 74386 33518 74398 33521
rect 74450 33518 74462 33570
rect 72270 33506 72322 33518
rect 3614 33458 3666 33470
rect 3614 33394 3666 33406
rect 6750 33458 6802 33470
rect 6750 33394 6802 33406
rect 8766 33458 8818 33470
rect 8766 33394 8818 33406
rect 9774 33458 9826 33470
rect 9774 33394 9826 33406
rect 14366 33458 14418 33470
rect 14366 33394 14418 33406
rect 17278 33458 17330 33470
rect 17278 33394 17330 33406
rect 21982 33458 22034 33470
rect 21982 33394 22034 33406
rect 22430 33458 22482 33470
rect 22430 33394 22482 33406
rect 22766 33458 22818 33470
rect 22766 33394 22818 33406
rect 23326 33458 23378 33470
rect 23326 33394 23378 33406
rect 28366 33458 28418 33470
rect 32062 33458 32114 33470
rect 42590 33458 42642 33470
rect 47294 33458 47346 33470
rect 29922 33406 29934 33458
rect 29986 33406 29998 33458
rect 34962 33406 34974 33458
rect 35026 33406 35038 33458
rect 37874 33406 37886 33458
rect 37938 33406 37950 33458
rect 40114 33406 40126 33458
rect 40178 33406 40190 33458
rect 43922 33406 43934 33458
rect 43986 33406 43998 33458
rect 28366 33394 28418 33406
rect 32062 33394 32114 33406
rect 42590 33394 42642 33406
rect 47294 33394 47346 33406
rect 47742 33458 47794 33470
rect 55694 33458 55746 33470
rect 49298 33406 49310 33458
rect 49362 33406 49374 33458
rect 53778 33406 53790 33458
rect 53842 33406 53854 33458
rect 47742 33394 47794 33406
rect 55694 33394 55746 33406
rect 71150 33458 71202 33470
rect 71150 33394 71202 33406
rect 73166 33458 73218 33470
rect 73166 33394 73218 33406
rect 74398 33458 74450 33470
rect 74398 33394 74450 33406
rect 75630 33458 75682 33470
rect 75630 33394 75682 33406
rect 3166 33346 3218 33358
rect 9662 33346 9714 33358
rect 8194 33294 8206 33346
rect 8258 33294 8270 33346
rect 3166 33282 3218 33294
rect 9662 33282 9714 33294
rect 10334 33346 10386 33358
rect 12686 33346 12738 33358
rect 12002 33294 12014 33346
rect 12066 33294 12078 33346
rect 10334 33282 10386 33294
rect 12686 33282 12738 33294
rect 12910 33346 12962 33358
rect 12910 33282 12962 33294
rect 17950 33346 18002 33358
rect 20414 33346 20466 33358
rect 18162 33294 18174 33346
rect 18226 33294 18238 33346
rect 19730 33294 19742 33346
rect 19794 33294 19806 33346
rect 17950 33282 18002 33294
rect 20414 33282 20466 33294
rect 28254 33346 28306 33358
rect 28254 33282 28306 33294
rect 28926 33346 28978 33358
rect 33518 33346 33570 33358
rect 48190 33346 48242 33358
rect 49870 33346 49922 33358
rect 50766 33346 50818 33358
rect 29810 33294 29822 33346
rect 29874 33294 29886 33346
rect 32834 33294 32846 33346
rect 32898 33294 32910 33346
rect 34178 33294 34190 33346
rect 34242 33294 34254 33346
rect 37986 33294 37998 33346
rect 38050 33294 38062 33346
rect 39330 33294 39342 33346
rect 39394 33294 39406 33346
rect 43138 33294 43150 33346
rect 43202 33294 43214 33346
rect 44258 33294 44270 33346
rect 44322 33294 44334 33346
rect 48402 33294 48414 33346
rect 48466 33294 48478 33346
rect 49634 33294 49646 33346
rect 49698 33294 49710 33346
rect 50418 33294 50430 33346
rect 50482 33294 50494 33346
rect 28926 33282 28978 33294
rect 33518 33282 33570 33294
rect 48190 33282 48242 33294
rect 49870 33282 49922 33294
rect 50766 33282 50818 33294
rect 50990 33346 51042 33358
rect 54574 33346 54626 33358
rect 56590 33346 56642 33358
rect 54114 33294 54126 33346
rect 54178 33294 54190 33346
rect 56130 33294 56142 33346
rect 56194 33294 56206 33346
rect 50990 33282 51042 33294
rect 54574 33282 54626 33294
rect 56590 33282 56642 33294
rect 57150 33346 57202 33358
rect 57150 33282 57202 33294
rect 57710 33346 57762 33358
rect 57710 33282 57762 33294
rect 57822 33346 57874 33358
rect 57822 33282 57874 33294
rect 64206 33346 64258 33358
rect 64206 33282 64258 33294
rect 65438 33346 65490 33358
rect 67118 33346 67170 33358
rect 66546 33294 66558 33346
rect 66610 33294 66622 33346
rect 65438 33282 65490 33294
rect 67118 33282 67170 33294
rect 70254 33346 70306 33358
rect 71934 33346 71986 33358
rect 70578 33294 70590 33346
rect 70642 33294 70654 33346
rect 70254 33282 70306 33294
rect 71934 33282 71986 33294
rect 73950 33346 74002 33358
rect 75058 33294 75070 33346
rect 75122 33294 75134 33346
rect 76402 33294 76414 33346
rect 76466 33294 76478 33346
rect 77522 33294 77534 33346
rect 77586 33294 77598 33346
rect 73950 33282 74002 33294
rect 13694 33234 13746 33246
rect 7186 33182 7198 33234
rect 7250 33182 7262 33234
rect 13694 33170 13746 33182
rect 13806 33234 13858 33246
rect 13806 33170 13858 33182
rect 18846 33234 18898 33246
rect 18846 33170 18898 33182
rect 44718 33234 44770 33246
rect 44718 33170 44770 33182
rect 45502 33234 45554 33246
rect 45502 33170 45554 33182
rect 45614 33234 45666 33246
rect 45614 33170 45666 33182
rect 45838 33234 45890 33246
rect 45838 33170 45890 33182
rect 51774 33234 51826 33246
rect 51774 33170 51826 33182
rect 60510 33234 60562 33246
rect 60510 33170 60562 33182
rect 61630 33234 61682 33246
rect 61630 33170 61682 33182
rect 62526 33234 62578 33246
rect 62526 33170 62578 33182
rect 63086 33234 63138 33246
rect 63086 33170 63138 33182
rect 63870 33234 63922 33246
rect 63870 33170 63922 33182
rect 63982 33234 64034 33246
rect 63982 33170 64034 33182
rect 65662 33234 65714 33246
rect 65662 33170 65714 33182
rect 67230 33234 67282 33246
rect 67230 33170 67282 33182
rect 71710 33234 71762 33246
rect 71710 33170 71762 33182
rect 2830 33122 2882 33134
rect 2830 33058 2882 33070
rect 9438 33122 9490 33134
rect 9438 33058 9490 33070
rect 9886 33122 9938 33134
rect 9886 33058 9938 33070
rect 19966 33122 20018 33134
rect 19966 33058 20018 33070
rect 28478 33122 28530 33134
rect 28478 33058 28530 33070
rect 36878 33122 36930 33134
rect 36878 33058 36930 33070
rect 51438 33122 51490 33134
rect 51438 33058 51490 33070
rect 51662 33122 51714 33134
rect 51662 33058 51714 33070
rect 52334 33122 52386 33134
rect 52334 33058 52386 33070
rect 52782 33122 52834 33134
rect 52782 33058 52834 33070
rect 57598 33122 57650 33134
rect 57598 33058 57650 33070
rect 59166 33122 59218 33134
rect 59166 33058 59218 33070
rect 60622 33122 60674 33134
rect 60622 33058 60674 33070
rect 61518 33122 61570 33134
rect 61518 33058 61570 33070
rect 74846 33122 74898 33134
rect 74846 33058 74898 33070
rect 76190 33122 76242 33134
rect 76190 33058 76242 33070
rect 77310 33122 77362 33134
rect 77310 33058 77362 33070
rect 78094 33122 78146 33134
rect 78094 33058 78146 33070
rect 1344 32954 78784 32988
rect 1344 32902 20534 32954
rect 20586 32902 20638 32954
rect 20690 32902 20742 32954
rect 20794 32902 39854 32954
rect 39906 32902 39958 32954
rect 40010 32902 40062 32954
rect 40114 32902 59174 32954
rect 59226 32902 59278 32954
rect 59330 32902 59382 32954
rect 59434 32902 78494 32954
rect 78546 32902 78598 32954
rect 78650 32902 78702 32954
rect 78754 32902 78784 32954
rect 1344 32868 78784 32902
rect 3614 32786 3666 32798
rect 3614 32722 3666 32734
rect 7422 32786 7474 32798
rect 7422 32722 7474 32734
rect 7646 32786 7698 32798
rect 7646 32722 7698 32734
rect 8206 32786 8258 32798
rect 8206 32722 8258 32734
rect 8318 32786 8370 32798
rect 8318 32722 8370 32734
rect 8990 32786 9042 32798
rect 8990 32722 9042 32734
rect 13134 32786 13186 32798
rect 13134 32722 13186 32734
rect 17614 32786 17666 32798
rect 17614 32722 17666 32734
rect 17838 32786 17890 32798
rect 38558 32786 38610 32798
rect 29474 32734 29486 32786
rect 29538 32734 29550 32786
rect 34178 32734 34190 32786
rect 34242 32734 34254 32786
rect 17838 32722 17890 32734
rect 38558 32722 38610 32734
rect 38670 32786 38722 32798
rect 38670 32722 38722 32734
rect 39230 32786 39282 32798
rect 39230 32722 39282 32734
rect 42366 32786 42418 32798
rect 49870 32786 49922 32798
rect 48066 32734 48078 32786
rect 48130 32734 48142 32786
rect 42366 32722 42418 32734
rect 49870 32722 49922 32734
rect 50654 32786 50706 32798
rect 50654 32722 50706 32734
rect 56030 32786 56082 32798
rect 56030 32722 56082 32734
rect 57934 32786 57986 32798
rect 57934 32722 57986 32734
rect 58494 32786 58546 32798
rect 58494 32722 58546 32734
rect 63534 32786 63586 32798
rect 63534 32722 63586 32734
rect 67230 32786 67282 32798
rect 67230 32722 67282 32734
rect 69582 32786 69634 32798
rect 69582 32722 69634 32734
rect 74286 32786 74338 32798
rect 74286 32722 74338 32734
rect 2830 32674 2882 32686
rect 2830 32610 2882 32622
rect 3166 32674 3218 32686
rect 3166 32610 3218 32622
rect 7310 32674 7362 32686
rect 7310 32610 7362 32622
rect 8094 32674 8146 32686
rect 8094 32610 8146 32622
rect 12798 32674 12850 32686
rect 12798 32610 12850 32622
rect 14926 32674 14978 32686
rect 14926 32610 14978 32622
rect 17950 32674 18002 32686
rect 17950 32610 18002 32622
rect 19742 32674 19794 32686
rect 19742 32610 19794 32622
rect 22654 32674 22706 32686
rect 22654 32610 22706 32622
rect 24894 32674 24946 32686
rect 24894 32610 24946 32622
rect 33630 32674 33682 32686
rect 49758 32674 49810 32686
rect 46610 32622 46622 32674
rect 46674 32622 46686 32674
rect 33630 32610 33682 32622
rect 49758 32610 49810 32622
rect 50094 32674 50146 32686
rect 50094 32610 50146 32622
rect 52222 32674 52274 32686
rect 52222 32610 52274 32622
rect 55918 32674 55970 32686
rect 55918 32610 55970 32622
rect 57486 32674 57538 32686
rect 57486 32610 57538 32622
rect 58718 32674 58770 32686
rect 58718 32610 58770 32622
rect 58830 32674 58882 32686
rect 58830 32610 58882 32622
rect 59278 32674 59330 32686
rect 59278 32610 59330 32622
rect 60286 32674 60338 32686
rect 60286 32610 60338 32622
rect 66446 32674 66498 32686
rect 66446 32610 66498 32622
rect 67454 32674 67506 32686
rect 67454 32610 67506 32622
rect 70478 32674 70530 32686
rect 70478 32610 70530 32622
rect 74734 32674 74786 32686
rect 74734 32610 74786 32622
rect 76526 32674 76578 32686
rect 76526 32610 76578 32622
rect 77198 32674 77250 32686
rect 77198 32610 77250 32622
rect 77534 32674 77586 32686
rect 77534 32610 77586 32622
rect 77982 32674 78034 32686
rect 77982 32610 78034 32622
rect 13022 32562 13074 32574
rect 13022 32498 13074 32510
rect 13246 32562 13298 32574
rect 18846 32562 18898 32574
rect 28926 32562 28978 32574
rect 14018 32510 14030 32562
rect 14082 32510 14094 32562
rect 19058 32510 19070 32562
rect 19122 32510 19134 32562
rect 22418 32510 22430 32562
rect 22482 32510 22494 32562
rect 24434 32510 24446 32562
rect 24498 32510 24510 32562
rect 27458 32510 27470 32562
rect 27522 32510 27534 32562
rect 13246 32498 13298 32510
rect 18846 32498 18898 32510
rect 28926 32498 28978 32510
rect 31166 32562 31218 32574
rect 31166 32498 31218 32510
rect 31502 32562 31554 32574
rect 31502 32498 31554 32510
rect 31726 32562 31778 32574
rect 31726 32498 31778 32510
rect 33854 32562 33906 32574
rect 33854 32498 33906 32510
rect 37326 32562 37378 32574
rect 37326 32498 37378 32510
rect 38110 32562 38162 32574
rect 38110 32498 38162 32510
rect 38782 32562 38834 32574
rect 49534 32562 49586 32574
rect 55358 32562 55410 32574
rect 56366 32562 56418 32574
rect 47618 32510 47630 32562
rect 47682 32510 47694 32562
rect 51538 32510 51550 32562
rect 51602 32510 51614 32562
rect 55682 32510 55694 32562
rect 55746 32510 55758 32562
rect 38782 32498 38834 32510
rect 49534 32498 49586 32510
rect 55358 32498 55410 32510
rect 56366 32498 56418 32510
rect 57710 32562 57762 32574
rect 57710 32498 57762 32510
rect 58158 32562 58210 32574
rect 58158 32498 58210 32510
rect 60062 32562 60114 32574
rect 60062 32498 60114 32510
rect 60398 32562 60450 32574
rect 62190 32562 62242 32574
rect 61506 32510 61518 32562
rect 61570 32510 61582 32562
rect 60398 32498 60450 32510
rect 62190 32498 62242 32510
rect 63198 32562 63250 32574
rect 63198 32498 63250 32510
rect 63534 32562 63586 32574
rect 63534 32498 63586 32510
rect 63758 32562 63810 32574
rect 67566 32562 67618 32574
rect 66770 32510 66782 32562
rect 66834 32510 66846 32562
rect 63758 32498 63810 32510
rect 67566 32498 67618 32510
rect 69918 32562 69970 32574
rect 69918 32498 69970 32510
rect 70590 32562 70642 32574
rect 74846 32562 74898 32574
rect 71138 32510 71150 32562
rect 71202 32510 71214 32562
rect 75170 32510 75182 32562
rect 75234 32510 75246 32562
rect 70590 32498 70642 32510
rect 74846 32498 74898 32510
rect 4174 32450 4226 32462
rect 16046 32450 16098 32462
rect 14130 32398 14142 32450
rect 14194 32398 14206 32450
rect 4174 32386 4226 32398
rect 16046 32386 16098 32398
rect 23438 32450 23490 32462
rect 28254 32450 28306 32462
rect 23986 32398 23998 32450
rect 24050 32398 24062 32450
rect 27570 32398 27582 32450
rect 27634 32398 27646 32450
rect 23438 32386 23490 32398
rect 28254 32386 28306 32398
rect 31390 32450 31442 32462
rect 31390 32386 31442 32398
rect 37102 32450 37154 32462
rect 37102 32386 37154 32398
rect 37662 32450 37714 32462
rect 37662 32386 37714 32398
rect 42254 32450 42306 32462
rect 42254 32386 42306 32398
rect 45390 32450 45442 32462
rect 45390 32386 45442 32398
rect 46174 32450 46226 32462
rect 53790 32450 53842 32462
rect 51426 32398 51438 32450
rect 51490 32398 51502 32450
rect 46174 32386 46226 32398
rect 53790 32386 53842 32398
rect 54350 32450 54402 32462
rect 62638 32450 62690 32462
rect 61730 32398 61742 32450
rect 61794 32398 61806 32450
rect 66658 32398 66670 32450
rect 66722 32398 66734 32450
rect 54350 32386 54402 32398
rect 62638 32386 62690 32398
rect 4398 32338 4450 32350
rect 29150 32338 29202 32350
rect 4722 32286 4734 32338
rect 4786 32286 4798 32338
rect 4398 32274 4450 32286
rect 29150 32274 29202 32286
rect 54574 32338 54626 32350
rect 76302 32338 76354 32350
rect 54898 32286 54910 32338
rect 54962 32286 54974 32338
rect 54574 32274 54626 32286
rect 76302 32274 76354 32286
rect 76638 32338 76690 32350
rect 76638 32274 76690 32286
rect 1344 32170 78624 32204
rect 1344 32118 10874 32170
rect 10926 32118 10978 32170
rect 11030 32118 11082 32170
rect 11134 32118 30194 32170
rect 30246 32118 30298 32170
rect 30350 32118 30402 32170
rect 30454 32118 49514 32170
rect 49566 32118 49618 32170
rect 49670 32118 49722 32170
rect 49774 32118 68834 32170
rect 68886 32118 68938 32170
rect 68990 32118 69042 32170
rect 69094 32118 78624 32170
rect 1344 32084 78624 32118
rect 37774 32002 37826 32014
rect 14130 31950 14142 32002
rect 14194 31950 14206 32002
rect 27570 31950 27582 32002
rect 27634 31950 27646 32002
rect 37774 31938 37826 31950
rect 59166 32002 59218 32014
rect 59166 31938 59218 31950
rect 60398 32002 60450 32014
rect 73390 32002 73442 32014
rect 70242 31950 70254 32002
rect 70306 31950 70318 32002
rect 60398 31938 60450 31950
rect 73390 31938 73442 31950
rect 4958 31890 5010 31902
rect 17726 31890 17778 31902
rect 22654 31890 22706 31902
rect 9202 31838 9214 31890
rect 9266 31838 9278 31890
rect 11442 31838 11454 31890
rect 11506 31838 11518 31890
rect 16930 31838 16942 31890
rect 16994 31838 17006 31890
rect 20290 31838 20302 31890
rect 20354 31838 20366 31890
rect 4958 31826 5010 31838
rect 17726 31826 17778 31838
rect 22654 31826 22706 31838
rect 23998 31890 24050 31902
rect 33406 31890 33458 31902
rect 37550 31890 37602 31902
rect 44046 31890 44098 31902
rect 26898 31838 26910 31890
rect 26962 31838 26974 31890
rect 31602 31838 31614 31890
rect 31666 31838 31678 31890
rect 33730 31838 33742 31890
rect 33794 31838 33806 31890
rect 38098 31838 38110 31890
rect 38162 31838 38174 31890
rect 40114 31838 40126 31890
rect 40178 31838 40190 31890
rect 41794 31838 41806 31890
rect 41858 31838 41870 31890
rect 23998 31826 24050 31838
rect 33406 31826 33458 31838
rect 37550 31826 37602 31838
rect 44046 31826 44098 31838
rect 46510 31890 46562 31902
rect 46510 31826 46562 31838
rect 61742 31890 61794 31902
rect 65886 31890 65938 31902
rect 63858 31838 63870 31890
rect 63922 31838 63934 31890
rect 61742 31826 61794 31838
rect 65886 31826 65938 31838
rect 74286 31890 74338 31902
rect 77310 31890 77362 31902
rect 75506 31838 75518 31890
rect 75570 31838 75582 31890
rect 74286 31826 74338 31838
rect 77310 31826 77362 31838
rect 78094 31890 78146 31902
rect 78094 31826 78146 31838
rect 4622 31778 4674 31790
rect 2930 31726 2942 31778
rect 2994 31726 3006 31778
rect 4622 31714 4674 31726
rect 5630 31778 5682 31790
rect 13918 31778 13970 31790
rect 20638 31778 20690 31790
rect 9314 31726 9326 31778
rect 9378 31726 9390 31778
rect 10658 31726 10670 31778
rect 10722 31726 10734 31778
rect 14130 31726 14142 31778
rect 14194 31726 14206 31778
rect 17042 31726 17054 31778
rect 17106 31726 17118 31778
rect 5630 31714 5682 31726
rect 13918 31714 13970 31726
rect 20638 31714 20690 31726
rect 20862 31778 20914 31790
rect 20862 31714 20914 31726
rect 21758 31778 21810 31790
rect 24894 31778 24946 31790
rect 32174 31778 32226 31790
rect 21970 31726 21982 31778
rect 22034 31726 22046 31778
rect 27234 31726 27246 31778
rect 27298 31726 27310 31778
rect 31266 31726 31278 31778
rect 31330 31726 31342 31778
rect 21758 31714 21810 31726
rect 24894 31714 24946 31726
rect 32174 31714 32226 31726
rect 33182 31778 33234 31790
rect 46398 31778 46450 31790
rect 39666 31726 39678 31778
rect 39730 31726 39742 31778
rect 41010 31726 41022 31778
rect 41074 31726 41086 31778
rect 43586 31726 43598 31778
rect 43650 31726 43662 31778
rect 43810 31726 43822 31778
rect 43874 31726 43886 31778
rect 46162 31726 46174 31778
rect 46226 31726 46238 31778
rect 33182 31714 33234 31726
rect 46398 31714 46450 31726
rect 47630 31778 47682 31790
rect 47630 31714 47682 31726
rect 49758 31778 49810 31790
rect 49758 31714 49810 31726
rect 49982 31778 50034 31790
rect 49982 31714 50034 31726
rect 54126 31778 54178 31790
rect 59502 31778 59554 31790
rect 55346 31726 55358 31778
rect 55410 31726 55422 31778
rect 56130 31726 56142 31778
rect 56194 31726 56206 31778
rect 54126 31714 54178 31726
rect 59502 31714 59554 31726
rect 60286 31778 60338 31790
rect 60286 31714 60338 31726
rect 61518 31778 61570 31790
rect 61518 31714 61570 31726
rect 61854 31778 61906 31790
rect 61854 31714 61906 31726
rect 63310 31778 63362 31790
rect 69794 31726 69806 31778
rect 69858 31726 69870 31778
rect 70802 31726 70814 31778
rect 70866 31726 70878 31778
rect 76178 31726 76190 31778
rect 76242 31726 76254 31778
rect 63310 31714 63362 31726
rect 3502 31666 3554 31678
rect 1922 31614 1934 31666
rect 1986 31614 1998 31666
rect 3502 31602 3554 31614
rect 4398 31666 4450 31678
rect 4398 31602 4450 31614
rect 6190 31666 6242 31678
rect 6190 31602 6242 31614
rect 15486 31666 15538 31678
rect 15486 31602 15538 31614
rect 15710 31666 15762 31678
rect 15710 31602 15762 31614
rect 24558 31666 24610 31678
rect 24558 31602 24610 31614
rect 46846 31666 46898 31678
rect 46846 31602 46898 31614
rect 47294 31666 47346 31678
rect 47294 31602 47346 31614
rect 51102 31666 51154 31678
rect 51102 31602 51154 31614
rect 52222 31666 52274 31678
rect 52222 31602 52274 31614
rect 53790 31666 53842 31678
rect 56814 31666 56866 31678
rect 54898 31614 54910 31666
rect 54962 31614 54974 31666
rect 53790 31602 53842 31614
rect 56814 31602 56866 31614
rect 59726 31666 59778 31678
rect 59726 31602 59778 31614
rect 60398 31666 60450 31678
rect 60398 31602 60450 31614
rect 62526 31666 62578 31678
rect 62526 31602 62578 31614
rect 65998 31666 66050 31678
rect 65998 31602 66050 31614
rect 66782 31666 66834 31678
rect 66782 31602 66834 31614
rect 69582 31666 69634 31678
rect 69582 31602 69634 31614
rect 71262 31666 71314 31678
rect 71262 31602 71314 31614
rect 72046 31666 72098 31678
rect 72046 31602 72098 31614
rect 73502 31666 73554 31678
rect 73502 31602 73554 31614
rect 74398 31666 74450 31678
rect 74398 31602 74450 31614
rect 77422 31666 77474 31678
rect 77422 31602 77474 31614
rect 6078 31554 6130 31566
rect 6078 31490 6130 31502
rect 6302 31554 6354 31566
rect 6302 31490 6354 31502
rect 11902 31554 11954 31566
rect 11902 31490 11954 31502
rect 15598 31554 15650 31566
rect 15598 31490 15650 31502
rect 16158 31554 16210 31566
rect 16158 31490 16210 31502
rect 24670 31554 24722 31566
rect 24670 31490 24722 31502
rect 25342 31554 25394 31566
rect 25342 31490 25394 31502
rect 30606 31554 30658 31566
rect 30606 31490 30658 31502
rect 39006 31554 39058 31566
rect 39006 31490 39058 31502
rect 46622 31554 46674 31566
rect 46622 31490 46674 31502
rect 47518 31554 47570 31566
rect 47518 31490 47570 31502
rect 48078 31554 48130 31566
rect 51214 31554 51266 31566
rect 50306 31502 50318 31554
rect 50370 31502 50382 31554
rect 48078 31490 48130 31502
rect 51214 31490 51266 31502
rect 51438 31554 51490 31566
rect 51438 31490 51490 31502
rect 51774 31554 51826 31566
rect 51774 31490 51826 31502
rect 53902 31554 53954 31566
rect 53902 31490 53954 31502
rect 57262 31554 57314 31566
rect 57262 31490 57314 31502
rect 57710 31554 57762 31566
rect 57710 31490 57762 31502
rect 58270 31554 58322 31566
rect 58270 31490 58322 31502
rect 61854 31554 61906 31566
rect 61854 31490 61906 31502
rect 62638 31554 62690 31566
rect 62638 31490 62690 31502
rect 63646 31554 63698 31566
rect 63646 31490 63698 31502
rect 63870 31554 63922 31566
rect 63870 31490 63922 31502
rect 64318 31554 64370 31566
rect 64318 31490 64370 31502
rect 65774 31554 65826 31566
rect 65774 31490 65826 31502
rect 66670 31554 66722 31566
rect 66670 31490 66722 31502
rect 67230 31554 67282 31566
rect 67230 31490 67282 31502
rect 68574 31554 68626 31566
rect 68574 31490 68626 31502
rect 71934 31554 71986 31566
rect 71934 31490 71986 31502
rect 73390 31554 73442 31566
rect 73390 31490 73442 31502
rect 74174 31554 74226 31566
rect 74174 31490 74226 31502
rect 77534 31554 77586 31566
rect 77534 31490 77586 31502
rect 1344 31386 78784 31420
rect 1344 31334 20534 31386
rect 20586 31334 20638 31386
rect 20690 31334 20742 31386
rect 20794 31334 39854 31386
rect 39906 31334 39958 31386
rect 40010 31334 40062 31386
rect 40114 31334 59174 31386
rect 59226 31334 59278 31386
rect 59330 31334 59382 31386
rect 59434 31334 78494 31386
rect 78546 31334 78598 31386
rect 78650 31334 78702 31386
rect 78754 31334 78784 31386
rect 1344 31300 78784 31334
rect 8878 31218 8930 31230
rect 8878 31154 8930 31166
rect 13470 31218 13522 31230
rect 13470 31154 13522 31166
rect 13694 31218 13746 31230
rect 13694 31154 13746 31166
rect 14702 31218 14754 31230
rect 14702 31154 14754 31166
rect 14814 31218 14866 31230
rect 14814 31154 14866 31166
rect 14926 31218 14978 31230
rect 14926 31154 14978 31166
rect 18622 31218 18674 31230
rect 18622 31154 18674 31166
rect 27694 31218 27746 31230
rect 48414 31218 48466 31230
rect 31714 31166 31726 31218
rect 31778 31166 31790 31218
rect 44146 31166 44158 31218
rect 44210 31166 44222 31218
rect 46498 31166 46510 31218
rect 46562 31166 46574 31218
rect 27694 31154 27746 31166
rect 48414 31154 48466 31166
rect 54350 31218 54402 31230
rect 54350 31154 54402 31166
rect 58494 31218 58546 31230
rect 67342 31218 67394 31230
rect 65538 31166 65550 31218
rect 65602 31166 65614 31218
rect 58494 31154 58546 31166
rect 67342 31154 67394 31166
rect 68238 31218 68290 31230
rect 68238 31154 68290 31166
rect 69582 31218 69634 31230
rect 69582 31154 69634 31166
rect 71822 31218 71874 31230
rect 71822 31154 71874 31166
rect 71934 31218 71986 31230
rect 71934 31154 71986 31166
rect 72270 31218 72322 31230
rect 72270 31154 72322 31166
rect 74622 31218 74674 31230
rect 74622 31154 74674 31166
rect 2718 31106 2770 31118
rect 2718 31042 2770 31054
rect 3054 31106 3106 31118
rect 3054 31042 3106 31054
rect 5966 31106 6018 31118
rect 5966 31042 6018 31054
rect 7086 31106 7138 31118
rect 7086 31042 7138 31054
rect 8206 31106 8258 31118
rect 8206 31042 8258 31054
rect 16942 31106 16994 31118
rect 16942 31042 16994 31054
rect 20638 31106 20690 31118
rect 20638 31042 20690 31054
rect 24334 31106 24386 31118
rect 24334 31042 24386 31054
rect 26686 31106 26738 31118
rect 26686 31042 26738 31054
rect 27806 31106 27858 31118
rect 27806 31042 27858 31054
rect 31166 31106 31218 31118
rect 37102 31106 37154 31118
rect 35522 31054 35534 31106
rect 35586 31054 35598 31106
rect 31166 31042 31218 31054
rect 37102 31042 37154 31054
rect 42030 31106 42082 31118
rect 42030 31042 42082 31054
rect 43598 31106 43650 31118
rect 55358 31106 55410 31118
rect 50418 31054 50430 31106
rect 50482 31054 50494 31106
rect 43598 31042 43650 31054
rect 55358 31042 55410 31054
rect 58606 31106 58658 31118
rect 58606 31042 58658 31054
rect 60734 31106 60786 31118
rect 60734 31042 60786 31054
rect 65998 31106 66050 31118
rect 65998 31042 66050 31054
rect 66894 31106 66946 31118
rect 66894 31042 66946 31054
rect 68462 31106 68514 31118
rect 68462 31042 68514 31054
rect 70254 31106 70306 31118
rect 70254 31042 70306 31054
rect 74846 31106 74898 31118
rect 74846 31042 74898 31054
rect 76862 31106 76914 31118
rect 76862 31042 76914 31054
rect 4510 30994 4562 31006
rect 6638 30994 6690 31006
rect 4162 30942 4174 30994
rect 4226 30942 4238 30994
rect 5170 30942 5182 30994
rect 5234 30942 5246 30994
rect 4510 30930 4562 30942
rect 6638 30930 6690 30942
rect 6862 30994 6914 31006
rect 6862 30930 6914 30942
rect 6974 30994 7026 31006
rect 13806 30994 13858 31006
rect 9762 30942 9774 30994
rect 9826 30942 9838 30994
rect 10434 30942 10446 30994
rect 10498 30942 10510 30994
rect 6974 30930 7026 30942
rect 13806 30930 13858 30942
rect 15374 30994 15426 31006
rect 18510 30994 18562 31006
rect 16034 30942 16046 30994
rect 16098 30942 16110 30994
rect 15374 30930 15426 30942
rect 18510 30930 18562 30942
rect 18734 30994 18786 31006
rect 18734 30930 18786 30942
rect 19182 30994 19234 31006
rect 27246 30994 27298 31006
rect 19954 30942 19966 30994
rect 20018 30942 20030 30994
rect 23874 30942 23886 30994
rect 23938 30942 23950 30994
rect 26002 30942 26014 30994
rect 26066 30942 26078 30994
rect 19182 30930 19234 30942
rect 27246 30930 27298 30942
rect 27470 30994 27522 31006
rect 31054 30994 31106 31006
rect 39342 30994 39394 31006
rect 30482 30942 30494 30994
rect 30546 30942 30558 30994
rect 36418 30942 36430 30994
rect 36482 30942 36494 30994
rect 27470 30930 27522 30942
rect 31054 30930 31106 30942
rect 39342 30930 39394 30942
rect 40462 30994 40514 31006
rect 41582 30994 41634 31006
rect 40786 30942 40798 30994
rect 40850 30942 40862 30994
rect 40462 30930 40514 30942
rect 41582 30930 41634 30942
rect 41806 30994 41858 31006
rect 41806 30930 41858 30942
rect 42142 30994 42194 31006
rect 42142 30930 42194 30942
rect 43822 30994 43874 31006
rect 43822 30930 43874 30942
rect 48750 30994 48802 31006
rect 54238 30994 54290 31006
rect 50306 30942 50318 30994
rect 50370 30942 50382 30994
rect 51538 30942 51550 30994
rect 51602 30942 51614 30994
rect 51874 30942 51886 30994
rect 51938 30942 51950 30994
rect 48750 30930 48802 30942
rect 54238 30930 54290 30942
rect 54462 30994 54514 31006
rect 54462 30930 54514 30942
rect 54910 30994 54962 31006
rect 54910 30930 54962 30942
rect 61070 30994 61122 31006
rect 61070 30930 61122 30942
rect 61630 30994 61682 31006
rect 61630 30930 61682 30942
rect 63198 30994 63250 31006
rect 63198 30930 63250 30942
rect 66110 30994 66162 31006
rect 67118 30994 67170 31006
rect 66322 30942 66334 30994
rect 66386 30942 66398 30994
rect 66110 30930 66162 30942
rect 67118 30930 67170 30942
rect 67566 30994 67618 31006
rect 67566 30930 67618 30942
rect 68574 30994 68626 31006
rect 69470 30994 69522 31006
rect 69122 30942 69134 30994
rect 69186 30942 69198 30994
rect 68574 30930 68626 30942
rect 69470 30930 69522 30942
rect 69694 30994 69746 31006
rect 72046 30994 72098 31006
rect 70690 30942 70702 30994
rect 70754 30942 70766 30994
rect 69694 30930 69746 30942
rect 72046 30930 72098 30942
rect 74958 30994 75010 31006
rect 74958 30930 75010 30942
rect 75966 30994 76018 31006
rect 75966 30930 76018 30942
rect 76078 30994 76130 31006
rect 76078 30930 76130 30942
rect 76190 30994 76242 31006
rect 77646 30994 77698 31006
rect 77074 30942 77086 30994
rect 77138 30942 77150 30994
rect 76190 30930 76242 30942
rect 77646 30930 77698 30942
rect 17614 30882 17666 30894
rect 22878 30882 22930 30894
rect 24894 30882 24946 30894
rect 29598 30882 29650 30894
rect 8978 30830 8990 30882
rect 9042 30830 9054 30882
rect 10098 30830 10110 30882
rect 10162 30830 10174 30882
rect 10322 30830 10334 30882
rect 10386 30830 10398 30882
rect 16706 30830 16718 30882
rect 16770 30830 16782 30882
rect 19730 30830 19742 30882
rect 19794 30830 19806 30882
rect 23426 30830 23438 30882
rect 23490 30830 23502 30882
rect 25890 30830 25902 30882
rect 25954 30830 25966 30882
rect 17614 30818 17666 30830
rect 22878 30818 22930 30830
rect 24894 30818 24946 30830
rect 29598 30818 29650 30830
rect 32286 30882 32338 30894
rect 32286 30818 32338 30830
rect 32734 30882 32786 30894
rect 32734 30818 32786 30830
rect 33854 30882 33906 30894
rect 33854 30818 33906 30830
rect 34414 30882 34466 30894
rect 39118 30882 39170 30894
rect 34962 30830 34974 30882
rect 35026 30830 35038 30882
rect 34414 30818 34466 30830
rect 39118 30818 39170 30830
rect 39678 30882 39730 30894
rect 39678 30818 39730 30830
rect 40238 30882 40290 30894
rect 40238 30818 40290 30830
rect 45390 30882 45442 30894
rect 45390 30818 45442 30830
rect 45950 30882 46002 30894
rect 45950 30818 46002 30830
rect 46174 30882 46226 30894
rect 46174 30818 46226 30830
rect 50990 30882 51042 30894
rect 50990 30818 51042 30830
rect 52446 30882 52498 30894
rect 52446 30818 52498 30830
rect 53566 30882 53618 30894
rect 53566 30818 53618 30830
rect 54686 30882 54738 30894
rect 54686 30818 54738 30830
rect 55806 30882 55858 30894
rect 55806 30818 55858 30830
rect 56254 30882 56306 30894
rect 56254 30818 56306 30830
rect 59726 30882 59778 30894
rect 59726 30818 59778 30830
rect 60174 30882 60226 30894
rect 63870 30882 63922 30894
rect 61954 30830 61966 30882
rect 62018 30830 62030 30882
rect 71138 30830 71150 30882
rect 71202 30830 71214 30882
rect 75506 30830 75518 30882
rect 75570 30830 75582 30882
rect 60174 30818 60226 30830
rect 63870 30818 63922 30830
rect 8654 30770 8706 30782
rect 8654 30706 8706 30718
rect 32062 30770 32114 30782
rect 32062 30706 32114 30718
rect 58382 30770 58434 30782
rect 63310 30770 63362 30782
rect 62178 30718 62190 30770
rect 62242 30718 62254 30770
rect 58382 30706 58434 30718
rect 63310 30706 63362 30718
rect 1344 30602 78624 30636
rect 1344 30550 10874 30602
rect 10926 30550 10978 30602
rect 11030 30550 11082 30602
rect 11134 30550 30194 30602
rect 30246 30550 30298 30602
rect 30350 30550 30402 30602
rect 30454 30550 49514 30602
rect 49566 30550 49618 30602
rect 49670 30550 49722 30602
rect 49774 30550 68834 30602
rect 68886 30550 68938 30602
rect 68990 30550 69042 30602
rect 69094 30550 78624 30602
rect 1344 30516 78624 30550
rect 4174 30434 4226 30446
rect 54798 30434 54850 30446
rect 19170 30382 19182 30434
rect 19234 30382 19246 30434
rect 4174 30370 4226 30382
rect 54798 30370 54850 30382
rect 55582 30434 55634 30446
rect 55582 30370 55634 30382
rect 57486 30434 57538 30446
rect 70702 30434 70754 30446
rect 70130 30382 70142 30434
rect 70194 30382 70206 30434
rect 57486 30370 57538 30382
rect 70702 30370 70754 30382
rect 71038 30434 71090 30446
rect 71698 30382 71710 30434
rect 71762 30382 71774 30434
rect 76402 30382 76414 30434
rect 76466 30431 76478 30434
rect 76738 30431 76750 30434
rect 76466 30385 76750 30431
rect 76466 30382 76478 30385
rect 76738 30382 76750 30385
rect 76802 30382 76814 30434
rect 71038 30370 71090 30382
rect 16606 30322 16658 30334
rect 23998 30322 24050 30334
rect 11554 30270 11566 30322
rect 11618 30270 11630 30322
rect 19282 30270 19294 30322
rect 19346 30270 19358 30322
rect 16606 30258 16658 30270
rect 23998 30258 24050 30270
rect 26014 30322 26066 30334
rect 26014 30258 26066 30270
rect 30942 30322 30994 30334
rect 30942 30258 30994 30270
rect 33854 30322 33906 30334
rect 35422 30322 35474 30334
rect 47854 30322 47906 30334
rect 34738 30270 34750 30322
rect 34802 30270 34814 30322
rect 44706 30270 44718 30322
rect 44770 30270 44782 30322
rect 33854 30258 33906 30270
rect 35422 30258 35474 30270
rect 47854 30258 47906 30270
rect 48302 30322 48354 30334
rect 48302 30258 48354 30270
rect 49758 30322 49810 30334
rect 57150 30322 57202 30334
rect 61406 30322 61458 30334
rect 72270 30322 72322 30334
rect 50530 30270 50542 30322
rect 50594 30270 50606 30322
rect 58370 30270 58382 30322
rect 58434 30270 58446 30322
rect 61730 30270 61742 30322
rect 61794 30270 61806 30322
rect 66994 30270 67006 30322
rect 67058 30270 67070 30322
rect 49758 30258 49810 30270
rect 57150 30258 57202 30270
rect 61406 30258 61458 30270
rect 72270 30258 72322 30270
rect 74398 30322 74450 30334
rect 74398 30258 74450 30270
rect 74510 30322 74562 30334
rect 75394 30270 75406 30322
rect 75458 30270 75470 30322
rect 74510 30258 74562 30270
rect 4062 30210 4114 30222
rect 4062 30146 4114 30158
rect 6750 30210 6802 30222
rect 7646 30210 7698 30222
rect 6962 30158 6974 30210
rect 7026 30158 7038 30210
rect 6750 30146 6802 30158
rect 7646 30146 7698 30158
rect 9438 30210 9490 30222
rect 9438 30146 9490 30158
rect 9774 30210 9826 30222
rect 9774 30146 9826 30158
rect 10334 30210 10386 30222
rect 10334 30146 10386 30158
rect 10558 30210 10610 30222
rect 10558 30146 10610 30158
rect 11006 30210 11058 30222
rect 12462 30210 12514 30222
rect 11778 30158 11790 30210
rect 11842 30158 11854 30210
rect 11006 30146 11058 30158
rect 12462 30146 12514 30158
rect 14030 30210 14082 30222
rect 14030 30146 14082 30158
rect 14366 30210 14418 30222
rect 14366 30146 14418 30158
rect 14814 30210 14866 30222
rect 14814 30146 14866 30158
rect 15038 30210 15090 30222
rect 15038 30146 15090 30158
rect 15822 30210 15874 30222
rect 15822 30146 15874 30158
rect 16158 30210 16210 30222
rect 23886 30210 23938 30222
rect 18946 30158 18958 30210
rect 19010 30158 19022 30210
rect 16158 30146 16210 30158
rect 23886 30146 23938 30158
rect 25790 30210 25842 30222
rect 30046 30210 30098 30222
rect 31502 30210 31554 30222
rect 26338 30158 26350 30210
rect 26402 30158 26414 30210
rect 30258 30158 30270 30210
rect 30322 30158 30334 30210
rect 25790 30146 25842 30158
rect 30046 30146 30098 30158
rect 31502 30146 31554 30158
rect 31838 30210 31890 30222
rect 31838 30146 31890 30158
rect 35310 30210 35362 30222
rect 35310 30146 35362 30158
rect 35982 30210 36034 30222
rect 35982 30146 36034 30158
rect 36318 30210 36370 30222
rect 36318 30146 36370 30158
rect 36654 30210 36706 30222
rect 36654 30146 36706 30158
rect 37438 30210 37490 30222
rect 53902 30210 53954 30222
rect 46050 30158 46062 30210
rect 46114 30158 46126 30210
rect 46946 30158 46958 30210
rect 47010 30158 47022 30210
rect 50418 30158 50430 30210
rect 50482 30158 50494 30210
rect 37438 30146 37490 30158
rect 53902 30146 53954 30158
rect 54238 30210 54290 30222
rect 66110 30210 66162 30222
rect 67566 30210 67618 30222
rect 58482 30158 58494 30210
rect 58546 30158 58558 30210
rect 62066 30158 62078 30210
rect 62130 30158 62142 30210
rect 66770 30158 66782 30210
rect 66834 30158 66846 30210
rect 54238 30146 54290 30158
rect 66110 30146 66162 30158
rect 67566 30146 67618 30158
rect 72046 30210 72098 30222
rect 72046 30146 72098 30158
rect 75070 30210 75122 30222
rect 77310 30210 77362 30222
rect 75506 30158 75518 30210
rect 75570 30158 75582 30210
rect 75070 30146 75122 30158
rect 77310 30146 77362 30158
rect 3166 30098 3218 30110
rect 3166 30034 3218 30046
rect 9550 30098 9602 30110
rect 9550 30034 9602 30046
rect 10446 30098 10498 30110
rect 10446 30034 10498 30046
rect 23550 30098 23602 30110
rect 23550 30034 23602 30046
rect 24110 30098 24162 30110
rect 24110 30034 24162 30046
rect 31614 30098 31666 30110
rect 31614 30034 31666 30046
rect 32174 30098 32226 30110
rect 32174 30034 32226 30046
rect 32734 30098 32786 30110
rect 32734 30034 32786 30046
rect 34414 30098 34466 30110
rect 34414 30034 34466 30046
rect 41694 30098 41746 30110
rect 41694 30034 41746 30046
rect 44382 30098 44434 30110
rect 47742 30098 47794 30110
rect 47170 30046 47182 30098
rect 47234 30046 47246 30098
rect 44382 30034 44434 30046
rect 47742 30034 47794 30046
rect 54686 30098 54738 30110
rect 54686 30034 54738 30046
rect 55694 30098 55746 30110
rect 55694 30034 55746 30046
rect 58158 30098 58210 30110
rect 58158 30034 58210 30046
rect 67790 30098 67842 30110
rect 67790 30034 67842 30046
rect 67902 30098 67954 30110
rect 67902 30034 67954 30046
rect 68462 30098 68514 30110
rect 68462 30034 68514 30046
rect 68574 30098 68626 30110
rect 68574 30034 68626 30046
rect 69470 30098 69522 30110
rect 69470 30034 69522 30046
rect 69582 30098 69634 30110
rect 69582 30034 69634 30046
rect 69694 30098 69746 30110
rect 69694 30034 69746 30046
rect 77534 30098 77586 30110
rect 77534 30034 77586 30046
rect 77758 30098 77810 30110
rect 77758 30034 77810 30046
rect 77870 30098 77922 30110
rect 77870 30034 77922 30046
rect 2382 29986 2434 29998
rect 2382 29922 2434 29934
rect 2830 29986 2882 29998
rect 2830 29922 2882 29934
rect 4174 29986 4226 29998
rect 4174 29922 4226 29934
rect 4846 29986 4898 29998
rect 4846 29922 4898 29934
rect 12910 29986 12962 29998
rect 12910 29922 12962 29934
rect 14142 29986 14194 29998
rect 16046 29986 16098 29998
rect 15362 29934 15374 29986
rect 15426 29934 15438 29986
rect 14142 29922 14194 29934
rect 16046 29922 16098 29934
rect 17166 29986 17218 29998
rect 17166 29922 17218 29934
rect 22990 29986 23042 29998
rect 22990 29922 23042 29934
rect 24894 29986 24946 29998
rect 24894 29922 24946 29934
rect 25230 29986 25282 29998
rect 25230 29922 25282 29934
rect 26910 29986 26962 29998
rect 26910 29922 26962 29934
rect 27358 29986 27410 29998
rect 27358 29922 27410 29934
rect 28142 29986 28194 29998
rect 28142 29922 28194 29934
rect 28814 29986 28866 29998
rect 28814 29922 28866 29934
rect 32846 29986 32898 29998
rect 32846 29922 32898 29934
rect 33070 29986 33122 29998
rect 33070 29922 33122 29934
rect 33406 29986 33458 29998
rect 33406 29922 33458 29934
rect 34638 29986 34690 29998
rect 34638 29922 34690 29934
rect 35534 29986 35586 29998
rect 35534 29922 35586 29934
rect 36542 29986 36594 29998
rect 36542 29922 36594 29934
rect 41358 29986 41410 29998
rect 41358 29922 41410 29934
rect 43822 29986 43874 29998
rect 43822 29922 43874 29934
rect 44606 29986 44658 29998
rect 53454 29986 53506 29998
rect 46274 29934 46286 29986
rect 46338 29934 46350 29986
rect 44606 29922 44658 29934
rect 53454 29922 53506 29934
rect 54014 29986 54066 29998
rect 54014 29922 54066 29934
rect 54798 29986 54850 29998
rect 54798 29922 54850 29934
rect 55582 29986 55634 29998
rect 55582 29922 55634 29934
rect 56254 29986 56306 29998
rect 56254 29922 56306 29934
rect 56702 29986 56754 29998
rect 56702 29922 56754 29934
rect 57374 29986 57426 29998
rect 57374 29922 57426 29934
rect 60622 29986 60674 29998
rect 60622 29922 60674 29934
rect 70814 29986 70866 29998
rect 70814 29922 70866 29934
rect 72718 29986 72770 29998
rect 72718 29922 72770 29934
rect 74286 29986 74338 29998
rect 74286 29922 74338 29934
rect 76638 29986 76690 29998
rect 76638 29922 76690 29934
rect 1344 29818 78784 29852
rect 1344 29766 20534 29818
rect 20586 29766 20638 29818
rect 20690 29766 20742 29818
rect 20794 29766 39854 29818
rect 39906 29766 39958 29818
rect 40010 29766 40062 29818
rect 40114 29766 59174 29818
rect 59226 29766 59278 29818
rect 59330 29766 59382 29818
rect 59434 29766 78494 29818
rect 78546 29766 78598 29818
rect 78650 29766 78702 29818
rect 78754 29766 78784 29818
rect 1344 29732 78784 29766
rect 9886 29650 9938 29662
rect 9886 29586 9938 29598
rect 12126 29650 12178 29662
rect 12126 29586 12178 29598
rect 13918 29650 13970 29662
rect 13918 29586 13970 29598
rect 16382 29650 16434 29662
rect 28590 29650 28642 29662
rect 19506 29598 19518 29650
rect 19570 29598 19582 29650
rect 16382 29586 16434 29598
rect 28590 29586 28642 29598
rect 28814 29650 28866 29662
rect 28814 29586 28866 29598
rect 29822 29650 29874 29662
rect 29822 29586 29874 29598
rect 33966 29650 34018 29662
rect 33966 29586 34018 29598
rect 36094 29650 36146 29662
rect 36094 29586 36146 29598
rect 40462 29650 40514 29662
rect 40462 29586 40514 29598
rect 51102 29650 51154 29662
rect 51102 29586 51154 29598
rect 60734 29650 60786 29662
rect 60734 29586 60786 29598
rect 63646 29650 63698 29662
rect 63646 29586 63698 29598
rect 70702 29650 70754 29662
rect 70702 29586 70754 29598
rect 71710 29650 71762 29662
rect 71710 29586 71762 29598
rect 4622 29538 4674 29550
rect 4622 29474 4674 29486
rect 6526 29538 6578 29550
rect 6526 29474 6578 29486
rect 12350 29538 12402 29550
rect 12350 29474 12402 29486
rect 15486 29538 15538 29550
rect 15486 29474 15538 29486
rect 18286 29538 18338 29550
rect 18286 29474 18338 29486
rect 21310 29538 21362 29550
rect 21310 29474 21362 29486
rect 23998 29538 24050 29550
rect 23998 29474 24050 29486
rect 26910 29538 26962 29550
rect 26910 29474 26962 29486
rect 33630 29538 33682 29550
rect 33630 29474 33682 29486
rect 33742 29538 33794 29550
rect 33742 29474 33794 29486
rect 37886 29538 37938 29550
rect 45950 29538 46002 29550
rect 43698 29486 43710 29538
rect 43762 29486 43774 29538
rect 37886 29474 37938 29486
rect 45950 29474 46002 29486
rect 46510 29538 46562 29550
rect 46510 29474 46562 29486
rect 51326 29538 51378 29550
rect 51326 29474 51378 29486
rect 53006 29538 53058 29550
rect 53006 29474 53058 29486
rect 54910 29538 54962 29550
rect 54910 29474 54962 29486
rect 59726 29538 59778 29550
rect 59726 29474 59778 29486
rect 59838 29538 59890 29550
rect 59838 29474 59890 29486
rect 63870 29538 63922 29550
rect 63870 29474 63922 29486
rect 67790 29538 67842 29550
rect 67790 29474 67842 29486
rect 68238 29538 68290 29550
rect 68238 29474 68290 29486
rect 71486 29538 71538 29550
rect 71486 29474 71538 29486
rect 4510 29426 4562 29438
rect 12462 29426 12514 29438
rect 18062 29426 18114 29438
rect 2818 29374 2830 29426
rect 2882 29374 2894 29426
rect 4162 29374 4174 29426
rect 4226 29374 4238 29426
rect 7186 29374 7198 29426
rect 7250 29374 7262 29426
rect 11442 29374 11454 29426
rect 11506 29374 11518 29426
rect 14802 29374 14814 29426
rect 14866 29374 14878 29426
rect 4510 29362 4562 29374
rect 12462 29362 12514 29374
rect 18062 29362 18114 29374
rect 18398 29426 18450 29438
rect 23102 29426 23154 29438
rect 22418 29374 22430 29426
rect 22482 29374 22494 29426
rect 18398 29362 18450 29374
rect 23102 29362 23154 29374
rect 23662 29426 23714 29438
rect 27806 29426 27858 29438
rect 27346 29374 27358 29426
rect 27410 29374 27422 29426
rect 23662 29362 23714 29374
rect 27806 29362 27858 29374
rect 28478 29426 28530 29438
rect 40126 29426 40178 29438
rect 32386 29374 32398 29426
rect 32450 29374 32462 29426
rect 37314 29374 37326 29426
rect 37378 29374 37390 29426
rect 28478 29362 28530 29374
rect 40126 29362 40178 29374
rect 40574 29426 40626 29438
rect 40574 29362 40626 29374
rect 40686 29426 40738 29438
rect 46846 29426 46898 29438
rect 41794 29374 41806 29426
rect 41858 29374 41870 29426
rect 43138 29374 43150 29426
rect 43202 29374 43214 29426
rect 45266 29374 45278 29426
rect 45330 29374 45342 29426
rect 40686 29362 40738 29374
rect 46846 29362 46898 29374
rect 49646 29426 49698 29438
rect 51438 29426 51490 29438
rect 50194 29374 50206 29426
rect 50258 29374 50270 29426
rect 49646 29362 49698 29374
rect 51438 29362 51490 29374
rect 54574 29426 54626 29438
rect 54574 29362 54626 29374
rect 54686 29426 54738 29438
rect 54686 29362 54738 29374
rect 55134 29426 55186 29438
rect 59502 29426 59554 29438
rect 56242 29374 56254 29426
rect 56306 29374 56318 29426
rect 58594 29374 58606 29426
rect 58658 29374 58670 29426
rect 55134 29362 55186 29374
rect 59502 29362 59554 29374
rect 63982 29426 64034 29438
rect 63982 29362 64034 29374
rect 64542 29426 64594 29438
rect 64542 29362 64594 29374
rect 70814 29426 70866 29438
rect 70814 29362 70866 29374
rect 71374 29426 71426 29438
rect 75170 29374 75182 29426
rect 75234 29374 75246 29426
rect 71374 29362 71426 29374
rect 5070 29314 5122 29326
rect 7982 29314 8034 29326
rect 1922 29262 1934 29314
rect 1986 29262 1998 29314
rect 6850 29262 6862 29314
rect 6914 29262 6926 29314
rect 5070 29250 5122 29262
rect 7982 29250 8034 29262
rect 10670 29314 10722 29326
rect 12910 29314 12962 29326
rect 11330 29262 11342 29314
rect 11394 29262 11406 29314
rect 10670 29250 10722 29262
rect 12910 29250 12962 29262
rect 13358 29314 13410 29326
rect 18958 29314 19010 29326
rect 21534 29314 21586 29326
rect 24558 29314 24610 29326
rect 15026 29262 15038 29314
rect 15090 29262 15102 29314
rect 21186 29262 21198 29314
rect 21250 29262 21262 29314
rect 22194 29262 22206 29314
rect 22258 29262 22270 29314
rect 13358 29250 13410 29262
rect 18958 29250 19010 29262
rect 21534 29250 21586 29262
rect 24558 29250 24610 29262
rect 25902 29314 25954 29326
rect 25902 29250 25954 29262
rect 26350 29314 26402 29326
rect 26350 29250 26402 29262
rect 29374 29314 29426 29326
rect 32734 29314 32786 29326
rect 38558 29314 38610 29326
rect 32050 29262 32062 29314
rect 32114 29262 32126 29314
rect 37090 29262 37102 29314
rect 37154 29262 37166 29314
rect 29374 29250 29426 29262
rect 32734 29250 32786 29262
rect 38558 29250 38610 29262
rect 39118 29314 39170 29326
rect 39118 29250 39170 29262
rect 39678 29314 39730 29326
rect 44382 29314 44434 29326
rect 48190 29314 48242 29326
rect 56590 29314 56642 29326
rect 60286 29314 60338 29326
rect 41682 29262 41694 29314
rect 41746 29262 41758 29314
rect 45042 29262 45054 29314
rect 45106 29262 45118 29314
rect 50418 29262 50430 29314
rect 50482 29262 50494 29314
rect 55906 29262 55918 29314
rect 55970 29262 55982 29314
rect 58146 29262 58158 29314
rect 58210 29262 58222 29314
rect 39678 29250 39730 29262
rect 44382 29250 44434 29262
rect 48190 29250 48242 29262
rect 56590 29250 56642 29262
rect 60286 29250 60338 29262
rect 64654 29314 64706 29326
rect 64654 29250 64706 29262
rect 67342 29314 67394 29326
rect 67342 29250 67394 29262
rect 68798 29314 68850 29326
rect 68798 29250 68850 29262
rect 70030 29314 70082 29326
rect 70030 29250 70082 29262
rect 72046 29314 72098 29326
rect 76750 29314 76802 29326
rect 76066 29262 76078 29314
rect 76130 29262 76142 29314
rect 72046 29250 72098 29262
rect 76750 29250 76802 29262
rect 77086 29314 77138 29326
rect 77086 29250 77138 29262
rect 77646 29314 77698 29326
rect 77646 29250 77698 29262
rect 77982 29314 78034 29326
rect 77982 29250 78034 29262
rect 19182 29202 19234 29214
rect 19182 29138 19234 29150
rect 39342 29202 39394 29214
rect 39342 29138 39394 29150
rect 48414 29202 48466 29214
rect 48414 29138 48466 29150
rect 48750 29202 48802 29214
rect 48750 29138 48802 29150
rect 52782 29202 52834 29214
rect 52782 29138 52834 29150
rect 53118 29202 53170 29214
rect 70702 29202 70754 29214
rect 58930 29150 58942 29202
rect 58994 29150 59006 29202
rect 76626 29150 76638 29202
rect 76690 29199 76702 29202
rect 77634 29199 77646 29202
rect 76690 29153 77646 29199
rect 76690 29150 76702 29153
rect 77634 29150 77646 29153
rect 77698 29150 77710 29202
rect 53118 29138 53170 29150
rect 70702 29138 70754 29150
rect 1344 29034 78624 29068
rect 1344 28982 10874 29034
rect 10926 28982 10978 29034
rect 11030 28982 11082 29034
rect 11134 28982 30194 29034
rect 30246 28982 30298 29034
rect 30350 28982 30402 29034
rect 30454 28982 49514 29034
rect 49566 28982 49618 29034
rect 49670 28982 49722 29034
rect 49774 28982 68834 29034
rect 68886 28982 68938 29034
rect 68990 28982 69042 29034
rect 69094 28982 78624 29034
rect 1344 28948 78624 28982
rect 14254 28866 14306 28878
rect 6738 28814 6750 28866
rect 6802 28814 6814 28866
rect 10658 28814 10670 28866
rect 10722 28814 10734 28866
rect 14254 28802 14306 28814
rect 28814 28866 28866 28878
rect 28814 28802 28866 28814
rect 33742 28866 33794 28878
rect 40910 28866 40962 28878
rect 40562 28814 40574 28866
rect 40626 28814 40638 28866
rect 33742 28802 33794 28814
rect 40910 28802 40962 28814
rect 69470 28866 69522 28878
rect 77298 28814 77310 28866
rect 77362 28814 77374 28866
rect 69470 28802 69522 28814
rect 3614 28754 3666 28766
rect 14814 28754 14866 28766
rect 4946 28702 4958 28754
rect 5010 28702 5022 28754
rect 10434 28702 10446 28754
rect 10498 28702 10510 28754
rect 3614 28690 3666 28702
rect 14814 28690 14866 28702
rect 17838 28754 17890 28766
rect 22878 28754 22930 28766
rect 30606 28754 30658 28766
rect 18610 28702 18622 28754
rect 18674 28702 18686 28754
rect 20850 28702 20862 28754
rect 20914 28702 20926 28754
rect 24770 28702 24782 28754
rect 24834 28702 24846 28754
rect 27010 28702 27022 28754
rect 27074 28702 27086 28754
rect 17838 28690 17890 28702
rect 22878 28690 22930 28702
rect 30606 28690 30658 28702
rect 32062 28754 32114 28766
rect 40014 28754 40066 28766
rect 32386 28702 32398 28754
rect 32450 28702 32462 28754
rect 32062 28690 32114 28702
rect 40014 28690 40066 28702
rect 41134 28754 41186 28766
rect 52334 28754 52386 28766
rect 46386 28702 46398 28754
rect 46450 28702 46462 28754
rect 41134 28690 41186 28702
rect 52334 28690 52386 28702
rect 65102 28754 65154 28766
rect 73838 28754 73890 28766
rect 77870 28754 77922 28766
rect 65762 28702 65774 28754
rect 65826 28702 65838 28754
rect 71474 28702 71486 28754
rect 71538 28702 71550 28754
rect 74610 28702 74622 28754
rect 74674 28702 74686 28754
rect 76178 28702 76190 28754
rect 76242 28702 76254 28754
rect 65102 28690 65154 28702
rect 73838 28690 73890 28702
rect 77870 28690 77922 28702
rect 7086 28642 7138 28654
rect 7086 28578 7138 28590
rect 7310 28642 7362 28654
rect 7310 28578 7362 28590
rect 7758 28642 7810 28654
rect 12126 28642 12178 28654
rect 10322 28590 10334 28642
rect 10386 28590 10398 28642
rect 7758 28578 7810 28590
rect 12126 28578 12178 28590
rect 12574 28642 12626 28654
rect 12574 28578 12626 28590
rect 14590 28642 14642 28654
rect 14590 28578 14642 28590
rect 15374 28642 15426 28654
rect 15374 28578 15426 28590
rect 17726 28642 17778 28654
rect 23998 28642 24050 28654
rect 25566 28642 25618 28654
rect 18834 28590 18846 28642
rect 18898 28590 18910 28642
rect 20178 28590 20190 28642
rect 20242 28590 20254 28642
rect 24434 28590 24446 28642
rect 24498 28590 24510 28642
rect 17726 28578 17778 28590
rect 23998 28578 24050 28590
rect 25566 28578 25618 28590
rect 26462 28642 26514 28654
rect 26462 28578 26514 28590
rect 28478 28642 28530 28654
rect 28478 28578 28530 28590
rect 29710 28642 29762 28654
rect 31614 28642 31666 28654
rect 34302 28642 34354 28654
rect 29922 28590 29934 28642
rect 29986 28590 29998 28642
rect 32498 28590 32510 28642
rect 32562 28590 32574 28642
rect 29710 28578 29762 28590
rect 31614 28578 31666 28590
rect 34302 28578 34354 28590
rect 36878 28642 36930 28654
rect 36878 28578 36930 28590
rect 37438 28642 37490 28654
rect 48302 28642 48354 28654
rect 46610 28590 46622 28642
rect 46674 28590 46686 28642
rect 37438 28578 37490 28590
rect 48302 28578 48354 28590
rect 48638 28642 48690 28654
rect 48638 28578 48690 28590
rect 49870 28642 49922 28654
rect 49870 28578 49922 28590
rect 50318 28642 50370 28654
rect 50318 28578 50370 28590
rect 54014 28642 54066 28654
rect 54014 28578 54066 28590
rect 56030 28642 56082 28654
rect 56030 28578 56082 28590
rect 58830 28642 58882 28654
rect 58830 28578 58882 28590
rect 59726 28642 59778 28654
rect 64206 28642 64258 28654
rect 67342 28642 67394 28654
rect 71934 28642 71986 28654
rect 75406 28642 75458 28654
rect 77646 28642 77698 28654
rect 60162 28590 60174 28642
rect 60226 28590 60238 28642
rect 61954 28590 61966 28642
rect 62018 28590 62030 28642
rect 64642 28590 64654 28642
rect 64706 28590 64718 28642
rect 65986 28590 65998 28642
rect 66050 28590 66062 28642
rect 67554 28590 67566 28642
rect 67618 28590 67630 28642
rect 71026 28590 71038 28642
rect 71090 28590 71102 28642
rect 74498 28590 74510 28642
rect 74562 28590 74574 28642
rect 76290 28590 76302 28642
rect 76354 28590 76366 28642
rect 59726 28578 59778 28590
rect 64206 28578 64258 28590
rect 67342 28578 67394 28590
rect 71934 28578 71986 28590
rect 75406 28578 75458 28590
rect 77646 28578 77698 28590
rect 2830 28530 2882 28542
rect 2830 28466 2882 28478
rect 3166 28530 3218 28542
rect 3166 28466 3218 28478
rect 4622 28530 4674 28542
rect 4622 28466 4674 28478
rect 13806 28530 13858 28542
rect 13806 28466 13858 28478
rect 17390 28530 17442 28542
rect 17390 28466 17442 28478
rect 17950 28530 18002 28542
rect 17950 28466 18002 28478
rect 25902 28530 25954 28542
rect 25902 28466 25954 28478
rect 27582 28530 27634 28542
rect 27582 28466 27634 28478
rect 28702 28530 28754 28542
rect 28702 28466 28754 28478
rect 33630 28530 33682 28542
rect 33630 28466 33682 28478
rect 33742 28530 33794 28542
rect 33742 28466 33794 28478
rect 36542 28530 36594 28542
rect 36542 28466 36594 28478
rect 37998 28530 38050 28542
rect 37998 28466 38050 28478
rect 47294 28530 47346 28542
rect 47294 28466 47346 28478
rect 48414 28530 48466 28542
rect 48414 28466 48466 28478
rect 50430 28530 50482 28542
rect 50430 28466 50482 28478
rect 50542 28530 50594 28542
rect 50542 28466 50594 28478
rect 53454 28530 53506 28542
rect 53454 28466 53506 28478
rect 54574 28530 54626 28542
rect 54574 28466 54626 28478
rect 54798 28530 54850 28542
rect 54798 28466 54850 28478
rect 55246 28530 55298 28542
rect 55246 28466 55298 28478
rect 55582 28530 55634 28542
rect 55582 28466 55634 28478
rect 58158 28530 58210 28542
rect 58158 28466 58210 28478
rect 60622 28530 60674 28542
rect 60622 28466 60674 28478
rect 61406 28530 61458 28542
rect 61406 28466 61458 28478
rect 61518 28530 61570 28542
rect 61518 28466 61570 28478
rect 66670 28530 66722 28542
rect 66670 28466 66722 28478
rect 68238 28530 68290 28542
rect 68238 28466 68290 28478
rect 69470 28530 69522 28542
rect 69470 28466 69522 28478
rect 69582 28530 69634 28542
rect 69582 28466 69634 28478
rect 4846 28418 4898 28430
rect 4846 28354 4898 28366
rect 5630 28418 5682 28430
rect 5630 28354 5682 28366
rect 16942 28418 16994 28430
rect 16942 28354 16994 28366
rect 22430 28418 22482 28430
rect 22430 28354 22482 28366
rect 22990 28418 23042 28430
rect 22990 28354 23042 28366
rect 23438 28418 23490 28430
rect 23438 28354 23490 28366
rect 25790 28418 25842 28430
rect 25790 28354 25842 28366
rect 26798 28418 26850 28430
rect 26798 28354 26850 28366
rect 27022 28418 27074 28430
rect 27022 28354 27074 28366
rect 27694 28418 27746 28430
rect 27694 28354 27746 28366
rect 27918 28418 27970 28430
rect 27918 28354 27970 28366
rect 31166 28418 31218 28430
rect 31166 28354 31218 28366
rect 35646 28418 35698 28430
rect 35646 28354 35698 28366
rect 36094 28418 36146 28430
rect 36094 28354 36146 28366
rect 36654 28418 36706 28430
rect 36654 28354 36706 28366
rect 37886 28418 37938 28430
rect 37886 28354 37938 28366
rect 38110 28418 38162 28430
rect 38110 28354 38162 28366
rect 52446 28418 52498 28430
rect 52446 28354 52498 28366
rect 53678 28418 53730 28430
rect 53678 28354 53730 28366
rect 53902 28418 53954 28430
rect 53902 28354 53954 28366
rect 54686 28418 54738 28430
rect 54686 28354 54738 28366
rect 55470 28418 55522 28430
rect 55470 28354 55522 28366
rect 58270 28418 58322 28430
rect 58270 28354 58322 28366
rect 58494 28418 58546 28430
rect 58494 28354 58546 28366
rect 61630 28418 61682 28430
rect 61630 28354 61682 28366
rect 1344 28250 78784 28284
rect 1344 28198 20534 28250
rect 20586 28198 20638 28250
rect 20690 28198 20742 28250
rect 20794 28198 39854 28250
rect 39906 28198 39958 28250
rect 40010 28198 40062 28250
rect 40114 28198 59174 28250
rect 59226 28198 59278 28250
rect 59330 28198 59382 28250
rect 59434 28198 78494 28250
rect 78546 28198 78598 28250
rect 78650 28198 78702 28250
rect 78754 28198 78784 28250
rect 1344 28164 78784 28198
rect 5294 28082 5346 28094
rect 5294 28018 5346 28030
rect 5406 28082 5458 28094
rect 5406 28018 5458 28030
rect 6526 28082 6578 28094
rect 6526 28018 6578 28030
rect 13918 28082 13970 28094
rect 13918 28018 13970 28030
rect 14702 28082 14754 28094
rect 19070 28082 19122 28094
rect 18274 28030 18286 28082
rect 18338 28030 18350 28082
rect 14702 28018 14754 28030
rect 19070 28018 19122 28030
rect 23662 28082 23714 28094
rect 23662 28018 23714 28030
rect 24894 28082 24946 28094
rect 24894 28018 24946 28030
rect 28702 28082 28754 28094
rect 56814 28082 56866 28094
rect 42130 28030 42142 28082
rect 42194 28030 42206 28082
rect 28702 28018 28754 28030
rect 56814 28018 56866 28030
rect 61966 28082 62018 28094
rect 71486 28082 71538 28094
rect 76526 28082 76578 28094
rect 65426 28030 65438 28082
rect 65490 28030 65502 28082
rect 75058 28030 75070 28082
rect 75122 28030 75134 28082
rect 61966 28018 62018 28030
rect 71486 28018 71538 28030
rect 76526 28018 76578 28030
rect 4734 27970 4786 27982
rect 3154 27918 3166 27970
rect 3218 27918 3230 27970
rect 4734 27906 4786 27918
rect 8766 27970 8818 27982
rect 8766 27906 8818 27918
rect 13358 27970 13410 27982
rect 13358 27906 13410 27918
rect 14142 27970 14194 27982
rect 14142 27906 14194 27918
rect 14926 27970 14978 27982
rect 14926 27906 14978 27918
rect 19182 27970 19234 27982
rect 19182 27906 19234 27918
rect 22430 27970 22482 27982
rect 22430 27906 22482 27918
rect 26798 27970 26850 27982
rect 26798 27906 26850 27918
rect 28142 27970 28194 27982
rect 28142 27906 28194 27918
rect 28590 27970 28642 27982
rect 28590 27906 28642 27918
rect 30718 27970 30770 27982
rect 30718 27906 30770 27918
rect 37214 27970 37266 27982
rect 37214 27906 37266 27918
rect 40798 27970 40850 27982
rect 40798 27906 40850 27918
rect 46286 27970 46338 27982
rect 54574 27970 54626 27982
rect 53778 27918 53790 27970
rect 53842 27918 53854 27970
rect 46286 27906 46338 27918
rect 54574 27906 54626 27918
rect 56590 27970 56642 27982
rect 56590 27906 56642 27918
rect 59278 27970 59330 27982
rect 59278 27906 59330 27918
rect 61406 27970 61458 27982
rect 61406 27906 61458 27918
rect 61854 27970 61906 27982
rect 61854 27906 61906 27918
rect 62862 27970 62914 27982
rect 62862 27906 62914 27918
rect 65998 27970 66050 27982
rect 65998 27906 66050 27918
rect 70030 27970 70082 27982
rect 70030 27906 70082 27918
rect 71374 27970 71426 27982
rect 71374 27906 71426 27918
rect 71598 27970 71650 27982
rect 71598 27906 71650 27918
rect 75518 27970 75570 27982
rect 75518 27906 75570 27918
rect 75742 27970 75794 27982
rect 75742 27906 75794 27918
rect 76750 27970 76802 27982
rect 76750 27906 76802 27918
rect 77758 27970 77810 27982
rect 77758 27906 77810 27918
rect 5518 27858 5570 27870
rect 3378 27806 3390 27858
rect 3442 27806 3454 27858
rect 4274 27806 4286 27858
rect 4338 27806 4350 27858
rect 5518 27794 5570 27806
rect 5966 27858 6018 27870
rect 5966 27794 6018 27806
rect 6302 27858 6354 27870
rect 6302 27794 6354 27806
rect 6638 27858 6690 27870
rect 13246 27858 13298 27870
rect 8306 27806 8318 27858
rect 8370 27806 8382 27858
rect 10994 27806 11006 27858
rect 11058 27806 11070 27858
rect 6638 27794 6690 27806
rect 13246 27794 13298 27806
rect 13582 27858 13634 27870
rect 13582 27794 13634 27806
rect 14254 27858 14306 27870
rect 14254 27794 14306 27806
rect 15038 27858 15090 27870
rect 21870 27858 21922 27870
rect 28030 27858 28082 27870
rect 18834 27806 18846 27858
rect 18898 27806 18910 27858
rect 22642 27806 22654 27858
rect 22706 27806 22718 27858
rect 22866 27806 22878 27858
rect 22930 27806 22942 27858
rect 26562 27806 26574 27858
rect 26626 27806 26638 27858
rect 27346 27806 27358 27858
rect 27410 27806 27422 27858
rect 15038 27794 15090 27806
rect 21870 27794 21922 27806
rect 28030 27794 28082 27806
rect 28926 27858 28978 27870
rect 28926 27794 28978 27806
rect 29038 27858 29090 27870
rect 29038 27794 29090 27806
rect 30046 27858 30098 27870
rect 30046 27794 30098 27806
rect 30830 27858 30882 27870
rect 45278 27858 45330 27870
rect 31602 27806 31614 27858
rect 31666 27806 31678 27858
rect 36306 27806 36318 27858
rect 36370 27806 36382 27858
rect 40114 27806 40126 27858
rect 40178 27806 40190 27858
rect 45042 27806 45054 27858
rect 45106 27806 45118 27858
rect 30830 27794 30882 27806
rect 45278 27794 45330 27806
rect 46062 27858 46114 27870
rect 46062 27794 46114 27806
rect 46622 27858 46674 27870
rect 54686 27858 54738 27870
rect 49858 27806 49870 27858
rect 49922 27806 49934 27858
rect 52546 27806 52558 27858
rect 52610 27806 52622 27858
rect 52882 27806 52894 27858
rect 52946 27806 52958 27858
rect 53554 27806 53566 27858
rect 53618 27806 53630 27858
rect 54338 27806 54350 27858
rect 54402 27806 54414 27858
rect 46622 27794 46674 27806
rect 54686 27794 54738 27806
rect 56478 27858 56530 27870
rect 60398 27858 60450 27870
rect 62750 27858 62802 27870
rect 58482 27806 58494 27858
rect 58546 27806 58558 27858
rect 61618 27806 61630 27858
rect 61682 27806 61694 27858
rect 56478 27794 56530 27806
rect 60398 27794 60450 27806
rect 62750 27794 62802 27806
rect 63086 27858 63138 27870
rect 63086 27794 63138 27806
rect 65774 27858 65826 27870
rect 75630 27858 75682 27870
rect 69458 27806 69470 27858
rect 69522 27806 69534 27858
rect 65774 27794 65826 27806
rect 75630 27794 75682 27806
rect 76414 27858 76466 27870
rect 76414 27794 76466 27806
rect 76974 27858 77026 27870
rect 76974 27794 77026 27806
rect 7086 27746 7138 27758
rect 10446 27746 10498 27758
rect 12014 27746 12066 27758
rect 7858 27694 7870 27746
rect 7922 27694 7934 27746
rect 11106 27694 11118 27746
rect 11170 27694 11182 27746
rect 7086 27682 7138 27694
rect 10446 27682 10498 27694
rect 12014 27682 12066 27694
rect 12686 27746 12738 27758
rect 12686 27682 12738 27694
rect 15598 27746 15650 27758
rect 15598 27682 15650 27694
rect 15934 27746 15986 27758
rect 15934 27682 15986 27694
rect 16494 27746 16546 27758
rect 16494 27682 16546 27694
rect 17054 27746 17106 27758
rect 17054 27682 17106 27694
rect 17726 27746 17778 27758
rect 17726 27682 17778 27694
rect 19742 27746 19794 27758
rect 19742 27682 19794 27694
rect 20078 27746 20130 27758
rect 20078 27682 20130 27694
rect 20526 27746 20578 27758
rect 20526 27682 20578 27694
rect 21086 27746 21138 27758
rect 21086 27682 21138 27694
rect 21422 27746 21474 27758
rect 21422 27682 21474 27694
rect 22766 27746 22818 27758
rect 22766 27682 22818 27694
rect 24222 27746 24274 27758
rect 24222 27682 24274 27694
rect 25566 27746 25618 27758
rect 25566 27682 25618 27694
rect 26014 27746 26066 27758
rect 32398 27746 32450 27758
rect 32050 27694 32062 27746
rect 32114 27694 32126 27746
rect 26014 27682 26066 27694
rect 32398 27682 32450 27694
rect 35086 27746 35138 27758
rect 35086 27682 35138 27694
rect 35534 27746 35586 27758
rect 39342 27746 39394 27758
rect 41582 27746 41634 27758
rect 36418 27694 36430 27746
rect 36482 27694 36494 27746
rect 39890 27694 39902 27746
rect 39954 27694 39966 27746
rect 35534 27682 35586 27694
rect 39342 27682 39394 27694
rect 41582 27682 41634 27694
rect 45390 27746 45442 27758
rect 45390 27682 45442 27694
rect 46510 27746 46562 27758
rect 55918 27746 55970 27758
rect 49746 27694 49758 27746
rect 49810 27694 49822 27746
rect 46510 27682 46562 27694
rect 55918 27682 55970 27694
rect 57374 27746 57426 27758
rect 59838 27746 59890 27758
rect 59378 27694 59390 27746
rect 59442 27694 59454 27746
rect 57374 27682 57426 27694
rect 59838 27682 59890 27694
rect 60846 27746 60898 27758
rect 72046 27746 72098 27758
rect 69570 27694 69582 27746
rect 69634 27694 69646 27746
rect 60846 27682 60898 27694
rect 72046 27682 72098 27694
rect 74174 27746 74226 27758
rect 74174 27682 74226 27694
rect 74510 27746 74562 27758
rect 77858 27694 77870 27746
rect 77922 27694 77934 27746
rect 74510 27682 74562 27694
rect 17950 27634 18002 27646
rect 17950 27570 18002 27582
rect 23438 27634 23490 27646
rect 23438 27570 23490 27582
rect 23774 27634 23826 27646
rect 23774 27570 23826 27582
rect 30718 27634 30770 27646
rect 30718 27570 30770 27582
rect 41806 27634 41858 27646
rect 58158 27634 58210 27646
rect 50194 27582 50206 27634
rect 50258 27582 50270 27634
rect 52658 27582 52670 27634
rect 52722 27582 52734 27634
rect 55122 27582 55134 27634
rect 55186 27582 55198 27634
rect 41806 27570 41858 27582
rect 58158 27570 58210 27582
rect 58494 27634 58546 27646
rect 58494 27570 58546 27582
rect 59054 27634 59106 27646
rect 77534 27634 77586 27646
rect 60610 27582 60622 27634
rect 60674 27631 60686 27634
rect 60834 27631 60846 27634
rect 60674 27585 60846 27631
rect 60674 27582 60686 27585
rect 60834 27582 60846 27585
rect 60898 27631 60910 27634
rect 61170 27631 61182 27634
rect 60898 27585 61182 27631
rect 60898 27582 60910 27585
rect 61170 27582 61182 27585
rect 61234 27582 61246 27634
rect 59054 27570 59106 27582
rect 77534 27570 77586 27582
rect 1344 27466 78624 27500
rect 1344 27414 10874 27466
rect 10926 27414 10978 27466
rect 11030 27414 11082 27466
rect 11134 27414 30194 27466
rect 30246 27414 30298 27466
rect 30350 27414 30402 27466
rect 30454 27414 49514 27466
rect 49566 27414 49618 27466
rect 49670 27414 49722 27466
rect 49774 27414 68834 27466
rect 68886 27414 68938 27466
rect 68990 27414 69042 27466
rect 69094 27414 78624 27466
rect 1344 27380 78624 27414
rect 10110 27298 10162 27310
rect 18958 27298 19010 27310
rect 16930 27246 16942 27298
rect 16994 27295 17006 27298
rect 17378 27295 17390 27298
rect 16994 27249 17390 27295
rect 16994 27246 17006 27249
rect 17378 27246 17390 27249
rect 17442 27295 17454 27298
rect 17714 27295 17726 27298
rect 17442 27249 17726 27295
rect 17442 27246 17454 27249
rect 17714 27246 17726 27249
rect 17778 27246 17790 27298
rect 10110 27234 10162 27246
rect 18958 27234 19010 27246
rect 28366 27298 28418 27310
rect 39678 27298 39730 27310
rect 36306 27246 36318 27298
rect 36370 27246 36382 27298
rect 28366 27234 28418 27246
rect 39678 27234 39730 27246
rect 45950 27298 46002 27310
rect 45950 27234 46002 27246
rect 48078 27298 48130 27310
rect 48078 27234 48130 27246
rect 48302 27298 48354 27310
rect 48302 27234 48354 27246
rect 48750 27298 48802 27310
rect 48750 27234 48802 27246
rect 54574 27298 54626 27310
rect 54574 27234 54626 27246
rect 54910 27298 54962 27310
rect 54910 27234 54962 27246
rect 56142 27298 56194 27310
rect 56142 27234 56194 27246
rect 56478 27298 56530 27310
rect 56478 27234 56530 27246
rect 57598 27298 57650 27310
rect 57598 27234 57650 27246
rect 62974 27298 63026 27310
rect 62974 27234 63026 27246
rect 63982 27298 64034 27310
rect 63982 27234 64034 27246
rect 65998 27298 66050 27310
rect 65998 27234 66050 27246
rect 66334 27298 66386 27310
rect 77310 27298 77362 27310
rect 73042 27246 73054 27298
rect 73106 27246 73118 27298
rect 76402 27246 76414 27298
rect 76466 27246 76478 27298
rect 66334 27234 66386 27246
rect 77310 27234 77362 27246
rect 4174 27186 4226 27198
rect 4174 27122 4226 27134
rect 4958 27186 5010 27198
rect 4958 27122 5010 27134
rect 5854 27186 5906 27198
rect 9550 27186 9602 27198
rect 28254 27186 28306 27198
rect 8866 27134 8878 27186
rect 8930 27134 8942 27186
rect 23090 27134 23102 27186
rect 23154 27134 23166 27186
rect 5854 27122 5906 27134
rect 9550 27122 9602 27134
rect 28254 27122 28306 27134
rect 30942 27186 30994 27198
rect 30942 27122 30994 27134
rect 31838 27186 31890 27198
rect 31838 27122 31890 27134
rect 34638 27186 34690 27198
rect 39230 27186 39282 27198
rect 35634 27134 35646 27186
rect 35698 27134 35710 27186
rect 34638 27122 34690 27134
rect 39230 27122 39282 27134
rect 42142 27186 42194 27198
rect 42142 27122 42194 27134
rect 44718 27186 44770 27198
rect 44718 27122 44770 27134
rect 57038 27186 57090 27198
rect 74846 27186 74898 27198
rect 58258 27134 58270 27186
rect 58322 27134 58334 27186
rect 57038 27122 57090 27134
rect 74846 27122 74898 27134
rect 78094 27186 78146 27198
rect 78094 27122 78146 27134
rect 4062 27074 4114 27086
rect 3714 27022 3726 27074
rect 3778 27022 3790 27074
rect 4062 27010 4114 27022
rect 5742 27074 5794 27086
rect 10558 27074 10610 27086
rect 6066 27022 6078 27074
rect 6130 27022 6142 27074
rect 10434 27022 10446 27074
rect 10498 27022 10510 27074
rect 5742 27010 5794 27022
rect 10558 27010 10610 27022
rect 11342 27074 11394 27086
rect 11342 27010 11394 27022
rect 14030 27074 14082 27086
rect 14030 27010 14082 27022
rect 14814 27074 14866 27086
rect 14814 27010 14866 27022
rect 17502 27074 17554 27086
rect 17502 27010 17554 27022
rect 19070 27074 19122 27086
rect 19070 27010 19122 27022
rect 19966 27074 20018 27086
rect 24334 27074 24386 27086
rect 23202 27022 23214 27074
rect 23266 27022 23278 27074
rect 23874 27022 23886 27074
rect 23938 27022 23950 27074
rect 19966 27010 20018 27022
rect 24334 27010 24386 27022
rect 25230 27074 25282 27086
rect 25230 27010 25282 27022
rect 26574 27074 26626 27086
rect 32062 27074 32114 27086
rect 27682 27022 27694 27074
rect 27746 27022 27758 27074
rect 26574 27010 26626 27022
rect 32062 27010 32114 27022
rect 34302 27074 34354 27086
rect 34302 27010 34354 27022
rect 34862 27074 34914 27086
rect 38558 27074 38610 27086
rect 41246 27074 41298 27086
rect 44606 27074 44658 27086
rect 35970 27022 35982 27074
rect 36034 27022 36046 27074
rect 39778 27022 39790 27074
rect 39842 27022 39854 27074
rect 40562 27022 40574 27074
rect 40626 27022 40638 27074
rect 44034 27022 44046 27074
rect 44098 27022 44110 27074
rect 34862 27010 34914 27022
rect 38558 27010 38610 27022
rect 41246 27010 41298 27022
rect 44606 27010 44658 27022
rect 45502 27074 45554 27086
rect 48526 27074 48578 27086
rect 45714 27022 45726 27074
rect 45778 27022 45790 27074
rect 46050 27022 46062 27074
rect 46114 27022 46126 27074
rect 45502 27010 45554 27022
rect 48526 27010 48578 27022
rect 48974 27074 49026 27086
rect 53902 27074 53954 27086
rect 49410 27022 49422 27074
rect 49474 27022 49486 27074
rect 48974 27010 49026 27022
rect 53902 27010 53954 27022
rect 57262 27074 57314 27086
rect 63870 27074 63922 27086
rect 58594 27022 58606 27074
rect 58658 27022 58670 27074
rect 57262 27010 57314 27022
rect 63870 27010 63922 27022
rect 64878 27074 64930 27086
rect 64878 27010 64930 27022
rect 68350 27074 68402 27086
rect 68350 27010 68402 27022
rect 69470 27074 69522 27086
rect 71038 27074 71090 27086
rect 71934 27074 71986 27086
rect 69906 27022 69918 27074
rect 69970 27022 69982 27074
rect 71250 27022 71262 27074
rect 71314 27022 71326 27074
rect 69470 27010 69522 27022
rect 71038 27010 71090 27022
rect 71934 27010 71986 27022
rect 72494 27074 72546 27086
rect 72494 27010 72546 27022
rect 72718 27074 72770 27086
rect 75618 27022 75630 27074
rect 75682 27022 75694 27074
rect 77298 27022 77310 27074
rect 77362 27022 77374 27074
rect 72718 27010 72770 27022
rect 8654 26962 8706 26974
rect 8654 26898 8706 26910
rect 8878 26962 8930 26974
rect 8878 26898 8930 26910
rect 9102 26962 9154 26974
rect 9102 26898 9154 26910
rect 10670 26962 10722 26974
rect 10670 26898 10722 26910
rect 11678 26962 11730 26974
rect 11678 26898 11730 26910
rect 13694 26962 13746 26974
rect 13694 26898 13746 26910
rect 14366 26962 14418 26974
rect 14366 26898 14418 26910
rect 15150 26962 15202 26974
rect 15150 26898 15202 26910
rect 16158 26962 16210 26974
rect 16158 26898 16210 26910
rect 16718 26962 16770 26974
rect 16718 26898 16770 26910
rect 17054 26962 17106 26974
rect 17054 26898 17106 26910
rect 18062 26962 18114 26974
rect 18062 26898 18114 26910
rect 20750 26962 20802 26974
rect 20750 26898 20802 26910
rect 22542 26962 22594 26974
rect 22542 26898 22594 26910
rect 22766 26962 22818 26974
rect 22766 26898 22818 26910
rect 24782 26962 24834 26974
rect 24782 26898 24834 26910
rect 26686 26962 26738 26974
rect 26686 26898 26738 26910
rect 27358 26962 27410 26974
rect 27358 26898 27410 26910
rect 28814 26962 28866 26974
rect 28814 26898 28866 26910
rect 31502 26962 31554 26974
rect 31502 26898 31554 26910
rect 31726 26962 31778 26974
rect 31726 26898 31778 26910
rect 32398 26962 32450 26974
rect 32398 26898 32450 26910
rect 34414 26962 34466 26974
rect 52670 26962 52722 26974
rect 39890 26910 39902 26962
rect 39954 26910 39966 26962
rect 34414 26898 34466 26910
rect 52670 26898 52722 26910
rect 54686 26962 54738 26974
rect 54686 26898 54738 26910
rect 56366 26962 56418 26974
rect 56366 26898 56418 26910
rect 59166 26962 59218 26974
rect 59166 26898 59218 26910
rect 61630 26962 61682 26974
rect 61630 26898 61682 26910
rect 63310 26962 63362 26974
rect 63310 26898 63362 26910
rect 65214 26962 65266 26974
rect 65214 26898 65266 26910
rect 65774 26962 65826 26974
rect 65774 26898 65826 26910
rect 70366 26962 70418 26974
rect 70366 26898 70418 26910
rect 74174 26962 74226 26974
rect 74174 26898 74226 26910
rect 74734 26962 74786 26974
rect 74734 26898 74786 26910
rect 75854 26962 75906 26974
rect 75854 26898 75906 26910
rect 75966 26962 76018 26974
rect 75966 26898 76018 26910
rect 77646 26962 77698 26974
rect 77646 26898 77698 26910
rect 7086 26850 7138 26862
rect 7086 26786 7138 26798
rect 8206 26850 8258 26862
rect 8206 26786 8258 26798
rect 10782 26850 10834 26862
rect 10782 26786 10834 26798
rect 11566 26850 11618 26862
rect 11566 26786 11618 26798
rect 12462 26850 12514 26862
rect 12462 26786 12514 26798
rect 12910 26850 12962 26862
rect 12910 26786 12962 26798
rect 14254 26850 14306 26862
rect 14254 26786 14306 26798
rect 15038 26850 15090 26862
rect 15038 26786 15090 26798
rect 15598 26850 15650 26862
rect 15598 26786 15650 26798
rect 18174 26850 18226 26862
rect 18174 26786 18226 26798
rect 18398 26850 18450 26862
rect 18398 26786 18450 26798
rect 18958 26850 19010 26862
rect 18958 26786 19010 26798
rect 19630 26850 19682 26862
rect 19630 26786 19682 26798
rect 19854 26850 19906 26862
rect 19854 26786 19906 26798
rect 21534 26850 21586 26862
rect 21534 26786 21586 26798
rect 21982 26850 22034 26862
rect 21982 26786 22034 26798
rect 22990 26850 23042 26862
rect 22990 26786 23042 26798
rect 26014 26850 26066 26862
rect 26014 26786 26066 26798
rect 26910 26850 26962 26862
rect 26910 26786 26962 26798
rect 27470 26850 27522 26862
rect 27470 26786 27522 26798
rect 33742 26850 33794 26862
rect 33742 26786 33794 26798
rect 39118 26850 39170 26862
rect 39118 26786 39170 26798
rect 41694 26850 41746 26862
rect 41694 26786 41746 26798
rect 46286 26850 46338 26862
rect 46286 26786 46338 26798
rect 49422 26850 49474 26862
rect 49422 26786 49474 26798
rect 52334 26850 52386 26862
rect 52334 26786 52386 26798
rect 53566 26850 53618 26862
rect 53566 26786 53618 26798
rect 53790 26850 53842 26862
rect 53790 26786 53842 26798
rect 54014 26850 54066 26862
rect 54014 26786 54066 26798
rect 61742 26850 61794 26862
rect 61742 26786 61794 26798
rect 61966 26850 62018 26862
rect 61966 26786 62018 26798
rect 63086 26850 63138 26862
rect 63086 26786 63138 26798
rect 63982 26850 64034 26862
rect 63982 26786 64034 26798
rect 65102 26850 65154 26862
rect 65102 26786 65154 26798
rect 68462 26850 68514 26862
rect 68462 26786 68514 26798
rect 68686 26850 68738 26862
rect 68686 26786 68738 26798
rect 74958 26850 75010 26862
rect 74958 26786 75010 26798
rect 1344 26682 78784 26716
rect 1344 26630 20534 26682
rect 20586 26630 20638 26682
rect 20690 26630 20742 26682
rect 20794 26630 39854 26682
rect 39906 26630 39958 26682
rect 40010 26630 40062 26682
rect 40114 26630 59174 26682
rect 59226 26630 59278 26682
rect 59330 26630 59382 26682
rect 59434 26630 78494 26682
rect 78546 26630 78598 26682
rect 78650 26630 78702 26682
rect 78754 26630 78784 26682
rect 1344 26596 78784 26630
rect 5406 26514 5458 26526
rect 5406 26450 5458 26462
rect 6190 26514 6242 26526
rect 6190 26450 6242 26462
rect 6302 26514 6354 26526
rect 6302 26450 6354 26462
rect 7646 26514 7698 26526
rect 7646 26450 7698 26462
rect 8654 26514 8706 26526
rect 8654 26450 8706 26462
rect 10446 26514 10498 26526
rect 10446 26450 10498 26462
rect 12910 26514 12962 26526
rect 12910 26450 12962 26462
rect 13582 26514 13634 26526
rect 13582 26450 13634 26462
rect 13806 26514 13858 26526
rect 22990 26514 23042 26526
rect 19618 26462 19630 26514
rect 19682 26462 19694 26514
rect 13806 26450 13858 26462
rect 22990 26450 23042 26462
rect 24558 26514 24610 26526
rect 24558 26450 24610 26462
rect 25566 26514 25618 26526
rect 43150 26514 43202 26526
rect 45502 26514 45554 26526
rect 49646 26514 49698 26526
rect 36530 26462 36542 26514
rect 36594 26462 36606 26514
rect 45042 26462 45054 26514
rect 45106 26462 45118 26514
rect 48738 26462 48750 26514
rect 48802 26462 48814 26514
rect 25566 26450 25618 26462
rect 43150 26450 43202 26462
rect 45502 26450 45554 26462
rect 49646 26450 49698 26462
rect 57934 26514 57986 26526
rect 57934 26450 57986 26462
rect 65438 26514 65490 26526
rect 65438 26450 65490 26462
rect 69694 26514 69746 26526
rect 69694 26450 69746 26462
rect 69806 26514 69858 26526
rect 69806 26450 69858 26462
rect 70478 26514 70530 26526
rect 70478 26450 70530 26462
rect 74286 26514 74338 26526
rect 74286 26450 74338 26462
rect 6526 26402 6578 26414
rect 6526 26338 6578 26350
rect 7422 26402 7474 26414
rect 7422 26338 7474 26350
rect 7982 26402 8034 26414
rect 7982 26338 8034 26350
rect 8878 26402 8930 26414
rect 8878 26338 8930 26350
rect 12014 26402 12066 26414
rect 12014 26338 12066 26350
rect 13694 26402 13746 26414
rect 13694 26338 13746 26350
rect 16718 26402 16770 26414
rect 16718 26338 16770 26350
rect 16830 26402 16882 26414
rect 20638 26402 20690 26414
rect 18386 26350 18398 26402
rect 18450 26350 18462 26402
rect 16830 26338 16882 26350
rect 20638 26338 20690 26350
rect 28366 26402 28418 26414
rect 28366 26338 28418 26350
rect 31390 26402 31442 26414
rect 31390 26338 31442 26350
rect 35422 26402 35474 26414
rect 35422 26338 35474 26350
rect 38670 26402 38722 26414
rect 38670 26338 38722 26350
rect 41918 26402 41970 26414
rect 41918 26338 41970 26350
rect 43822 26402 43874 26414
rect 43822 26338 43874 26350
rect 43934 26402 43986 26414
rect 43934 26338 43986 26350
rect 49758 26402 49810 26414
rect 49758 26338 49810 26350
rect 50430 26402 50482 26414
rect 50430 26338 50482 26350
rect 60062 26402 60114 26414
rect 60062 26338 60114 26350
rect 63758 26402 63810 26414
rect 63758 26338 63810 26350
rect 65550 26402 65602 26414
rect 65550 26338 65602 26350
rect 67006 26402 67058 26414
rect 67006 26338 67058 26350
rect 67902 26402 67954 26414
rect 67902 26338 67954 26350
rect 70366 26402 70418 26414
rect 70366 26338 70418 26350
rect 73838 26402 73890 26414
rect 73838 26338 73890 26350
rect 4062 26290 4114 26302
rect 2818 26238 2830 26290
rect 2882 26238 2894 26290
rect 4062 26226 4114 26238
rect 4510 26290 4562 26302
rect 4510 26226 4562 26238
rect 4846 26290 4898 26302
rect 4846 26226 4898 26238
rect 5294 26290 5346 26302
rect 5294 26226 5346 26238
rect 5518 26290 5570 26302
rect 5518 26226 5570 26238
rect 6078 26290 6130 26302
rect 6078 26226 6130 26238
rect 7310 26290 7362 26302
rect 7310 26226 7362 26238
rect 8990 26290 9042 26302
rect 8990 26226 9042 26238
rect 10334 26290 10386 26302
rect 10334 26226 10386 26238
rect 10558 26290 10610 26302
rect 10558 26226 10610 26238
rect 11006 26290 11058 26302
rect 11006 26226 11058 26238
rect 11454 26290 11506 26302
rect 13918 26290 13970 26302
rect 15262 26290 15314 26302
rect 11778 26238 11790 26290
rect 11842 26238 11854 26290
rect 14130 26238 14142 26290
rect 14194 26238 14206 26290
rect 14802 26238 14814 26290
rect 14866 26238 14878 26290
rect 11454 26226 11506 26238
rect 13918 26226 13970 26238
rect 15262 26226 15314 26238
rect 17054 26290 17106 26302
rect 20750 26290 20802 26302
rect 19506 26238 19518 26290
rect 19570 26238 19582 26290
rect 17054 26226 17106 26238
rect 20750 26226 20802 26238
rect 23550 26290 23602 26302
rect 23550 26226 23602 26238
rect 27470 26290 27522 26302
rect 29822 26290 29874 26302
rect 32286 26290 32338 26302
rect 27682 26238 27694 26290
rect 27746 26238 27758 26290
rect 30930 26238 30942 26290
rect 30994 26238 31006 26290
rect 31938 26238 31950 26290
rect 32002 26238 32014 26290
rect 27470 26226 27522 26238
rect 29822 26226 29874 26238
rect 32286 26226 32338 26238
rect 32510 26290 32562 26302
rect 36206 26290 36258 26302
rect 41470 26290 41522 26302
rect 34738 26238 34750 26290
rect 34802 26238 34814 26290
rect 38322 26238 38334 26290
rect 38386 26238 38398 26290
rect 39890 26238 39902 26290
rect 39954 26238 39966 26290
rect 32510 26226 32562 26238
rect 36206 26226 36258 26238
rect 41470 26226 41522 26238
rect 42030 26290 42082 26302
rect 42030 26226 42082 26238
rect 42142 26290 42194 26302
rect 42142 26226 42194 26238
rect 44494 26290 44546 26302
rect 44494 26226 44546 26238
rect 50766 26290 50818 26302
rect 50766 26226 50818 26238
rect 52670 26290 52722 26302
rect 53566 26290 53618 26302
rect 57710 26290 57762 26302
rect 61294 26290 61346 26302
rect 62190 26290 62242 26302
rect 53106 26238 53118 26290
rect 53170 26238 53182 26290
rect 57474 26238 57486 26290
rect 57538 26238 57550 26290
rect 58146 26238 58158 26290
rect 58210 26238 58222 26290
rect 61506 26238 61518 26290
rect 61570 26238 61582 26290
rect 52670 26226 52722 26238
rect 53566 26226 53618 26238
rect 57710 26226 57762 26238
rect 61294 26226 61346 26238
rect 62190 26226 62242 26238
rect 62862 26290 62914 26302
rect 69134 26290 69186 26302
rect 63074 26238 63086 26290
rect 63138 26238 63150 26290
rect 62862 26226 62914 26238
rect 69134 26226 69186 26238
rect 69582 26290 69634 26302
rect 72382 26290 72434 26302
rect 71922 26238 71934 26290
rect 71986 26238 71998 26290
rect 69582 26226 69634 26238
rect 72382 26226 72434 26238
rect 74174 26290 74226 26302
rect 74174 26226 74226 26238
rect 74398 26290 74450 26302
rect 76178 26238 76190 26290
rect 76242 26238 76254 26290
rect 77410 26238 77422 26290
rect 77474 26238 77486 26290
rect 74398 26226 74450 26238
rect 3614 26178 3666 26190
rect 1922 26126 1934 26178
rect 1986 26126 1998 26178
rect 3614 26114 3666 26126
rect 9662 26178 9714 26190
rect 9662 26114 9714 26126
rect 11678 26178 11730 26190
rect 11678 26114 11730 26126
rect 12462 26178 12514 26190
rect 12462 26114 12514 26126
rect 15710 26178 15762 26190
rect 15710 26114 15762 26126
rect 16158 26178 16210 26190
rect 16158 26114 16210 26126
rect 17950 26178 18002 26190
rect 17950 26114 18002 26126
rect 21534 26178 21586 26190
rect 21534 26114 21586 26126
rect 21982 26178 22034 26190
rect 21982 26114 22034 26126
rect 22430 26178 22482 26190
rect 22430 26114 22482 26126
rect 24110 26178 24162 26190
rect 24110 26114 24162 26126
rect 29710 26178 29762 26190
rect 32398 26178 32450 26190
rect 30482 26126 30494 26178
rect 30546 26126 30558 26178
rect 29710 26114 29762 26126
rect 32398 26114 32450 26126
rect 33854 26178 33906 26190
rect 35982 26178 36034 26190
rect 40238 26178 40290 26190
rect 34962 26126 34974 26178
rect 35026 26126 35038 26178
rect 39442 26126 39454 26178
rect 39506 26126 39518 26178
rect 33854 26114 33906 26126
rect 35982 26114 36034 26126
rect 40238 26114 40290 26126
rect 48190 26178 48242 26190
rect 48190 26114 48242 26126
rect 56254 26178 56306 26190
rect 56254 26114 56306 26126
rect 56702 26178 56754 26190
rect 58606 26178 58658 26190
rect 57586 26126 57598 26178
rect 57650 26126 57662 26178
rect 56702 26114 56754 26126
rect 58606 26114 58658 26126
rect 59054 26178 59106 26190
rect 59054 26114 59106 26126
rect 60622 26178 60674 26190
rect 60622 26114 60674 26126
rect 64654 26178 64706 26190
rect 64654 26114 64706 26126
rect 65998 26178 66050 26190
rect 77758 26178 77810 26190
rect 68002 26126 68014 26178
rect 68066 26126 68078 26178
rect 75506 26126 75518 26178
rect 75570 26126 75582 26178
rect 77298 26126 77310 26178
rect 77362 26126 77374 26178
rect 65998 26114 66050 26126
rect 77758 26114 77810 26126
rect 3838 26066 3890 26078
rect 3838 26002 3890 26014
rect 20638 26066 20690 26078
rect 38334 26066 38386 26078
rect 21522 26014 21534 26066
rect 21586 26063 21598 26066
rect 21970 26063 21982 26066
rect 21586 26017 21982 26063
rect 21586 26014 21598 26017
rect 21970 26014 21982 26017
rect 22034 26014 22046 26066
rect 20638 26002 20690 26014
rect 38334 26002 38386 26014
rect 43822 26066 43874 26078
rect 43822 26002 43874 26014
rect 44718 26066 44770 26078
rect 44718 26002 44770 26014
rect 48414 26066 48466 26078
rect 48414 26002 48466 26014
rect 49534 26066 49586 26078
rect 49534 26002 49586 26014
rect 66782 26066 66834 26078
rect 66782 26002 66834 26014
rect 67118 26066 67170 26078
rect 67118 26002 67170 26014
rect 67678 26066 67730 26078
rect 72258 26014 72270 26066
rect 72322 26014 72334 26066
rect 67678 26002 67730 26014
rect 1344 25898 78624 25932
rect 1344 25846 10874 25898
rect 10926 25846 10978 25898
rect 11030 25846 11082 25898
rect 11134 25846 30194 25898
rect 30246 25846 30298 25898
rect 30350 25846 30402 25898
rect 30454 25846 49514 25898
rect 49566 25846 49618 25898
rect 49670 25846 49722 25898
rect 49774 25846 68834 25898
rect 68886 25846 68938 25898
rect 68990 25846 69042 25898
rect 69094 25846 78624 25898
rect 1344 25812 78624 25846
rect 23662 25730 23714 25742
rect 18274 25678 18286 25730
rect 18338 25678 18350 25730
rect 23662 25666 23714 25678
rect 27470 25730 27522 25742
rect 27470 25666 27522 25678
rect 57150 25730 57202 25742
rect 72382 25730 72434 25742
rect 66770 25678 66782 25730
rect 66834 25678 66846 25730
rect 57150 25666 57202 25678
rect 72382 25666 72434 25678
rect 77310 25730 77362 25742
rect 77310 25666 77362 25678
rect 4398 25618 4450 25630
rect 7086 25618 7138 25630
rect 3266 25566 3278 25618
rect 3330 25566 3342 25618
rect 6178 25566 6190 25618
rect 6242 25566 6254 25618
rect 4398 25554 4450 25566
rect 7086 25554 7138 25566
rect 7758 25618 7810 25630
rect 14702 25618 14754 25630
rect 10322 25566 10334 25618
rect 10386 25566 10398 25618
rect 7758 25554 7810 25566
rect 14702 25554 14754 25566
rect 15150 25618 15202 25630
rect 25678 25618 25730 25630
rect 19282 25566 19294 25618
rect 19346 25566 19358 25618
rect 15150 25554 15202 25566
rect 25678 25554 25730 25566
rect 27694 25618 27746 25630
rect 27694 25554 27746 25566
rect 28030 25618 28082 25630
rect 28030 25554 28082 25566
rect 34750 25618 34802 25630
rect 34750 25554 34802 25566
rect 38670 25618 38722 25630
rect 38670 25554 38722 25566
rect 39118 25618 39170 25630
rect 40798 25618 40850 25630
rect 39778 25566 39790 25618
rect 39842 25566 39854 25618
rect 39118 25554 39170 25566
rect 40798 25554 40850 25566
rect 43374 25618 43426 25630
rect 43374 25554 43426 25566
rect 53454 25618 53506 25630
rect 58382 25618 58434 25630
rect 54226 25566 54238 25618
rect 54290 25566 54302 25618
rect 53454 25554 53506 25566
rect 58382 25554 58434 25566
rect 61294 25618 61346 25630
rect 64206 25618 64258 25630
rect 62738 25566 62750 25618
rect 62802 25566 62814 25618
rect 61294 25554 61346 25566
rect 64206 25554 64258 25566
rect 64654 25618 64706 25630
rect 69806 25618 69858 25630
rect 66098 25566 66110 25618
rect 66162 25566 66174 25618
rect 67778 25566 67790 25618
rect 67842 25566 67854 25618
rect 64654 25554 64706 25566
rect 69806 25554 69858 25566
rect 76526 25618 76578 25630
rect 76526 25554 76578 25566
rect 77422 25618 77474 25630
rect 77422 25554 77474 25566
rect 77870 25618 77922 25630
rect 77870 25554 77922 25566
rect 3726 25506 3778 25518
rect 17950 25506 18002 25518
rect 20190 25506 20242 25518
rect 3154 25454 3166 25506
rect 3218 25454 3230 25506
rect 4610 25454 4622 25506
rect 4674 25454 4686 25506
rect 6626 25454 6638 25506
rect 6690 25454 6702 25506
rect 7970 25454 7982 25506
rect 8034 25454 8046 25506
rect 10770 25454 10782 25506
rect 10834 25454 10846 25506
rect 18386 25454 18398 25506
rect 18450 25454 18462 25506
rect 19394 25454 19406 25506
rect 19458 25454 19470 25506
rect 3726 25442 3778 25454
rect 17950 25442 18002 25454
rect 20190 25442 20242 25454
rect 21982 25506 22034 25518
rect 21982 25442 22034 25454
rect 23438 25506 23490 25518
rect 23438 25442 23490 25454
rect 27022 25506 27074 25518
rect 27022 25442 27074 25454
rect 27918 25506 27970 25518
rect 27918 25442 27970 25454
rect 33854 25506 33906 25518
rect 39902 25506 39954 25518
rect 34290 25454 34302 25506
rect 34354 25454 34366 25506
rect 39666 25454 39678 25506
rect 39730 25454 39742 25506
rect 33854 25442 33906 25454
rect 39902 25442 39954 25454
rect 40126 25506 40178 25518
rect 40126 25442 40178 25454
rect 43486 25506 43538 25518
rect 45838 25506 45890 25518
rect 57822 25506 57874 25518
rect 43810 25454 43822 25506
rect 43874 25454 43886 25506
rect 53890 25454 53902 25506
rect 53954 25454 53966 25506
rect 43486 25442 43538 25454
rect 45838 25442 45890 25454
rect 57822 25442 57874 25454
rect 58046 25506 58098 25518
rect 58046 25442 58098 25454
rect 59054 25506 59106 25518
rect 59054 25442 59106 25454
rect 62414 25506 62466 25518
rect 62414 25442 62466 25454
rect 62638 25506 62690 25518
rect 63310 25506 63362 25518
rect 69246 25506 69298 25518
rect 76414 25506 76466 25518
rect 62850 25454 62862 25506
rect 62914 25454 62926 25506
rect 65986 25454 65998 25506
rect 66050 25454 66062 25506
rect 67666 25454 67678 25506
rect 67730 25454 67742 25506
rect 75842 25454 75854 25506
rect 75906 25454 75918 25506
rect 62638 25442 62690 25454
rect 63310 25442 63362 25454
rect 69246 25442 69298 25454
rect 76414 25442 76466 25454
rect 4286 25394 4338 25406
rect 4286 25330 4338 25342
rect 7646 25394 7698 25406
rect 7646 25330 7698 25342
rect 11230 25394 11282 25406
rect 11230 25330 11282 25342
rect 20414 25394 20466 25406
rect 20414 25330 20466 25342
rect 20526 25394 20578 25406
rect 20526 25330 20578 25342
rect 21870 25394 21922 25406
rect 21870 25330 21922 25342
rect 22318 25394 22370 25406
rect 24558 25394 24610 25406
rect 23986 25342 23998 25394
rect 24050 25342 24062 25394
rect 22318 25330 22370 25342
rect 24558 25330 24610 25342
rect 24894 25394 24946 25406
rect 24894 25330 24946 25342
rect 26238 25394 26290 25406
rect 26238 25330 26290 25342
rect 26686 25394 26738 25406
rect 26686 25330 26738 25342
rect 26798 25394 26850 25406
rect 26798 25330 26850 25342
rect 33070 25394 33122 25406
rect 33070 25330 33122 25342
rect 33182 25394 33234 25406
rect 33182 25330 33234 25342
rect 40350 25394 40402 25406
rect 40350 25330 40402 25342
rect 41246 25394 41298 25406
rect 41246 25330 41298 25342
rect 45502 25394 45554 25406
rect 45502 25330 45554 25342
rect 57038 25394 57090 25406
rect 57038 25330 57090 25342
rect 57150 25394 57202 25406
rect 57150 25330 57202 25342
rect 62190 25394 62242 25406
rect 62190 25330 62242 25342
rect 63870 25394 63922 25406
rect 63870 25330 63922 25342
rect 68574 25394 68626 25406
rect 68574 25330 68626 25342
rect 69918 25394 69970 25406
rect 69918 25330 69970 25342
rect 72494 25394 72546 25406
rect 72494 25330 72546 25342
rect 8654 25282 8706 25294
rect 8654 25218 8706 25230
rect 9214 25282 9266 25294
rect 9214 25218 9266 25230
rect 9774 25282 9826 25294
rect 9774 25218 9826 25230
rect 11790 25282 11842 25294
rect 11790 25218 11842 25230
rect 12126 25282 12178 25294
rect 12126 25218 12178 25230
rect 12574 25282 12626 25294
rect 12574 25218 12626 25230
rect 17390 25282 17442 25294
rect 17390 25218 17442 25230
rect 21758 25282 21810 25294
rect 21758 25218 21810 25230
rect 22094 25282 22146 25294
rect 22094 25218 22146 25230
rect 22878 25282 22930 25294
rect 22878 25218 22930 25230
rect 28142 25282 28194 25294
rect 28142 25218 28194 25230
rect 32846 25282 32898 25294
rect 32846 25218 32898 25230
rect 38110 25282 38162 25294
rect 38110 25218 38162 25230
rect 45614 25282 45666 25294
rect 45614 25218 45666 25230
rect 56478 25282 56530 25294
rect 56478 25218 56530 25230
rect 58270 25282 58322 25294
rect 58270 25218 58322 25230
rect 58494 25282 58546 25294
rect 58494 25218 58546 25230
rect 59502 25282 59554 25294
rect 59502 25218 59554 25230
rect 59950 25282 60002 25294
rect 59950 25218 60002 25230
rect 69694 25282 69746 25294
rect 69694 25218 69746 25230
rect 72382 25282 72434 25294
rect 72382 25218 72434 25230
rect 1344 25114 78784 25148
rect 1344 25062 20534 25114
rect 20586 25062 20638 25114
rect 20690 25062 20742 25114
rect 20794 25062 39854 25114
rect 39906 25062 39958 25114
rect 40010 25062 40062 25114
rect 40114 25062 59174 25114
rect 59226 25062 59278 25114
rect 59330 25062 59382 25114
rect 59434 25062 78494 25114
rect 78546 25062 78598 25114
rect 78650 25062 78702 25114
rect 78754 25062 78784 25114
rect 1344 25028 78784 25062
rect 4286 24946 4338 24958
rect 4286 24882 4338 24894
rect 10446 24946 10498 24958
rect 10446 24882 10498 24894
rect 11454 24946 11506 24958
rect 11454 24882 11506 24894
rect 15934 24946 15986 24958
rect 15934 24882 15986 24894
rect 22654 24946 22706 24958
rect 22654 24882 22706 24894
rect 27582 24946 27634 24958
rect 27582 24882 27634 24894
rect 27694 24946 27746 24958
rect 27694 24882 27746 24894
rect 44494 24946 44546 24958
rect 44494 24882 44546 24894
rect 44606 24946 44658 24958
rect 44606 24882 44658 24894
rect 44942 24946 44994 24958
rect 59054 24946 59106 24958
rect 46834 24894 46846 24946
rect 46898 24894 46910 24946
rect 44942 24882 44994 24894
rect 59054 24882 59106 24894
rect 63422 24946 63474 24958
rect 63422 24882 63474 24894
rect 64542 24946 64594 24958
rect 64542 24882 64594 24894
rect 64766 24946 64818 24958
rect 64766 24882 64818 24894
rect 65550 24946 65602 24958
rect 65550 24882 65602 24894
rect 65774 24946 65826 24958
rect 65774 24882 65826 24894
rect 66670 24946 66722 24958
rect 66670 24882 66722 24894
rect 66782 24946 66834 24958
rect 66782 24882 66834 24894
rect 72270 24946 72322 24958
rect 72270 24882 72322 24894
rect 73278 24946 73330 24958
rect 73278 24882 73330 24894
rect 74958 24946 75010 24958
rect 74958 24882 75010 24894
rect 3614 24834 3666 24846
rect 3614 24770 3666 24782
rect 4398 24834 4450 24846
rect 4398 24770 4450 24782
rect 6414 24834 6466 24846
rect 6414 24770 6466 24782
rect 8094 24834 8146 24846
rect 8094 24770 8146 24782
rect 9886 24834 9938 24846
rect 9886 24770 9938 24782
rect 10670 24834 10722 24846
rect 10670 24770 10722 24782
rect 10782 24834 10834 24846
rect 10782 24770 10834 24782
rect 12014 24834 12066 24846
rect 12014 24770 12066 24782
rect 14254 24834 14306 24846
rect 24446 24834 24498 24846
rect 18610 24782 18622 24834
rect 18674 24782 18686 24834
rect 14254 24770 14306 24782
rect 24446 24770 24498 24782
rect 26126 24834 26178 24846
rect 26126 24770 26178 24782
rect 26686 24834 26738 24846
rect 26686 24770 26738 24782
rect 30942 24834 30994 24846
rect 30942 24770 30994 24782
rect 32734 24834 32786 24846
rect 32734 24770 32786 24782
rect 32846 24834 32898 24846
rect 32846 24770 32898 24782
rect 35422 24834 35474 24846
rect 35422 24770 35474 24782
rect 37774 24834 37826 24846
rect 37774 24770 37826 24782
rect 39454 24834 39506 24846
rect 39454 24770 39506 24782
rect 43486 24834 43538 24846
rect 43486 24770 43538 24782
rect 44046 24834 44098 24846
rect 53342 24834 53394 24846
rect 48066 24782 48078 24834
rect 48130 24782 48142 24834
rect 44046 24770 44098 24782
rect 53342 24770 53394 24782
rect 53902 24834 53954 24846
rect 53902 24770 53954 24782
rect 59278 24834 59330 24846
rect 59278 24770 59330 24782
rect 59390 24834 59442 24846
rect 59390 24770 59442 24782
rect 62414 24834 62466 24846
rect 62414 24770 62466 24782
rect 64430 24834 64482 24846
rect 64430 24770 64482 24782
rect 66558 24834 66610 24846
rect 66558 24770 66610 24782
rect 69022 24834 69074 24846
rect 69022 24770 69074 24782
rect 69806 24834 69858 24846
rect 69806 24770 69858 24782
rect 72046 24834 72098 24846
rect 72046 24770 72098 24782
rect 73502 24834 73554 24846
rect 73502 24770 73554 24782
rect 75182 24834 75234 24846
rect 75182 24770 75234 24782
rect 76862 24834 76914 24846
rect 76862 24770 76914 24782
rect 77534 24834 77586 24846
rect 77534 24770 77586 24782
rect 77646 24834 77698 24846
rect 77646 24770 77698 24782
rect 4062 24722 4114 24734
rect 9662 24722 9714 24734
rect 2930 24670 2942 24722
rect 2994 24670 3006 24722
rect 7074 24670 7086 24722
rect 7138 24670 7150 24722
rect 4062 24658 4114 24670
rect 9662 24658 9714 24670
rect 9998 24722 10050 24734
rect 9998 24658 10050 24670
rect 11566 24722 11618 24734
rect 13582 24722 13634 24734
rect 13010 24670 13022 24722
rect 13074 24670 13086 24722
rect 11566 24658 11618 24670
rect 13582 24658 13634 24670
rect 13694 24722 13746 24734
rect 13694 24658 13746 24670
rect 14366 24722 14418 24734
rect 15822 24722 15874 24734
rect 14914 24670 14926 24722
rect 14978 24670 14990 24722
rect 14366 24658 14418 24670
rect 15822 24658 15874 24670
rect 16046 24722 16098 24734
rect 16046 24658 16098 24670
rect 16494 24722 16546 24734
rect 19854 24722 19906 24734
rect 22766 24722 22818 24734
rect 19170 24670 19182 24722
rect 19234 24670 19246 24722
rect 20290 24670 20302 24722
rect 20354 24670 20366 24722
rect 16494 24658 16546 24670
rect 19854 24658 19906 24670
rect 22766 24658 22818 24670
rect 22990 24722 23042 24734
rect 22990 24658 23042 24670
rect 23102 24722 23154 24734
rect 23102 24658 23154 24670
rect 26350 24722 26402 24734
rect 26350 24658 26402 24670
rect 26574 24722 26626 24734
rect 32510 24722 32562 24734
rect 34526 24722 34578 24734
rect 30482 24670 30494 24722
rect 30546 24670 30558 24722
rect 33842 24670 33854 24722
rect 33906 24670 33918 24722
rect 26574 24658 26626 24670
rect 32510 24658 32562 24670
rect 34526 24658 34578 24670
rect 35310 24722 35362 24734
rect 37662 24722 37714 24734
rect 54014 24722 54066 24734
rect 57710 24722 57762 24734
rect 65438 24722 65490 24734
rect 37090 24670 37102 24722
rect 37154 24670 37166 24722
rect 38882 24670 38894 24722
rect 38946 24670 38958 24722
rect 42578 24670 42590 24722
rect 42642 24670 42654 24722
rect 44258 24670 44270 24722
rect 44322 24670 44334 24722
rect 46946 24670 46958 24722
rect 47010 24670 47022 24722
rect 47842 24670 47854 24722
rect 47906 24670 47918 24722
rect 52546 24670 52558 24722
rect 52610 24670 52622 24722
rect 54338 24670 54350 24722
rect 54402 24670 54414 24722
rect 58034 24670 58046 24722
rect 58098 24670 58110 24722
rect 61842 24670 61854 24722
rect 61906 24670 61918 24722
rect 35310 24658 35362 24670
rect 37662 24658 37714 24670
rect 54014 24658 54066 24670
rect 57710 24658 57762 24670
rect 65438 24658 65490 24670
rect 67790 24722 67842 24734
rect 71374 24722 71426 24734
rect 70690 24670 70702 24722
rect 70754 24670 70766 24722
rect 67790 24658 67842 24670
rect 71374 24658 71426 24670
rect 71934 24722 71986 24734
rect 71934 24658 71986 24670
rect 73614 24722 73666 24734
rect 73614 24658 73666 24670
rect 75294 24722 75346 24734
rect 76290 24670 76302 24722
rect 76354 24670 76366 24722
rect 75294 24658 75346 24670
rect 4846 24610 4898 24622
rect 9102 24610 9154 24622
rect 3154 24558 3166 24610
rect 3218 24558 3230 24610
rect 7298 24558 7310 24610
rect 7362 24558 7374 24610
rect 7970 24558 7982 24610
rect 8034 24558 8046 24610
rect 4846 24546 4898 24558
rect 9102 24546 9154 24558
rect 21534 24610 21586 24622
rect 21534 24546 21586 24558
rect 21982 24610 22034 24622
rect 21982 24546 22034 24558
rect 22878 24610 22930 24622
rect 22878 24546 22930 24558
rect 23998 24610 24050 24622
rect 23998 24546 24050 24558
rect 24894 24610 24946 24622
rect 24894 24546 24946 24558
rect 25566 24610 25618 24622
rect 28254 24610 28306 24622
rect 34638 24610 34690 24622
rect 45390 24610 45442 24622
rect 59950 24610 60002 24622
rect 26674 24558 26686 24610
rect 26738 24558 26750 24610
rect 30034 24558 30046 24610
rect 30098 24558 30110 24610
rect 38770 24558 38782 24610
rect 38834 24558 38846 24610
rect 42690 24558 42702 24610
rect 42754 24558 42766 24610
rect 52434 24558 52446 24610
rect 52498 24558 52510 24610
rect 25566 24546 25618 24558
rect 28254 24546 28306 24558
rect 34638 24546 34690 24558
rect 45390 24546 45442 24558
rect 59950 24546 60002 24558
rect 60286 24610 60338 24622
rect 60286 24546 60338 24558
rect 60734 24610 60786 24622
rect 63870 24610 63922 24622
rect 61730 24558 61742 24610
rect 61794 24558 61806 24610
rect 60734 24546 60786 24558
rect 63870 24546 63922 24558
rect 67342 24610 67394 24622
rect 74062 24610 74114 24622
rect 70578 24558 70590 24610
rect 70642 24558 70654 24610
rect 76402 24558 76414 24610
rect 76466 24558 76478 24610
rect 67342 24546 67394 24558
rect 74062 24546 74114 24558
rect 8318 24498 8370 24510
rect 8318 24434 8370 24446
rect 11454 24498 11506 24510
rect 27806 24498 27858 24510
rect 21522 24446 21534 24498
rect 21586 24495 21598 24498
rect 21746 24495 21758 24498
rect 21586 24449 21758 24495
rect 21586 24446 21598 24449
rect 21746 24446 21758 24449
rect 21810 24495 21822 24498
rect 22306 24495 22318 24498
rect 21810 24449 22318 24495
rect 21810 24446 21822 24449
rect 22306 24446 22318 24449
rect 22370 24446 22382 24498
rect 11454 24434 11506 24446
rect 27806 24434 27858 24446
rect 35422 24498 35474 24510
rect 77534 24498 77586 24510
rect 57922 24446 57934 24498
rect 57986 24446 57998 24498
rect 63858 24446 63870 24498
rect 63922 24495 63934 24498
rect 64194 24495 64206 24498
rect 63922 24449 64206 24495
rect 63922 24446 63934 24449
rect 64194 24446 64206 24449
rect 64258 24446 64270 24498
rect 35422 24434 35474 24446
rect 77534 24434 77586 24446
rect 1344 24330 78624 24364
rect 1344 24278 10874 24330
rect 10926 24278 10978 24330
rect 11030 24278 11082 24330
rect 11134 24278 30194 24330
rect 30246 24278 30298 24330
rect 30350 24278 30402 24330
rect 30454 24278 49514 24330
rect 49566 24278 49618 24330
rect 49670 24278 49722 24330
rect 49774 24278 68834 24330
rect 68886 24278 68938 24330
rect 68990 24278 69042 24330
rect 69094 24278 78624 24330
rect 1344 24244 78624 24278
rect 7310 24162 7362 24174
rect 7310 24098 7362 24110
rect 7422 24162 7474 24174
rect 7422 24098 7474 24110
rect 7646 24162 7698 24174
rect 10110 24162 10162 24174
rect 9090 24110 9102 24162
rect 9154 24159 9166 24162
rect 9538 24159 9550 24162
rect 9154 24113 9550 24159
rect 9154 24110 9166 24113
rect 9538 24110 9550 24113
rect 9602 24159 9614 24162
rect 9874 24159 9886 24162
rect 9602 24113 9886 24159
rect 9602 24110 9614 24113
rect 9874 24110 9886 24113
rect 9938 24110 9950 24162
rect 7646 24098 7698 24110
rect 10110 24098 10162 24110
rect 19294 24162 19346 24174
rect 19294 24098 19346 24110
rect 40462 24162 40514 24174
rect 40462 24098 40514 24110
rect 41022 24162 41074 24174
rect 54002 24110 54014 24162
rect 54066 24110 54078 24162
rect 64418 24110 64430 24162
rect 64482 24159 64494 24162
rect 64754 24159 64766 24162
rect 64482 24113 64766 24159
rect 64482 24110 64494 24113
rect 64754 24110 64766 24113
rect 64818 24159 64830 24162
rect 65090 24159 65102 24162
rect 64818 24113 65102 24159
rect 64818 24110 64830 24113
rect 65090 24110 65102 24113
rect 65154 24110 65166 24162
rect 41022 24098 41074 24110
rect 4398 24050 4450 24062
rect 3938 23998 3950 24050
rect 4002 23998 4014 24050
rect 4398 23986 4450 23998
rect 8430 24050 8482 24062
rect 8430 23986 8482 23998
rect 11790 24050 11842 24062
rect 11790 23986 11842 23998
rect 12238 24050 12290 24062
rect 12238 23986 12290 23998
rect 12910 24050 12962 24062
rect 12910 23986 12962 23998
rect 14478 24050 14530 24062
rect 14478 23986 14530 23998
rect 17726 24050 17778 24062
rect 17726 23986 17778 23998
rect 19518 24050 19570 24062
rect 19518 23986 19570 23998
rect 19854 24050 19906 24062
rect 19854 23986 19906 23998
rect 20862 24050 20914 24062
rect 20862 23986 20914 23998
rect 21870 24050 21922 24062
rect 27246 24050 27298 24062
rect 22978 23998 22990 24050
rect 23042 23998 23054 24050
rect 26002 23998 26014 24050
rect 26066 23998 26078 24050
rect 21870 23986 21922 23998
rect 27246 23986 27298 23998
rect 34078 24050 34130 24062
rect 34078 23986 34130 23998
rect 38110 24050 38162 24062
rect 38110 23986 38162 23998
rect 39566 24050 39618 24062
rect 39566 23986 39618 23998
rect 42030 24050 42082 24062
rect 42030 23986 42082 23998
rect 44718 24050 44770 24062
rect 44718 23986 44770 23998
rect 48414 24050 48466 24062
rect 48414 23986 48466 23998
rect 49310 24050 49362 24062
rect 49310 23986 49362 23998
rect 49758 24050 49810 24062
rect 60398 24050 60450 24062
rect 57922 23998 57934 24050
rect 57986 23998 57998 24050
rect 49758 23986 49810 23998
rect 60398 23986 60450 23998
rect 64766 24050 64818 24062
rect 77310 24050 77362 24062
rect 71810 23998 71822 24050
rect 71874 23998 71886 24050
rect 75506 23998 75518 24050
rect 75570 23998 75582 24050
rect 64766 23986 64818 23998
rect 77310 23986 77362 23998
rect 11118 23938 11170 23950
rect 2818 23886 2830 23938
rect 2882 23886 2894 23938
rect 7858 23886 7870 23938
rect 7922 23886 7934 23938
rect 10546 23886 10558 23938
rect 10610 23886 10622 23938
rect 11118 23874 11170 23886
rect 13694 23938 13746 23950
rect 13694 23874 13746 23886
rect 14030 23938 14082 23950
rect 14030 23874 14082 23886
rect 18622 23938 18674 23950
rect 18622 23874 18674 23886
rect 19742 23938 19794 23950
rect 19742 23874 19794 23886
rect 23102 23938 23154 23950
rect 23102 23874 23154 23886
rect 23326 23938 23378 23950
rect 27470 23938 27522 23950
rect 26114 23886 26126 23938
rect 26178 23886 26190 23938
rect 23326 23874 23378 23886
rect 27470 23874 27522 23886
rect 30606 23938 30658 23950
rect 33966 23938 34018 23950
rect 33618 23886 33630 23938
rect 33682 23886 33694 23938
rect 30606 23874 30658 23886
rect 33966 23874 34018 23886
rect 34638 23938 34690 23950
rect 34638 23874 34690 23886
rect 35422 23938 35474 23950
rect 35422 23874 35474 23886
rect 35758 23938 35810 23950
rect 35758 23874 35810 23886
rect 37998 23938 38050 23950
rect 37998 23874 38050 23886
rect 38782 23938 38834 23950
rect 38782 23874 38834 23886
rect 39118 23938 39170 23950
rect 39118 23874 39170 23886
rect 41918 23938 41970 23950
rect 47518 23938 47570 23950
rect 52782 23938 52834 23950
rect 44258 23886 44270 23938
rect 44322 23886 44334 23938
rect 44482 23886 44494 23938
rect 44546 23886 44558 23938
rect 47730 23886 47742 23938
rect 47794 23886 47806 23938
rect 41918 23874 41970 23886
rect 47518 23874 47570 23886
rect 52782 23874 52834 23886
rect 53454 23938 53506 23950
rect 53454 23874 53506 23886
rect 53678 23938 53730 23950
rect 53678 23874 53730 23886
rect 56814 23938 56866 23950
rect 58382 23938 58434 23950
rect 57810 23886 57822 23938
rect 57874 23886 57886 23938
rect 56814 23874 56866 23886
rect 58382 23874 58434 23886
rect 58942 23938 58994 23950
rect 58942 23874 58994 23886
rect 61742 23938 61794 23950
rect 61742 23874 61794 23886
rect 62078 23938 62130 23950
rect 62078 23874 62130 23886
rect 65326 23938 65378 23950
rect 65326 23874 65378 23886
rect 66334 23938 66386 23950
rect 66334 23874 66386 23886
rect 66670 23938 66722 23950
rect 72146 23886 72158 23938
rect 72210 23886 72222 23938
rect 76178 23886 76190 23938
rect 76242 23886 76254 23938
rect 66670 23874 66722 23886
rect 3614 23826 3666 23838
rect 13918 23826 13970 23838
rect 1922 23774 1934 23826
rect 1986 23774 1998 23826
rect 10658 23774 10670 23826
rect 10722 23774 10734 23826
rect 10994 23774 11006 23826
rect 11058 23774 11070 23826
rect 3614 23762 3666 23774
rect 13918 23762 13970 23774
rect 18286 23826 18338 23838
rect 18286 23762 18338 23774
rect 18398 23826 18450 23838
rect 18398 23762 18450 23774
rect 23550 23826 23602 23838
rect 23550 23762 23602 23774
rect 23998 23826 24050 23838
rect 23998 23762 24050 23774
rect 24894 23826 24946 23838
rect 24894 23762 24946 23774
rect 25454 23826 25506 23838
rect 25454 23762 25506 23774
rect 27918 23826 27970 23838
rect 27918 23762 27970 23774
rect 30270 23826 30322 23838
rect 30270 23762 30322 23774
rect 38894 23826 38946 23838
rect 38894 23762 38946 23774
rect 40126 23826 40178 23838
rect 40126 23762 40178 23774
rect 41134 23826 41186 23838
rect 41134 23762 41186 23774
rect 42366 23826 42418 23838
rect 42366 23762 42418 23774
rect 52446 23826 52498 23838
rect 52446 23762 52498 23774
rect 59054 23826 59106 23838
rect 59054 23762 59106 23774
rect 59726 23826 59778 23838
rect 59726 23762 59778 23774
rect 65438 23826 65490 23838
rect 65438 23762 65490 23774
rect 72606 23826 72658 23838
rect 72606 23762 72658 23774
rect 3838 23714 3890 23726
rect 3838 23650 3890 23662
rect 9214 23714 9266 23726
rect 9214 23650 9266 23662
rect 9662 23714 9714 23726
rect 9662 23650 9714 23662
rect 17278 23714 17330 23726
rect 17278 23650 17330 23662
rect 19966 23714 20018 23726
rect 19966 23650 20018 23662
rect 22318 23714 22370 23726
rect 22318 23650 22370 23662
rect 22990 23714 23042 23726
rect 22990 23650 23042 23662
rect 24446 23714 24498 23726
rect 24446 23650 24498 23662
rect 25678 23714 25730 23726
rect 25678 23650 25730 23662
rect 25902 23714 25954 23726
rect 25902 23650 25954 23662
rect 26798 23714 26850 23726
rect 26798 23650 26850 23662
rect 26910 23714 26962 23726
rect 26910 23650 26962 23662
rect 27022 23714 27074 23726
rect 27022 23650 27074 23662
rect 30382 23714 30434 23726
rect 30382 23650 30434 23662
rect 32622 23714 32674 23726
rect 32622 23650 32674 23662
rect 34750 23714 34802 23726
rect 34750 23650 34802 23662
rect 34974 23714 35026 23726
rect 34974 23650 35026 23662
rect 35534 23714 35586 23726
rect 35534 23650 35586 23662
rect 36878 23714 36930 23726
rect 36878 23650 36930 23662
rect 37774 23714 37826 23726
rect 37774 23650 37826 23662
rect 38222 23714 38274 23726
rect 38222 23650 38274 23662
rect 40350 23714 40402 23726
rect 40350 23650 40402 23662
rect 41246 23714 41298 23726
rect 41246 23650 41298 23662
rect 42142 23714 42194 23726
rect 42142 23650 42194 23662
rect 50990 23714 51042 23726
rect 50990 23650 51042 23662
rect 52558 23714 52610 23726
rect 52558 23650 52610 23662
rect 59278 23714 59330 23726
rect 59278 23650 59330 23662
rect 59838 23714 59890 23726
rect 59838 23650 59890 23662
rect 60062 23714 60114 23726
rect 60062 23650 60114 23662
rect 61854 23714 61906 23726
rect 61854 23650 61906 23662
rect 65662 23714 65714 23726
rect 65662 23650 65714 23662
rect 66446 23714 66498 23726
rect 66446 23650 66498 23662
rect 67006 23714 67058 23726
rect 67006 23650 67058 23662
rect 67454 23714 67506 23726
rect 67454 23650 67506 23662
rect 67902 23714 67954 23726
rect 67902 23650 67954 23662
rect 1344 23546 78784 23580
rect 1344 23494 20534 23546
rect 20586 23494 20638 23546
rect 20690 23494 20742 23546
rect 20794 23494 39854 23546
rect 39906 23494 39958 23546
rect 40010 23494 40062 23546
rect 40114 23494 59174 23546
rect 59226 23494 59278 23546
rect 59330 23494 59382 23546
rect 59434 23494 78494 23546
rect 78546 23494 78598 23546
rect 78650 23494 78702 23546
rect 78754 23494 78784 23546
rect 1344 23460 78784 23494
rect 11342 23378 11394 23390
rect 11342 23314 11394 23326
rect 18062 23378 18114 23390
rect 18062 23314 18114 23326
rect 18510 23378 18562 23390
rect 18510 23314 18562 23326
rect 26798 23378 26850 23390
rect 26798 23314 26850 23326
rect 35086 23378 35138 23390
rect 35086 23314 35138 23326
rect 40462 23378 40514 23390
rect 40462 23314 40514 23326
rect 41694 23378 41746 23390
rect 41694 23314 41746 23326
rect 48078 23378 48130 23390
rect 48078 23314 48130 23326
rect 50094 23378 50146 23390
rect 50094 23314 50146 23326
rect 50318 23378 50370 23390
rect 50318 23314 50370 23326
rect 53454 23378 53506 23390
rect 53454 23314 53506 23326
rect 53566 23378 53618 23390
rect 53566 23314 53618 23326
rect 57598 23378 57650 23390
rect 57598 23314 57650 23326
rect 65326 23378 65378 23390
rect 65326 23314 65378 23326
rect 73502 23378 73554 23390
rect 73502 23314 73554 23326
rect 74846 23378 74898 23390
rect 74846 23314 74898 23326
rect 4286 23266 4338 23278
rect 4286 23202 4338 23214
rect 4510 23266 4562 23278
rect 4510 23202 4562 23214
rect 9886 23266 9938 23278
rect 19070 23266 19122 23278
rect 15026 23214 15038 23266
rect 15090 23214 15102 23266
rect 9886 23202 9938 23214
rect 19070 23202 19122 23214
rect 19182 23266 19234 23278
rect 25902 23266 25954 23278
rect 20066 23214 20078 23266
rect 20130 23214 20142 23266
rect 19182 23202 19234 23214
rect 25902 23202 25954 23214
rect 26462 23266 26514 23278
rect 26462 23202 26514 23214
rect 26574 23266 26626 23278
rect 29822 23266 29874 23278
rect 28242 23214 28254 23266
rect 28306 23214 28318 23266
rect 26574 23202 26626 23214
rect 29822 23202 29874 23214
rect 34638 23266 34690 23278
rect 47182 23266 47234 23278
rect 46162 23214 46174 23266
rect 46226 23214 46238 23266
rect 34638 23202 34690 23214
rect 47182 23202 47234 23214
rect 49870 23266 49922 23278
rect 49870 23202 49922 23214
rect 52894 23266 52946 23278
rect 52894 23202 52946 23214
rect 53678 23266 53730 23278
rect 53678 23202 53730 23214
rect 53790 23266 53842 23278
rect 76414 23266 76466 23278
rect 53890 23214 53902 23266
rect 53954 23214 53966 23266
rect 67442 23214 67454 23266
rect 67506 23214 67518 23266
rect 53790 23202 53842 23214
rect 76414 23202 76466 23214
rect 8206 23154 8258 23166
rect 3490 23102 3502 23154
rect 3554 23102 3566 23154
rect 6962 23102 6974 23154
rect 7026 23102 7038 23154
rect 8206 23090 8258 23102
rect 9774 23154 9826 23166
rect 19406 23154 19458 23166
rect 21310 23154 21362 23166
rect 24110 23154 24162 23166
rect 13458 23102 13470 23154
rect 13522 23102 13534 23154
rect 14802 23102 14814 23154
rect 14866 23102 14878 23154
rect 16594 23102 16606 23154
rect 16658 23102 16670 23154
rect 20290 23102 20302 23154
rect 20354 23102 20366 23154
rect 21634 23102 21646 23154
rect 21698 23102 21710 23154
rect 9774 23090 9826 23102
rect 19406 23090 19458 23102
rect 21310 23090 21362 23102
rect 24110 23090 24162 23102
rect 24670 23154 24722 23166
rect 36766 23154 36818 23166
rect 29138 23102 29150 23154
rect 29202 23102 29214 23154
rect 34066 23102 34078 23154
rect 34130 23102 34142 23154
rect 24670 23090 24722 23102
rect 36766 23090 36818 23102
rect 38670 23154 38722 23166
rect 40238 23154 40290 23166
rect 39554 23102 39566 23154
rect 39618 23102 39630 23154
rect 38670 23090 38722 23102
rect 40238 23090 40290 23102
rect 40574 23154 40626 23166
rect 50990 23154 51042 23166
rect 55582 23154 55634 23166
rect 41906 23102 41918 23154
rect 41970 23102 41982 23154
rect 44706 23102 44718 23154
rect 44770 23102 44782 23154
rect 45490 23102 45502 23154
rect 45554 23102 45566 23154
rect 47842 23102 47854 23154
rect 47906 23102 47918 23154
rect 50530 23102 50542 23154
rect 50594 23102 50606 23154
rect 52434 23102 52446 23154
rect 52498 23102 52510 23154
rect 40574 23090 40626 23102
rect 50990 23090 51042 23102
rect 55582 23090 55634 23102
rect 56142 23154 56194 23166
rect 56142 23090 56194 23102
rect 56702 23154 56754 23166
rect 56702 23090 56754 23102
rect 57486 23154 57538 23166
rect 57486 23090 57538 23102
rect 59950 23154 60002 23166
rect 59950 23090 60002 23102
rect 60062 23154 60114 23166
rect 60062 23090 60114 23102
rect 60174 23154 60226 23166
rect 60622 23154 60674 23166
rect 64094 23154 64146 23166
rect 60274 23102 60286 23154
rect 60338 23102 60350 23154
rect 61394 23102 61406 23154
rect 61458 23102 61470 23154
rect 62738 23102 62750 23154
rect 62802 23102 62814 23154
rect 60174 23090 60226 23102
rect 60622 23090 60674 23102
rect 64094 23090 64146 23102
rect 64654 23154 64706 23166
rect 64654 23090 64706 23102
rect 66110 23154 66162 23166
rect 72158 23154 72210 23166
rect 68562 23102 68574 23154
rect 68626 23102 68638 23154
rect 71250 23102 71262 23154
rect 71314 23102 71326 23154
rect 66110 23090 66162 23102
rect 72158 23090 72210 23102
rect 73390 23154 73442 23166
rect 73390 23090 73442 23102
rect 73614 23154 73666 23166
rect 73938 23102 73950 23154
rect 74002 23102 74014 23154
rect 75730 23102 75742 23154
rect 75794 23102 75806 23154
rect 73614 23090 73666 23102
rect 5070 23042 5122 23054
rect 7758 23042 7810 23054
rect 23550 23042 23602 23054
rect 3378 22990 3390 23042
rect 3442 22990 3454 23042
rect 6402 22990 6414 23042
rect 6466 22990 6478 23042
rect 13010 22990 13022 23042
rect 13074 22990 13086 23042
rect 16370 22990 16382 23042
rect 16434 22990 16446 23042
rect 5070 22978 5122 22990
rect 7758 22978 7810 22990
rect 23550 22978 23602 22990
rect 27806 23042 27858 23054
rect 36206 23042 36258 23054
rect 38110 23042 38162 23054
rect 48638 23042 48690 23054
rect 34178 22990 34190 23042
rect 34242 22990 34254 23042
rect 37202 22990 37214 23042
rect 37266 22990 37278 23042
rect 39442 22990 39454 23042
rect 39506 22990 39518 23042
rect 45602 22990 45614 23042
rect 45666 22990 45678 23042
rect 27806 22978 27858 22990
rect 36206 22978 36258 22990
rect 38110 22978 38162 22990
rect 48638 22978 48690 22990
rect 50206 23042 50258 23054
rect 58158 23042 58210 23054
rect 52546 22990 52558 23042
rect 52610 22990 52622 23042
rect 50206 22978 50258 22990
rect 58158 22978 58210 22990
rect 58718 23042 58770 23054
rect 58718 22978 58770 22990
rect 58942 23042 58994 23054
rect 65886 23042 65938 23054
rect 69246 23042 69298 23054
rect 61282 22990 61294 23042
rect 61346 22990 61358 23042
rect 63522 22990 63534 23042
rect 63586 22990 63598 23042
rect 67106 22990 67118 23042
rect 67170 22990 67182 23042
rect 58942 22978 58994 22990
rect 65886 22978 65938 22990
rect 69246 22978 69298 22990
rect 70590 23042 70642 23054
rect 74734 23042 74786 23054
rect 76862 23042 76914 23054
rect 71362 22990 71374 23042
rect 71426 22990 71438 23042
rect 75618 22990 75630 23042
rect 75682 22990 75694 23042
rect 70590 22978 70642 22990
rect 74734 22978 74786 22990
rect 76862 22978 76914 22990
rect 4622 22930 4674 22942
rect 9886 22930 9938 22942
rect 41582 22930 41634 22942
rect 3154 22878 3166 22930
rect 3218 22878 3230 22930
rect 6626 22878 6638 22930
rect 6690 22878 6702 22930
rect 16034 22878 16046 22930
rect 16098 22878 16110 22930
rect 40786 22878 40798 22930
rect 40850 22927 40862 22930
rect 41010 22927 41022 22930
rect 40850 22881 41022 22927
rect 40850 22878 40862 22881
rect 41010 22878 41022 22881
rect 41074 22878 41086 22930
rect 4622 22866 4674 22878
rect 9886 22866 9938 22878
rect 41582 22866 41634 22878
rect 46958 22930 47010 22942
rect 46958 22866 47010 22878
rect 47294 22930 47346 22942
rect 47294 22866 47346 22878
rect 48190 22930 48242 22942
rect 48190 22866 48242 22878
rect 57598 22930 57650 22942
rect 59266 22878 59278 22930
rect 59330 22878 59342 22930
rect 66434 22878 66446 22930
rect 66498 22878 66510 22930
rect 57598 22866 57650 22878
rect 1344 22762 78624 22796
rect 1344 22710 10874 22762
rect 10926 22710 10978 22762
rect 11030 22710 11082 22762
rect 11134 22710 30194 22762
rect 30246 22710 30298 22762
rect 30350 22710 30402 22762
rect 30454 22710 49514 22762
rect 49566 22710 49618 22762
rect 49670 22710 49722 22762
rect 49774 22710 68834 22762
rect 68886 22710 68938 22762
rect 68990 22710 69042 22762
rect 69094 22710 78624 22762
rect 1344 22676 78624 22710
rect 3502 22594 3554 22606
rect 3502 22530 3554 22542
rect 3838 22594 3890 22606
rect 12574 22594 12626 22606
rect 10098 22542 10110 22594
rect 10162 22542 10174 22594
rect 3838 22530 3890 22542
rect 12574 22530 12626 22542
rect 16494 22594 16546 22606
rect 16494 22530 16546 22542
rect 20638 22594 20690 22606
rect 49534 22594 49586 22606
rect 40114 22542 40126 22594
rect 40178 22542 40190 22594
rect 44482 22542 44494 22594
rect 44546 22542 44558 22594
rect 48066 22542 48078 22594
rect 48130 22542 48142 22594
rect 59490 22542 59502 22594
rect 59554 22591 59566 22594
rect 60274 22591 60286 22594
rect 59554 22545 60286 22591
rect 59554 22542 59566 22545
rect 60274 22542 60286 22545
rect 60338 22542 60350 22594
rect 20638 22530 20690 22542
rect 49534 22530 49586 22542
rect 2494 22482 2546 22494
rect 2494 22418 2546 22430
rect 3054 22482 3106 22494
rect 3054 22418 3106 22430
rect 5630 22482 5682 22494
rect 5630 22418 5682 22430
rect 6190 22482 6242 22494
rect 6190 22418 6242 22430
rect 8542 22482 8594 22494
rect 12126 22482 12178 22494
rect 13806 22482 13858 22494
rect 9426 22430 9438 22482
rect 9490 22430 9502 22482
rect 12898 22430 12910 22482
rect 12962 22430 12974 22482
rect 8542 22418 8594 22430
rect 12126 22418 12178 22430
rect 13806 22418 13858 22430
rect 24222 22482 24274 22494
rect 24222 22418 24274 22430
rect 25790 22482 25842 22494
rect 25790 22418 25842 22430
rect 38558 22482 38610 22494
rect 54910 22482 54962 22494
rect 40786 22430 40798 22482
rect 40850 22430 40862 22482
rect 43810 22430 43822 22482
rect 43874 22430 43886 22482
rect 48178 22430 48190 22482
rect 48242 22430 48254 22482
rect 54338 22430 54350 22482
rect 54402 22430 54414 22482
rect 38558 22418 38610 22430
rect 54910 22418 54962 22430
rect 55918 22482 55970 22494
rect 55918 22418 55970 22430
rect 56926 22482 56978 22494
rect 56926 22418 56978 22430
rect 59838 22482 59890 22494
rect 59838 22418 59890 22430
rect 60622 22482 60674 22494
rect 60622 22418 60674 22430
rect 64206 22482 64258 22494
rect 64206 22418 64258 22430
rect 66894 22482 66946 22494
rect 66894 22418 66946 22430
rect 70590 22482 70642 22494
rect 77422 22482 77474 22494
rect 72482 22430 72494 22482
rect 72546 22430 72558 22482
rect 70590 22418 70642 22430
rect 77422 22418 77474 22430
rect 4622 22370 4674 22382
rect 4622 22306 4674 22318
rect 6526 22370 6578 22382
rect 6526 22306 6578 22318
rect 6862 22370 6914 22382
rect 6862 22306 6914 22318
rect 7646 22370 7698 22382
rect 13694 22370 13746 22382
rect 8082 22318 8094 22370
rect 8146 22318 8158 22370
rect 9314 22318 9326 22370
rect 9378 22318 9390 22370
rect 7646 22306 7698 22318
rect 13694 22306 13746 22318
rect 13918 22370 13970 22382
rect 13918 22306 13970 22318
rect 14366 22370 14418 22382
rect 14366 22306 14418 22318
rect 14702 22370 14754 22382
rect 14702 22306 14754 22318
rect 16382 22370 16434 22382
rect 16382 22306 16434 22318
rect 20190 22370 20242 22382
rect 20190 22306 20242 22318
rect 20414 22370 20466 22382
rect 20414 22306 20466 22318
rect 26686 22370 26738 22382
rect 26686 22306 26738 22318
rect 32062 22370 32114 22382
rect 32958 22370 33010 22382
rect 32498 22318 32510 22370
rect 32562 22318 32574 22370
rect 32062 22306 32114 22318
rect 32958 22306 33010 22318
rect 33406 22370 33458 22382
rect 33406 22306 33458 22318
rect 33854 22370 33906 22382
rect 33854 22306 33906 22318
rect 34078 22370 34130 22382
rect 34078 22306 34130 22318
rect 37662 22370 37714 22382
rect 45502 22370 45554 22382
rect 37874 22318 37886 22370
rect 37938 22318 37950 22370
rect 40898 22318 40910 22370
rect 40962 22318 40974 22370
rect 44258 22318 44270 22370
rect 44322 22318 44334 22370
rect 37662 22306 37714 22318
rect 45502 22306 45554 22318
rect 45726 22370 45778 22382
rect 49422 22370 49474 22382
rect 45938 22318 45950 22370
rect 46002 22318 46014 22370
rect 45726 22306 45778 22318
rect 49422 22306 49474 22318
rect 52670 22370 52722 22382
rect 57822 22370 57874 22382
rect 53890 22318 53902 22370
rect 53954 22318 53966 22370
rect 52670 22306 52722 22318
rect 57822 22306 57874 22318
rect 64766 22370 64818 22382
rect 64766 22306 64818 22318
rect 65102 22370 65154 22382
rect 65102 22306 65154 22318
rect 66670 22370 66722 22382
rect 66670 22306 66722 22318
rect 67342 22370 67394 22382
rect 67342 22306 67394 22318
rect 71150 22370 71202 22382
rect 71150 22306 71202 22318
rect 71486 22370 71538 22382
rect 72942 22370 72994 22382
rect 75630 22370 75682 22382
rect 72258 22318 72270 22370
rect 72322 22318 72334 22370
rect 74386 22318 74398 22370
rect 74450 22318 74462 22370
rect 74610 22318 74622 22370
rect 74674 22318 74686 22370
rect 75842 22318 75854 22370
rect 75906 22318 75918 22370
rect 71486 22306 71538 22318
rect 72942 22306 72994 22318
rect 75630 22306 75682 22318
rect 3726 22258 3778 22270
rect 3726 22194 3778 22206
rect 4510 22258 4562 22270
rect 4510 22194 4562 22206
rect 6750 22258 6802 22270
rect 6750 22194 6802 22206
rect 12798 22258 12850 22270
rect 12798 22194 12850 22206
rect 14926 22258 14978 22270
rect 14926 22194 14978 22206
rect 15038 22258 15090 22270
rect 15038 22194 15090 22206
rect 16494 22258 16546 22270
rect 16494 22194 16546 22206
rect 20078 22258 20130 22270
rect 20078 22194 20130 22206
rect 24782 22258 24834 22270
rect 24782 22194 24834 22206
rect 25230 22258 25282 22270
rect 25230 22194 25282 22206
rect 26350 22258 26402 22270
rect 26350 22194 26402 22206
rect 27694 22258 27746 22270
rect 27694 22194 27746 22206
rect 43038 22258 43090 22270
rect 43038 22194 43090 22206
rect 47854 22258 47906 22270
rect 47854 22194 47906 22206
rect 51438 22258 51490 22270
rect 51438 22194 51490 22206
rect 51774 22258 51826 22270
rect 51774 22194 51826 22206
rect 52334 22258 52386 22270
rect 52334 22194 52386 22206
rect 53454 22258 53506 22270
rect 53454 22194 53506 22206
rect 57486 22258 57538 22270
rect 57486 22194 57538 22206
rect 58270 22258 58322 22270
rect 58270 22194 58322 22206
rect 58606 22258 58658 22270
rect 58606 22194 58658 22206
rect 59054 22258 59106 22270
rect 59054 22194 59106 22206
rect 59166 22258 59218 22270
rect 59166 22194 59218 22206
rect 63758 22258 63810 22270
rect 63758 22194 63810 22206
rect 64878 22258 64930 22270
rect 64878 22194 64930 22206
rect 65550 22258 65602 22270
rect 65550 22194 65602 22206
rect 65662 22258 65714 22270
rect 65662 22194 65714 22206
rect 68350 22258 68402 22270
rect 68350 22194 68402 22206
rect 71262 22258 71314 22270
rect 71262 22194 71314 22206
rect 74846 22258 74898 22270
rect 74846 22194 74898 22206
rect 75406 22258 75458 22270
rect 75406 22194 75458 22206
rect 77534 22258 77586 22270
rect 77534 22194 77586 22206
rect 2158 22146 2210 22158
rect 2158 22082 2210 22094
rect 4286 22146 4338 22158
rect 4286 22082 4338 22094
rect 15486 22146 15538 22158
rect 15486 22082 15538 22094
rect 17166 22146 17218 22158
rect 17166 22082 17218 22094
rect 19966 22146 20018 22158
rect 19966 22082 20018 22094
rect 21870 22146 21922 22158
rect 21870 22082 21922 22094
rect 22318 22146 22370 22158
rect 22318 22082 22370 22094
rect 26462 22146 26514 22158
rect 26462 22082 26514 22094
rect 27358 22146 27410 22158
rect 27358 22082 27410 22094
rect 27582 22146 27634 22158
rect 27582 22082 27634 22094
rect 28142 22146 28194 22158
rect 28142 22082 28194 22094
rect 28590 22146 28642 22158
rect 28590 22082 28642 22094
rect 33966 22146 34018 22158
rect 33966 22082 34018 22094
rect 36430 22146 36482 22158
rect 36430 22082 36482 22094
rect 36766 22146 36818 22158
rect 36766 22082 36818 22094
rect 41582 22146 41634 22158
rect 41582 22082 41634 22094
rect 47294 22146 47346 22158
rect 47294 22082 47346 22094
rect 52446 22146 52498 22158
rect 52446 22082 52498 22094
rect 55470 22146 55522 22158
rect 55470 22082 55522 22094
rect 56478 22146 56530 22158
rect 56478 22082 56530 22094
rect 57598 22146 57650 22158
rect 57598 22082 57650 22094
rect 58382 22146 58434 22158
rect 58382 22082 58434 22094
rect 59390 22146 59442 22158
rect 59390 22082 59442 22094
rect 60174 22146 60226 22158
rect 60174 22082 60226 22094
rect 61294 22146 61346 22158
rect 61294 22082 61346 22094
rect 65886 22146 65938 22158
rect 65886 22082 65938 22094
rect 67118 22146 67170 22158
rect 67118 22082 67170 22094
rect 67230 22146 67282 22158
rect 67230 22082 67282 22094
rect 67902 22146 67954 22158
rect 67902 22082 67954 22094
rect 77310 22146 77362 22158
rect 77310 22082 77362 22094
rect 77758 22146 77810 22158
rect 77758 22082 77810 22094
rect 1344 21978 78784 22012
rect 1344 21926 20534 21978
rect 20586 21926 20638 21978
rect 20690 21926 20742 21978
rect 20794 21926 39854 21978
rect 39906 21926 39958 21978
rect 40010 21926 40062 21978
rect 40114 21926 59174 21978
rect 59226 21926 59278 21978
rect 59330 21926 59382 21978
rect 59434 21926 78494 21978
rect 78546 21926 78598 21978
rect 78650 21926 78702 21978
rect 78754 21926 78784 21978
rect 1344 21892 78784 21926
rect 2718 21810 2770 21822
rect 2718 21746 2770 21758
rect 2942 21810 2994 21822
rect 7758 21810 7810 21822
rect 5506 21758 5518 21810
rect 5570 21758 5582 21810
rect 2942 21746 2994 21758
rect 7758 21746 7810 21758
rect 8990 21810 9042 21822
rect 8990 21746 9042 21758
rect 9774 21810 9826 21822
rect 9774 21746 9826 21758
rect 10222 21810 10274 21822
rect 10222 21746 10274 21758
rect 18286 21810 18338 21822
rect 18286 21746 18338 21758
rect 20638 21810 20690 21822
rect 20638 21746 20690 21758
rect 21198 21810 21250 21822
rect 21198 21746 21250 21758
rect 24446 21810 24498 21822
rect 24446 21746 24498 21758
rect 26238 21810 26290 21822
rect 26238 21746 26290 21758
rect 32958 21810 33010 21822
rect 37998 21810 38050 21822
rect 36642 21758 36654 21810
rect 36706 21758 36718 21810
rect 32958 21746 33010 21758
rect 37998 21746 38050 21758
rect 38446 21810 38498 21822
rect 38446 21746 38498 21758
rect 40350 21810 40402 21822
rect 40350 21746 40402 21758
rect 44494 21810 44546 21822
rect 44494 21746 44546 21758
rect 44830 21810 44882 21822
rect 44830 21746 44882 21758
rect 45390 21810 45442 21822
rect 45390 21746 45442 21758
rect 47854 21810 47906 21822
rect 47854 21746 47906 21758
rect 48078 21810 48130 21822
rect 48078 21746 48130 21758
rect 49982 21810 50034 21822
rect 49982 21746 50034 21758
rect 54238 21810 54290 21822
rect 54238 21746 54290 21758
rect 56366 21810 56418 21822
rect 56366 21746 56418 21758
rect 57822 21810 57874 21822
rect 57822 21746 57874 21758
rect 59502 21810 59554 21822
rect 59502 21746 59554 21758
rect 63198 21810 63250 21822
rect 63198 21746 63250 21758
rect 63758 21810 63810 21822
rect 63758 21746 63810 21758
rect 65774 21810 65826 21822
rect 65774 21746 65826 21758
rect 76862 21810 76914 21822
rect 76862 21746 76914 21758
rect 77086 21810 77138 21822
rect 77086 21746 77138 21758
rect 2606 21698 2658 21710
rect 6974 21698 7026 21710
rect 4050 21646 4062 21698
rect 4114 21646 4126 21698
rect 5394 21646 5406 21698
rect 5458 21646 5470 21698
rect 2606 21634 2658 21646
rect 6974 21634 7026 21646
rect 7198 21698 7250 21710
rect 7198 21634 7250 21646
rect 8206 21698 8258 21710
rect 8206 21634 8258 21646
rect 8878 21698 8930 21710
rect 8878 21634 8930 21646
rect 12574 21698 12626 21710
rect 12574 21634 12626 21646
rect 16830 21698 16882 21710
rect 16830 21634 16882 21646
rect 18174 21698 18226 21710
rect 18174 21634 18226 21646
rect 21422 21698 21474 21710
rect 21422 21634 21474 21646
rect 22094 21698 22146 21710
rect 22094 21634 22146 21646
rect 23662 21698 23714 21710
rect 23662 21634 23714 21646
rect 25678 21698 25730 21710
rect 25678 21634 25730 21646
rect 29710 21698 29762 21710
rect 29710 21634 29762 21646
rect 31950 21698 32002 21710
rect 31950 21634 32002 21646
rect 32734 21698 32786 21710
rect 37886 21698 37938 21710
rect 35746 21646 35758 21698
rect 35810 21646 35822 21698
rect 32734 21634 32786 21646
rect 37886 21634 37938 21646
rect 40126 21698 40178 21710
rect 40126 21634 40178 21646
rect 42478 21698 42530 21710
rect 42478 21634 42530 21646
rect 44270 21698 44322 21710
rect 44270 21634 44322 21646
rect 48638 21698 48690 21710
rect 48638 21634 48690 21646
rect 53566 21698 53618 21710
rect 53566 21634 53618 21646
rect 60510 21698 60562 21710
rect 60510 21634 60562 21646
rect 61518 21698 61570 21710
rect 61518 21634 61570 21646
rect 65550 21698 65602 21710
rect 65550 21634 65602 21646
rect 71710 21698 71762 21710
rect 71710 21634 71762 21646
rect 76750 21698 76802 21710
rect 76750 21634 76802 21646
rect 6638 21586 6690 21598
rect 4274 21534 4286 21586
rect 4338 21534 4350 21586
rect 6638 21522 6690 21534
rect 7310 21586 7362 21598
rect 7310 21522 7362 21534
rect 9998 21586 10050 21598
rect 16718 21586 16770 21598
rect 13010 21534 13022 21586
rect 13074 21534 13086 21586
rect 9998 21522 10050 21534
rect 16718 21522 16770 21534
rect 17054 21586 17106 21598
rect 18398 21586 18450 21598
rect 18050 21534 18062 21586
rect 18114 21534 18126 21586
rect 17054 21522 17106 21534
rect 18398 21522 18450 21534
rect 19518 21586 19570 21598
rect 19518 21522 19570 21534
rect 20750 21586 20802 21598
rect 20750 21522 20802 21534
rect 21534 21586 21586 21598
rect 21534 21522 21586 21534
rect 24894 21586 24946 21598
rect 24894 21522 24946 21534
rect 25902 21586 25954 21598
rect 25902 21522 25954 21534
rect 26126 21586 26178 21598
rect 32062 21586 32114 21598
rect 27570 21534 27582 21586
rect 27634 21534 27646 21586
rect 29138 21534 29150 21586
rect 29202 21534 29214 21586
rect 26126 21522 26178 21534
rect 32062 21522 32114 21534
rect 32622 21586 32674 21598
rect 37326 21586 37378 21598
rect 36082 21534 36094 21586
rect 36146 21534 36158 21586
rect 36642 21534 36654 21586
rect 36706 21534 36718 21586
rect 32622 21522 32674 21534
rect 37326 21522 37378 21534
rect 37774 21586 37826 21598
rect 37774 21522 37826 21534
rect 40014 21586 40066 21598
rect 40014 21522 40066 21534
rect 42142 21586 42194 21598
rect 42142 21522 42194 21534
rect 44158 21586 44210 21598
rect 44158 21522 44210 21534
rect 47742 21586 47794 21598
rect 47742 21522 47794 21534
rect 48526 21586 48578 21598
rect 48526 21522 48578 21534
rect 48862 21586 48914 21598
rect 48862 21522 48914 21534
rect 49422 21586 49474 21598
rect 49422 21522 49474 21534
rect 49870 21586 49922 21598
rect 49870 21522 49922 21534
rect 50094 21586 50146 21598
rect 50094 21522 50146 21534
rect 55918 21586 55970 21598
rect 59054 21586 59106 21598
rect 61294 21586 61346 21598
rect 58034 21534 58046 21586
rect 58098 21534 58110 21586
rect 60722 21534 60734 21586
rect 60786 21534 60798 21586
rect 55918 21522 55970 21534
rect 59054 21522 59106 21534
rect 61294 21522 61346 21534
rect 61630 21586 61682 21598
rect 61630 21522 61682 21534
rect 64318 21586 64370 21598
rect 64318 21522 64370 21534
rect 65438 21586 65490 21598
rect 65438 21522 65490 21534
rect 66558 21586 66610 21598
rect 74398 21586 74450 21598
rect 71138 21534 71150 21586
rect 71202 21534 71214 21586
rect 74946 21534 74958 21586
rect 75010 21534 75022 21586
rect 66558 21522 66610 21534
rect 74398 21522 74450 21534
rect 2158 21474 2210 21486
rect 2158 21410 2210 21422
rect 9886 21474 9938 21486
rect 15262 21474 15314 21486
rect 13458 21422 13470 21474
rect 13522 21422 13534 21474
rect 9886 21410 9938 21422
rect 15262 21410 15314 21422
rect 16158 21474 16210 21486
rect 16158 21410 16210 21422
rect 19966 21474 20018 21486
rect 23102 21474 23154 21486
rect 22530 21422 22542 21474
rect 22594 21422 22606 21474
rect 19966 21410 20018 21422
rect 23102 21410 23154 21422
rect 26014 21474 26066 21486
rect 26014 21410 26066 21422
rect 26798 21474 26850 21486
rect 39006 21474 39058 21486
rect 27458 21422 27470 21474
rect 27522 21422 27534 21474
rect 26798 21410 26850 21422
rect 39006 21410 39058 21422
rect 39454 21474 39506 21486
rect 39454 21410 39506 21422
rect 40686 21474 40738 21486
rect 45838 21474 45890 21486
rect 42018 21422 42030 21474
rect 42082 21422 42094 21474
rect 40686 21410 40738 21422
rect 45838 21410 45890 21422
rect 53678 21474 53730 21486
rect 53678 21410 53730 21422
rect 53790 21474 53842 21486
rect 53790 21410 53842 21422
rect 55470 21474 55522 21486
rect 55470 21410 55522 21422
rect 58606 21474 58658 21486
rect 58606 21410 58658 21422
rect 59950 21474 60002 21486
rect 59950 21410 60002 21422
rect 66334 21474 66386 21486
rect 66334 21410 66386 21422
rect 67454 21474 67506 21486
rect 67454 21410 67506 21422
rect 67790 21474 67842 21486
rect 67790 21410 67842 21422
rect 69470 21474 69522 21486
rect 69470 21410 69522 21422
rect 69806 21474 69858 21486
rect 70802 21422 70814 21474
rect 70866 21422 70878 21474
rect 76066 21422 76078 21474
rect 76130 21422 76142 21474
rect 69806 21410 69858 21422
rect 17726 21362 17778 21374
rect 17726 21298 17778 21310
rect 20638 21362 20690 21374
rect 55694 21362 55746 21374
rect 40450 21310 40462 21362
rect 40514 21359 40526 21362
rect 40674 21359 40686 21362
rect 40514 21313 40686 21359
rect 40514 21310 40526 21313
rect 40674 21310 40686 21313
rect 40738 21310 40750 21362
rect 66882 21310 66894 21362
rect 66946 21310 66958 21362
rect 20638 21298 20690 21310
rect 55694 21298 55746 21310
rect 1344 21194 78624 21228
rect 1344 21142 10874 21194
rect 10926 21142 10978 21194
rect 11030 21142 11082 21194
rect 11134 21142 30194 21194
rect 30246 21142 30298 21194
rect 30350 21142 30402 21194
rect 30454 21142 49514 21194
rect 49566 21142 49618 21194
rect 49670 21142 49722 21194
rect 49774 21142 68834 21194
rect 68886 21142 68938 21194
rect 68990 21142 69042 21194
rect 69094 21142 78624 21194
rect 1344 21108 78624 21142
rect 3950 21026 4002 21038
rect 26574 21026 26626 21038
rect 16370 20974 16382 21026
rect 16434 20974 16446 21026
rect 3950 20962 4002 20974
rect 26574 20962 26626 20974
rect 27246 21026 27298 21038
rect 41582 21026 41634 21038
rect 55806 21026 55858 21038
rect 69918 21026 69970 21038
rect 34962 20974 34974 21026
rect 35026 20974 35038 21026
rect 36530 20974 36542 21026
rect 36594 20974 36606 21026
rect 49858 20974 49870 21026
rect 49922 20974 49934 21026
rect 62290 20974 62302 21026
rect 62354 20974 62366 21026
rect 27246 20962 27298 20974
rect 41582 20962 41634 20974
rect 55806 20962 55858 20974
rect 69918 20962 69970 20974
rect 4174 20914 4226 20926
rect 1922 20862 1934 20914
rect 1986 20862 1998 20914
rect 4174 20850 4226 20862
rect 6526 20914 6578 20926
rect 6526 20850 6578 20862
rect 7646 20914 7698 20926
rect 7646 20850 7698 20862
rect 8654 20914 8706 20926
rect 8654 20850 8706 20862
rect 11118 20914 11170 20926
rect 11118 20850 11170 20862
rect 13806 20914 13858 20926
rect 22990 20914 23042 20926
rect 25902 20914 25954 20926
rect 17714 20862 17726 20914
rect 17778 20862 17790 20914
rect 21858 20862 21870 20914
rect 21922 20862 21934 20914
rect 23986 20862 23998 20914
rect 24050 20862 24062 20914
rect 13806 20850 13858 20862
rect 22990 20850 23042 20862
rect 25902 20850 25954 20862
rect 27470 20914 27522 20926
rect 27470 20850 27522 20862
rect 30270 20914 30322 20926
rect 38110 20914 38162 20926
rect 41918 20914 41970 20926
rect 46510 20914 46562 20926
rect 55022 20914 55074 20926
rect 57934 20914 57986 20926
rect 64542 20914 64594 20926
rect 71038 20914 71090 20926
rect 36082 20862 36094 20914
rect 36146 20862 36158 20914
rect 39218 20862 39230 20914
rect 39282 20862 39294 20914
rect 40674 20862 40686 20914
rect 40738 20862 40750 20914
rect 46050 20862 46062 20914
rect 46114 20862 46126 20914
rect 48626 20862 48638 20914
rect 48690 20862 48702 20914
rect 56130 20862 56142 20914
rect 56194 20862 56206 20914
rect 58706 20862 58718 20914
rect 58770 20862 58782 20914
rect 66098 20862 66110 20914
rect 66162 20862 66174 20914
rect 30270 20850 30322 20862
rect 38110 20850 38162 20862
rect 41918 20850 41970 20862
rect 46510 20850 46562 20862
rect 55022 20850 55074 20862
rect 57934 20850 57986 20862
rect 64542 20850 64594 20862
rect 71038 20850 71090 20862
rect 72158 20914 72210 20926
rect 72158 20850 72210 20862
rect 72718 20914 72770 20926
rect 72718 20850 72770 20862
rect 74062 20914 74114 20926
rect 77534 20914 77586 20926
rect 75506 20862 75518 20914
rect 75570 20862 75582 20914
rect 74062 20850 74114 20862
rect 77534 20850 77586 20862
rect 4622 20802 4674 20814
rect 8206 20802 8258 20814
rect 3042 20750 3054 20802
rect 3106 20750 3118 20802
rect 7186 20750 7198 20802
rect 7250 20750 7262 20802
rect 4622 20738 4674 20750
rect 8206 20738 8258 20750
rect 10670 20802 10722 20814
rect 10670 20738 10722 20750
rect 11566 20802 11618 20814
rect 11566 20738 11618 20750
rect 13694 20802 13746 20814
rect 13694 20738 13746 20750
rect 14366 20802 14418 20814
rect 22094 20802 22146 20814
rect 16594 20750 16606 20802
rect 16658 20750 16670 20802
rect 17938 20750 17950 20802
rect 18002 20750 18014 20802
rect 21634 20750 21646 20802
rect 21698 20750 21710 20802
rect 14366 20738 14418 20750
rect 22094 20738 22146 20750
rect 23550 20802 23602 20814
rect 23550 20738 23602 20750
rect 27694 20802 27746 20814
rect 27694 20738 27746 20750
rect 28478 20802 28530 20814
rect 28478 20738 28530 20750
rect 33854 20802 33906 20814
rect 33854 20738 33906 20750
rect 34414 20802 34466 20814
rect 34414 20738 34466 20750
rect 34638 20802 34690 20814
rect 54350 20802 54402 20814
rect 35746 20750 35758 20802
rect 35810 20750 35822 20802
rect 38658 20750 38670 20802
rect 38722 20750 38734 20802
rect 39330 20750 39342 20802
rect 39394 20750 39406 20802
rect 40338 20750 40350 20802
rect 40402 20750 40414 20802
rect 45826 20750 45838 20802
rect 45890 20750 45902 20802
rect 48290 20750 48302 20802
rect 48354 20750 48366 20802
rect 49634 20750 49646 20802
rect 49698 20750 49710 20802
rect 54114 20750 54126 20802
rect 54178 20750 54190 20802
rect 34638 20738 34690 20750
rect 54350 20738 54402 20750
rect 55582 20802 55634 20814
rect 60398 20802 60450 20814
rect 58594 20750 58606 20802
rect 58658 20750 58670 20802
rect 59826 20750 59838 20802
rect 59890 20750 59902 20802
rect 55582 20738 55634 20750
rect 60398 20738 60450 20750
rect 60622 20802 60674 20814
rect 60622 20738 60674 20750
rect 61742 20802 61794 20814
rect 63422 20802 63474 20814
rect 61954 20750 61966 20802
rect 62018 20750 62030 20802
rect 62962 20750 62974 20802
rect 63026 20750 63038 20802
rect 61742 20738 61794 20750
rect 63422 20738 63474 20750
rect 63870 20802 63922 20814
rect 63870 20738 63922 20750
rect 65214 20802 65266 20814
rect 65214 20738 65266 20750
rect 65550 20802 65602 20814
rect 71598 20802 71650 20814
rect 67554 20750 67566 20802
rect 67618 20750 67630 20802
rect 69570 20750 69582 20802
rect 69634 20750 69646 20802
rect 70354 20750 70366 20802
rect 70418 20750 70430 20802
rect 65550 20738 65602 20750
rect 71598 20738 71650 20750
rect 73726 20802 73778 20814
rect 73726 20738 73778 20750
rect 74286 20802 74338 20814
rect 77310 20802 77362 20814
rect 75170 20750 75182 20802
rect 75234 20750 75246 20802
rect 77858 20750 77870 20802
rect 77922 20750 77934 20802
rect 74286 20738 74338 20750
rect 77310 20738 77362 20750
rect 4958 20690 5010 20702
rect 4958 20626 5010 20638
rect 6078 20690 6130 20702
rect 6078 20626 6130 20638
rect 9214 20690 9266 20702
rect 9214 20626 9266 20638
rect 9326 20690 9378 20702
rect 9326 20626 9378 20638
rect 9886 20690 9938 20702
rect 9886 20626 9938 20638
rect 10558 20690 10610 20702
rect 10558 20626 10610 20638
rect 19630 20690 19682 20702
rect 19630 20626 19682 20638
rect 20526 20690 20578 20702
rect 20526 20626 20578 20638
rect 20750 20690 20802 20702
rect 20750 20626 20802 20638
rect 20862 20690 20914 20702
rect 20862 20626 20914 20638
rect 21870 20690 21922 20702
rect 21870 20626 21922 20638
rect 22318 20690 22370 20702
rect 22318 20626 22370 20638
rect 25566 20690 25618 20702
rect 25566 20626 25618 20638
rect 26462 20690 26514 20702
rect 26462 20626 26514 20638
rect 28814 20690 28866 20702
rect 39902 20690 39954 20702
rect 30594 20638 30606 20690
rect 30658 20638 30670 20690
rect 32050 20638 32062 20690
rect 32114 20638 32126 20690
rect 28814 20626 28866 20638
rect 39902 20626 39954 20638
rect 42142 20690 42194 20702
rect 42142 20626 42194 20638
rect 44606 20690 44658 20702
rect 44606 20626 44658 20638
rect 44718 20690 44770 20702
rect 44718 20626 44770 20638
rect 52334 20690 52386 20702
rect 52334 20626 52386 20638
rect 52670 20690 52722 20702
rect 52670 20626 52722 20638
rect 53454 20690 53506 20702
rect 53454 20626 53506 20638
rect 56142 20690 56194 20702
rect 56142 20626 56194 20638
rect 56366 20690 56418 20702
rect 56366 20626 56418 20638
rect 65326 20690 65378 20702
rect 68238 20690 68290 20702
rect 66322 20638 66334 20690
rect 66386 20638 66398 20690
rect 65326 20626 65378 20638
rect 68238 20626 68290 20638
rect 69358 20690 69410 20702
rect 69358 20626 69410 20638
rect 70814 20690 70866 20702
rect 70814 20626 70866 20638
rect 72270 20690 72322 20702
rect 72270 20626 72322 20638
rect 73838 20690 73890 20702
rect 73838 20626 73890 20638
rect 74734 20690 74786 20702
rect 74734 20626 74786 20638
rect 4846 20578 4898 20590
rect 3602 20526 3614 20578
rect 3666 20526 3678 20578
rect 4846 20514 4898 20526
rect 5630 20578 5682 20590
rect 5630 20514 5682 20526
rect 9550 20578 9602 20590
rect 9550 20514 9602 20526
rect 10334 20578 10386 20590
rect 10334 20514 10386 20526
rect 13918 20578 13970 20590
rect 13918 20514 13970 20526
rect 18734 20578 18786 20590
rect 18734 20514 18786 20526
rect 19182 20578 19234 20590
rect 19182 20514 19234 20526
rect 20078 20578 20130 20590
rect 20078 20514 20130 20526
rect 24558 20578 24610 20590
rect 24558 20514 24610 20526
rect 25118 20578 25170 20590
rect 25118 20514 25170 20526
rect 26574 20578 26626 20590
rect 26574 20514 26626 20526
rect 27806 20578 27858 20590
rect 27806 20514 27858 20526
rect 27918 20578 27970 20590
rect 27918 20514 27970 20526
rect 28702 20578 28754 20590
rect 28702 20514 28754 20526
rect 29598 20578 29650 20590
rect 37774 20578 37826 20590
rect 31938 20526 31950 20578
rect 32002 20526 32014 20578
rect 29598 20514 29650 20526
rect 37774 20514 37826 20526
rect 38894 20578 38946 20590
rect 38894 20514 38946 20526
rect 39118 20578 39170 20590
rect 39118 20514 39170 20526
rect 44382 20578 44434 20590
rect 44382 20514 44434 20526
rect 69806 20578 69858 20590
rect 69806 20514 69858 20526
rect 70926 20578 70978 20590
rect 70926 20514 70978 20526
rect 71150 20578 71202 20590
rect 71150 20514 71202 20526
rect 72046 20578 72098 20590
rect 72046 20514 72098 20526
rect 1344 20410 78784 20444
rect 1344 20358 20534 20410
rect 20586 20358 20638 20410
rect 20690 20358 20742 20410
rect 20794 20358 39854 20410
rect 39906 20358 39958 20410
rect 40010 20358 40062 20410
rect 40114 20358 59174 20410
rect 59226 20358 59278 20410
rect 59330 20358 59382 20410
rect 59434 20358 78494 20410
rect 78546 20358 78598 20410
rect 78650 20358 78702 20410
rect 78754 20358 78784 20410
rect 1344 20324 78784 20358
rect 14814 20242 14866 20254
rect 14814 20178 14866 20190
rect 20862 20242 20914 20254
rect 20862 20178 20914 20190
rect 27246 20242 27298 20254
rect 27246 20178 27298 20190
rect 27470 20242 27522 20254
rect 27470 20178 27522 20190
rect 29710 20242 29762 20254
rect 29710 20178 29762 20190
rect 39790 20242 39842 20254
rect 45390 20242 45442 20254
rect 44482 20190 44494 20242
rect 44546 20190 44558 20242
rect 39790 20178 39842 20190
rect 45390 20178 45442 20190
rect 54238 20242 54290 20254
rect 54238 20178 54290 20190
rect 55918 20242 55970 20254
rect 55918 20178 55970 20190
rect 59838 20242 59890 20254
rect 59838 20178 59890 20190
rect 65326 20242 65378 20254
rect 65326 20178 65378 20190
rect 67342 20242 67394 20254
rect 67342 20178 67394 20190
rect 74398 20242 74450 20254
rect 74398 20178 74450 20190
rect 4622 20130 4674 20142
rect 4622 20066 4674 20078
rect 5854 20130 5906 20142
rect 12014 20130 12066 20142
rect 10098 20078 10110 20130
rect 10162 20078 10174 20130
rect 11666 20078 11678 20130
rect 11730 20078 11742 20130
rect 5854 20066 5906 20078
rect 12014 20066 12066 20078
rect 15038 20130 15090 20142
rect 24222 20130 24274 20142
rect 17826 20078 17838 20130
rect 17890 20078 17902 20130
rect 15038 20066 15090 20078
rect 24222 20066 24274 20078
rect 25902 20130 25954 20142
rect 25902 20066 25954 20078
rect 28254 20130 28306 20142
rect 28254 20066 28306 20078
rect 35982 20130 36034 20142
rect 35982 20066 36034 20078
rect 39566 20130 39618 20142
rect 39566 20066 39618 20078
rect 40574 20130 40626 20142
rect 40574 20066 40626 20078
rect 41582 20130 41634 20142
rect 41582 20066 41634 20078
rect 41806 20130 41858 20142
rect 41806 20066 41858 20078
rect 46286 20130 46338 20142
rect 46286 20066 46338 20078
rect 46510 20130 46562 20142
rect 46510 20066 46562 20078
rect 48414 20130 48466 20142
rect 48414 20066 48466 20078
rect 48526 20130 48578 20142
rect 48526 20066 48578 20078
rect 48638 20130 48690 20142
rect 48638 20066 48690 20078
rect 60062 20130 60114 20142
rect 60062 20066 60114 20078
rect 63086 20130 63138 20142
rect 63086 20066 63138 20078
rect 67230 20130 67282 20142
rect 67230 20066 67282 20078
rect 70366 20130 70418 20142
rect 70366 20066 70418 20078
rect 76974 20130 77026 20142
rect 77522 20078 77534 20130
rect 77586 20078 77598 20130
rect 76974 20066 77026 20078
rect 1822 20018 1874 20030
rect 3502 20018 3554 20030
rect 2370 19966 2382 20018
rect 2434 19966 2446 20018
rect 1822 19954 1874 19966
rect 3502 19954 3554 19966
rect 3726 20018 3778 20030
rect 4174 20018 4226 20030
rect 3826 19966 3838 20018
rect 3890 19966 3902 20018
rect 3726 19954 3778 19966
rect 4174 19954 4226 19966
rect 5070 20018 5122 20030
rect 5070 19954 5122 19966
rect 5742 20018 5794 20030
rect 5742 19954 5794 19966
rect 5966 20018 6018 20030
rect 5966 19954 6018 19966
rect 6414 20018 6466 20030
rect 15150 20018 15202 20030
rect 19182 20018 19234 20030
rect 24110 20018 24162 20030
rect 14130 19966 14142 20018
rect 14194 19966 14206 20018
rect 18386 19966 18398 20018
rect 18450 19966 18462 20018
rect 19506 19966 19518 20018
rect 19570 19966 19582 20018
rect 22306 19966 22318 20018
rect 22370 19966 22382 20018
rect 6414 19954 6466 19966
rect 15150 19954 15202 19966
rect 19182 19954 19234 19966
rect 24110 19954 24162 19966
rect 24334 20018 24386 20030
rect 24334 19954 24386 19966
rect 24782 20018 24834 20030
rect 24782 19954 24834 19966
rect 27582 20018 27634 20030
rect 27582 19954 27634 19966
rect 28366 20018 28418 20030
rect 28366 19954 28418 19966
rect 29598 20018 29650 20030
rect 29598 19954 29650 19966
rect 29934 20018 29986 20030
rect 29934 19954 29986 19966
rect 30382 20018 30434 20030
rect 30830 20018 30882 20030
rect 30706 19966 30718 20018
rect 30770 19966 30782 20018
rect 30382 19954 30434 19966
rect 30830 19954 30882 19966
rect 31054 20018 31106 20030
rect 31054 19954 31106 19966
rect 33742 20018 33794 20030
rect 38670 20018 38722 20030
rect 35298 19966 35310 20018
rect 35362 19966 35374 20018
rect 33742 19954 33794 19966
rect 38670 19954 38722 19966
rect 39902 20018 39954 20030
rect 39902 19954 39954 19966
rect 40686 20018 40738 20030
rect 40686 19954 40738 19966
rect 44158 20018 44210 20030
rect 44158 19954 44210 19966
rect 44942 20018 44994 20030
rect 44942 19954 44994 19966
rect 45614 20018 45666 20030
rect 45614 19954 45666 19966
rect 46174 20018 46226 20030
rect 54126 20018 54178 20030
rect 55806 20018 55858 20030
rect 49522 19966 49534 20018
rect 49586 19966 49598 20018
rect 53554 19966 53566 20018
rect 53618 19966 53630 20018
rect 54450 19966 54462 20018
rect 54514 19966 54526 20018
rect 46174 19954 46226 19966
rect 54126 19954 54178 19966
rect 55806 19954 55858 19966
rect 56030 20018 56082 20030
rect 56030 19954 56082 19966
rect 56478 20018 56530 20030
rect 56478 19954 56530 19966
rect 59614 20018 59666 20030
rect 59614 19954 59666 19966
rect 60174 20018 60226 20030
rect 64206 20018 64258 20030
rect 61954 19966 61966 20018
rect 62018 19966 62030 20018
rect 60174 19954 60226 19966
rect 64206 19954 64258 19966
rect 66670 20018 66722 20030
rect 66670 19954 66722 19966
rect 66894 20018 66946 20030
rect 66894 19954 66946 19966
rect 67118 20018 67170 20030
rect 67118 19954 67170 19966
rect 69022 20018 69074 20030
rect 74062 20018 74114 20030
rect 71250 19966 71262 20018
rect 71314 19966 71326 20018
rect 71698 19966 71710 20018
rect 71762 19966 71774 20018
rect 69022 19954 69074 19966
rect 74062 19954 74114 19966
rect 74174 20018 74226 20030
rect 74174 19954 74226 19966
rect 74622 20018 74674 20030
rect 77086 20018 77138 20030
rect 75282 19966 75294 20018
rect 75346 19966 75358 20018
rect 76738 19966 76750 20018
rect 76802 19966 76814 20018
rect 74622 19954 74674 19966
rect 77086 19954 77138 19966
rect 3614 19906 3666 19918
rect 17054 19906 17106 19918
rect 2706 19854 2718 19906
rect 2770 19854 2782 19906
rect 9874 19854 9886 19906
rect 9938 19854 9950 19906
rect 13906 19854 13918 19906
rect 13970 19854 13982 19906
rect 3614 19842 3666 19854
rect 17054 19842 17106 19854
rect 21310 19906 21362 19918
rect 21310 19842 21362 19854
rect 22766 19906 22818 19918
rect 22766 19842 22818 19854
rect 23550 19906 23602 19918
rect 23550 19842 23602 19854
rect 26350 19906 26402 19918
rect 26350 19842 26402 19854
rect 26910 19906 26962 19918
rect 26910 19842 26962 19854
rect 29038 19906 29090 19918
rect 29038 19842 29090 19854
rect 30942 19906 30994 19918
rect 30942 19842 30994 19854
rect 34302 19906 34354 19918
rect 37102 19906 37154 19918
rect 35186 19854 35198 19906
rect 35250 19854 35262 19906
rect 34302 19842 34354 19854
rect 37102 19842 37154 19854
rect 39118 19906 39170 19918
rect 43374 19906 43426 19918
rect 41906 19854 41918 19906
rect 41970 19854 41982 19906
rect 39118 19842 39170 19854
rect 43374 19842 43426 19854
rect 43934 19906 43986 19918
rect 43934 19842 43986 19854
rect 45502 19906 45554 19918
rect 45502 19842 45554 19854
rect 46846 19906 46898 19918
rect 46846 19842 46898 19854
rect 53006 19906 53058 19918
rect 53006 19842 53058 19854
rect 61630 19906 61682 19918
rect 64766 19906 64818 19918
rect 62402 19854 62414 19906
rect 62466 19854 62478 19906
rect 61630 19842 61682 19854
rect 64766 19842 64818 19854
rect 65774 19906 65826 19918
rect 65774 19842 65826 19854
rect 67902 19906 67954 19918
rect 67902 19842 67954 19854
rect 68686 19906 68738 19918
rect 68686 19842 68738 19854
rect 69694 19906 69746 19918
rect 69694 19842 69746 19854
rect 70254 19906 70306 19918
rect 70254 19842 70306 19854
rect 71934 19906 71986 19918
rect 71934 19842 71986 19854
rect 73278 19906 73330 19918
rect 75394 19854 75406 19906
rect 75458 19854 75470 19906
rect 73278 19842 73330 19854
rect 28254 19794 28306 19806
rect 4386 19742 4398 19794
rect 4450 19791 4462 19794
rect 4946 19791 4958 19794
rect 4450 19745 4958 19791
rect 4450 19742 4462 19745
rect 4946 19742 4958 19745
rect 5010 19742 5022 19794
rect 13682 19742 13694 19794
rect 13746 19742 13758 19794
rect 28254 19730 28306 19742
rect 34414 19794 34466 19806
rect 34414 19730 34466 19742
rect 40798 19794 40850 19806
rect 40798 19730 40850 19742
rect 49534 19794 49586 19806
rect 49534 19730 49586 19742
rect 49870 19794 49922 19806
rect 49870 19730 49922 19742
rect 53230 19794 53282 19806
rect 65650 19742 65662 19794
rect 65714 19791 65726 19794
rect 65874 19791 65886 19794
rect 65714 19745 65886 19791
rect 65714 19742 65726 19745
rect 65874 19742 65886 19745
rect 65938 19742 65950 19794
rect 75618 19742 75630 19794
rect 75682 19742 75694 19794
rect 53230 19730 53282 19742
rect 1344 19626 78624 19660
rect 1344 19574 10874 19626
rect 10926 19574 10978 19626
rect 11030 19574 11082 19626
rect 11134 19574 30194 19626
rect 30246 19574 30298 19626
rect 30350 19574 30402 19626
rect 30454 19574 49514 19626
rect 49566 19574 49618 19626
rect 49670 19574 49722 19626
rect 49774 19574 68834 19626
rect 68886 19574 68938 19626
rect 68990 19574 69042 19626
rect 69094 19574 78624 19626
rect 1344 19540 78624 19574
rect 4958 19458 5010 19470
rect 4958 19394 5010 19406
rect 9438 19458 9490 19470
rect 26238 19458 26290 19470
rect 40462 19458 40514 19470
rect 24994 19406 25006 19458
rect 25058 19406 25070 19458
rect 30818 19406 30830 19458
rect 30882 19406 30894 19458
rect 37538 19406 37550 19458
rect 37602 19455 37614 19458
rect 38434 19455 38446 19458
rect 37602 19409 38446 19455
rect 37602 19406 37614 19409
rect 38434 19406 38446 19409
rect 38498 19406 38510 19458
rect 9438 19394 9490 19406
rect 26238 19394 26290 19406
rect 40462 19394 40514 19406
rect 43934 19458 43986 19470
rect 61854 19458 61906 19470
rect 54338 19406 54350 19458
rect 54402 19406 54414 19458
rect 60050 19406 60062 19458
rect 60114 19406 60126 19458
rect 43934 19394 43986 19406
rect 61854 19394 61906 19406
rect 64318 19458 64370 19470
rect 64318 19394 64370 19406
rect 69470 19458 69522 19470
rect 69470 19394 69522 19406
rect 4846 19346 4898 19358
rect 6750 19346 6802 19358
rect 5842 19294 5854 19346
rect 5906 19294 5918 19346
rect 4846 19282 4898 19294
rect 6750 19282 6802 19294
rect 8318 19346 8370 19358
rect 8318 19282 8370 19294
rect 14254 19346 14306 19358
rect 14254 19282 14306 19294
rect 14702 19346 14754 19358
rect 14702 19282 14754 19294
rect 16942 19346 16994 19358
rect 16942 19282 16994 19294
rect 17278 19346 17330 19358
rect 22206 19346 22258 19358
rect 18162 19294 18174 19346
rect 18226 19294 18238 19346
rect 19618 19294 19630 19346
rect 19682 19294 19694 19346
rect 17278 19282 17330 19294
rect 22206 19282 22258 19294
rect 22654 19346 22706 19358
rect 22654 19282 22706 19294
rect 28814 19346 28866 19358
rect 28814 19282 28866 19294
rect 30270 19346 30322 19358
rect 30270 19282 30322 19294
rect 35310 19346 35362 19358
rect 36766 19346 36818 19358
rect 36082 19294 36094 19346
rect 36146 19294 36158 19346
rect 35310 19282 35362 19294
rect 36766 19282 36818 19294
rect 37662 19346 37714 19358
rect 37662 19282 37714 19294
rect 38110 19346 38162 19358
rect 43598 19346 43650 19358
rect 52334 19346 52386 19358
rect 57822 19346 57874 19358
rect 63646 19346 63698 19358
rect 74398 19346 74450 19358
rect 77310 19346 77362 19358
rect 42690 19294 42702 19346
rect 42754 19294 42766 19346
rect 48066 19294 48078 19346
rect 48130 19294 48142 19346
rect 50306 19294 50318 19346
rect 50370 19294 50382 19346
rect 53778 19294 53790 19346
rect 53842 19294 53854 19346
rect 56578 19294 56590 19346
rect 56642 19294 56654 19346
rect 59714 19294 59726 19346
rect 59778 19294 59790 19346
rect 70466 19294 70478 19346
rect 70530 19294 70542 19346
rect 75506 19294 75518 19346
rect 75570 19294 75582 19346
rect 38110 19282 38162 19294
rect 43598 19282 43650 19294
rect 52334 19282 52386 19294
rect 57822 19282 57874 19294
rect 63646 19282 63698 19294
rect 74398 19282 74450 19294
rect 77310 19282 77362 19294
rect 3950 19234 4002 19246
rect 8542 19234 8594 19246
rect 9662 19234 9714 19246
rect 3042 19182 3054 19234
rect 3106 19182 3118 19234
rect 6066 19182 6078 19234
rect 6130 19182 6142 19234
rect 8866 19182 8878 19234
rect 8930 19182 8942 19234
rect 3950 19170 4002 19182
rect 8542 19170 8594 19182
rect 9662 19170 9714 19182
rect 9886 19234 9938 19246
rect 17054 19234 17106 19246
rect 13794 19182 13806 19234
rect 13858 19182 13870 19234
rect 9886 19170 9938 19182
rect 17054 19170 17106 19182
rect 17502 19234 17554 19246
rect 17502 19170 17554 19182
rect 18286 19234 18338 19246
rect 18286 19170 18338 19182
rect 19742 19234 19794 19246
rect 19742 19170 19794 19182
rect 21534 19234 21586 19246
rect 24110 19234 24162 19246
rect 26350 19234 26402 19246
rect 23426 19182 23438 19234
rect 23490 19182 23502 19234
rect 24994 19182 25006 19234
rect 25058 19182 25070 19234
rect 21534 19170 21586 19182
rect 24110 19170 24162 19182
rect 26350 19170 26402 19182
rect 27806 19234 27858 19246
rect 27806 19170 27858 19182
rect 30494 19234 30546 19246
rect 30494 19170 30546 19182
rect 31726 19234 31778 19246
rect 31726 19170 31778 19182
rect 33854 19234 33906 19246
rect 39006 19234 39058 19246
rect 51102 19234 51154 19246
rect 55806 19234 55858 19246
rect 61518 19234 61570 19246
rect 63198 19234 63250 19246
rect 34066 19182 34078 19234
rect 34130 19182 34142 19234
rect 35858 19182 35870 19234
rect 35922 19182 35934 19234
rect 48178 19182 48190 19234
rect 48242 19182 48254 19234
rect 49858 19182 49870 19234
rect 49922 19182 49934 19234
rect 53666 19182 53678 19234
rect 53730 19182 53742 19234
rect 56242 19182 56254 19234
rect 56306 19182 56318 19234
rect 58034 19182 58046 19234
rect 58098 19182 58110 19234
rect 59378 19182 59390 19234
rect 59442 19182 59454 19234
rect 61842 19182 61854 19234
rect 61906 19182 61918 19234
rect 33854 19170 33906 19182
rect 39006 19170 39058 19182
rect 51102 19170 51154 19182
rect 55806 19170 55858 19182
rect 61518 19170 61570 19182
rect 63198 19170 63250 19182
rect 64094 19234 64146 19246
rect 66110 19234 66162 19246
rect 71262 19234 71314 19246
rect 65426 19182 65438 19234
rect 65490 19182 65502 19234
rect 66770 19182 66782 19234
rect 66834 19182 66846 19234
rect 70354 19182 70366 19234
rect 70418 19182 70430 19234
rect 76178 19182 76190 19234
rect 76242 19182 76254 19234
rect 64094 19170 64146 19182
rect 66110 19170 66162 19182
rect 71262 19170 71314 19182
rect 3614 19122 3666 19134
rect 1922 19070 1934 19122
rect 1986 19070 1998 19122
rect 3614 19058 3666 19070
rect 18174 19122 18226 19134
rect 18174 19058 18226 19070
rect 18734 19122 18786 19134
rect 18734 19058 18786 19070
rect 20190 19122 20242 19134
rect 20190 19058 20242 19070
rect 26238 19122 26290 19134
rect 26238 19058 26290 19070
rect 26910 19122 26962 19134
rect 26910 19058 26962 19070
rect 27470 19122 27522 19134
rect 27470 19058 27522 19070
rect 31390 19122 31442 19134
rect 31390 19058 31442 19070
rect 34750 19122 34802 19134
rect 34750 19058 34802 19070
rect 39566 19122 39618 19134
rect 39566 19058 39618 19070
rect 39678 19122 39730 19134
rect 39678 19058 39730 19070
rect 40350 19122 40402 19134
rect 40350 19058 40402 19070
rect 40462 19122 40514 19134
rect 40462 19058 40514 19070
rect 41582 19122 41634 19134
rect 41582 19058 41634 19070
rect 42366 19122 42418 19134
rect 42366 19058 42418 19070
rect 50990 19122 51042 19134
rect 50990 19058 51042 19070
rect 57710 19122 57762 19134
rect 57710 19058 57762 19070
rect 67566 19122 67618 19134
rect 67566 19058 67618 19070
rect 69358 19122 69410 19134
rect 69358 19058 69410 19070
rect 9998 19010 10050 19022
rect 9998 18946 10050 18958
rect 10110 19010 10162 19022
rect 10110 18946 10162 18958
rect 16270 19010 16322 19022
rect 16270 18946 16322 18958
rect 16830 19010 16882 19022
rect 16830 18946 16882 18958
rect 18510 19010 18562 19022
rect 18510 18946 18562 18958
rect 19630 19010 19682 19022
rect 19630 18946 19682 18958
rect 19966 19010 20018 19022
rect 19966 18946 20018 18958
rect 20862 19010 20914 19022
rect 20862 18946 20914 18958
rect 27582 19010 27634 19022
rect 27582 18946 27634 18958
rect 28254 19010 28306 19022
rect 28254 18946 28306 18958
rect 29710 19010 29762 19022
rect 29710 18946 29762 18958
rect 31502 19010 31554 19022
rect 31502 18946 31554 18958
rect 32174 19010 32226 19022
rect 32174 18946 32226 18958
rect 38670 19010 38722 19022
rect 38670 18946 38722 18958
rect 39902 19010 39954 19022
rect 39902 18946 39954 18958
rect 41022 19010 41074 19022
rect 41022 18946 41074 18958
rect 42590 19010 42642 19022
rect 42590 18946 42642 18958
rect 43822 19010 43874 19022
rect 43822 18946 43874 18958
rect 44494 19010 44546 19022
rect 44494 18946 44546 18958
rect 45390 19010 45442 19022
rect 45390 18946 45442 18958
rect 50766 19010 50818 19022
rect 50766 18946 50818 18958
rect 51550 19010 51602 19022
rect 68014 19010 68066 19022
rect 64642 18958 64654 19010
rect 64706 18958 64718 19010
rect 51550 18946 51602 18958
rect 68014 18946 68066 18958
rect 68574 19010 68626 19022
rect 68574 18946 68626 18958
rect 69470 19010 69522 19022
rect 69470 18946 69522 18958
rect 71710 19010 71762 19022
rect 71710 18946 71762 18958
rect 1344 18842 78784 18876
rect 1344 18790 20534 18842
rect 20586 18790 20638 18842
rect 20690 18790 20742 18842
rect 20794 18790 39854 18842
rect 39906 18790 39958 18842
rect 40010 18790 40062 18842
rect 40114 18790 59174 18842
rect 59226 18790 59278 18842
rect 59330 18790 59382 18842
rect 59434 18790 78494 18842
rect 78546 18790 78598 18842
rect 78650 18790 78702 18842
rect 78754 18790 78784 18842
rect 1344 18756 78784 18790
rect 2382 18674 2434 18686
rect 2382 18610 2434 18622
rect 3838 18674 3890 18686
rect 3838 18610 3890 18622
rect 8878 18674 8930 18686
rect 8878 18610 8930 18622
rect 9886 18674 9938 18686
rect 9886 18610 9938 18622
rect 16606 18674 16658 18686
rect 16606 18610 16658 18622
rect 16830 18674 16882 18686
rect 16830 18610 16882 18622
rect 18062 18674 18114 18686
rect 18062 18610 18114 18622
rect 19854 18674 19906 18686
rect 19854 18610 19906 18622
rect 23438 18674 23490 18686
rect 23438 18610 23490 18622
rect 24222 18674 24274 18686
rect 24222 18610 24274 18622
rect 24334 18674 24386 18686
rect 34638 18674 34690 18686
rect 31378 18622 31390 18674
rect 31442 18622 31454 18674
rect 24334 18610 24386 18622
rect 34638 18610 34690 18622
rect 35646 18674 35698 18686
rect 35646 18610 35698 18622
rect 35870 18674 35922 18686
rect 35870 18610 35922 18622
rect 36654 18674 36706 18686
rect 36654 18610 36706 18622
rect 37550 18674 37602 18686
rect 37550 18610 37602 18622
rect 38894 18674 38946 18686
rect 38894 18610 38946 18622
rect 45838 18674 45890 18686
rect 45838 18610 45890 18622
rect 49534 18674 49586 18686
rect 49534 18610 49586 18622
rect 49646 18674 49698 18686
rect 49646 18610 49698 18622
rect 49758 18674 49810 18686
rect 49758 18610 49810 18622
rect 51326 18674 51378 18686
rect 51326 18610 51378 18622
rect 51662 18674 51714 18686
rect 65550 18674 65602 18686
rect 55346 18622 55358 18674
rect 55410 18622 55422 18674
rect 57586 18622 57598 18674
rect 57650 18622 57662 18674
rect 59378 18622 59390 18674
rect 59442 18622 59454 18674
rect 51662 18610 51714 18622
rect 65550 18610 65602 18622
rect 71710 18674 71762 18686
rect 71710 18610 71762 18622
rect 77646 18674 77698 18686
rect 77646 18610 77698 18622
rect 1934 18562 1986 18574
rect 1934 18498 1986 18510
rect 2830 18562 2882 18574
rect 2830 18498 2882 18510
rect 3166 18562 3218 18574
rect 3166 18498 3218 18510
rect 5854 18562 5906 18574
rect 5854 18498 5906 18510
rect 6526 18562 6578 18574
rect 6526 18498 6578 18510
rect 9774 18562 9826 18574
rect 15822 18562 15874 18574
rect 11554 18510 11566 18562
rect 11618 18510 11630 18562
rect 13234 18510 13246 18562
rect 13298 18510 13310 18562
rect 9774 18498 9826 18510
rect 15822 18498 15874 18510
rect 16942 18562 16994 18574
rect 16942 18498 16994 18510
rect 17726 18562 17778 18574
rect 17726 18498 17778 18510
rect 17838 18562 17890 18574
rect 17838 18498 17890 18510
rect 18622 18562 18674 18574
rect 18622 18498 18674 18510
rect 20078 18562 20130 18574
rect 20078 18498 20130 18510
rect 20190 18562 20242 18574
rect 20190 18498 20242 18510
rect 23550 18562 23602 18574
rect 23550 18498 23602 18510
rect 25678 18562 25730 18574
rect 25678 18498 25730 18510
rect 27806 18562 27858 18574
rect 34526 18562 34578 18574
rect 29922 18510 29934 18562
rect 29986 18510 29998 18562
rect 31266 18510 31278 18562
rect 31330 18510 31342 18562
rect 27806 18498 27858 18510
rect 34526 18498 34578 18510
rect 36542 18562 36594 18574
rect 36542 18498 36594 18510
rect 38446 18562 38498 18574
rect 38446 18498 38498 18510
rect 39006 18562 39058 18574
rect 39006 18498 39058 18510
rect 43710 18562 43762 18574
rect 43710 18498 43762 18510
rect 45614 18562 45666 18574
rect 45614 18498 45666 18510
rect 47630 18562 47682 18574
rect 47630 18498 47682 18510
rect 51886 18562 51938 18574
rect 51886 18498 51938 18510
rect 53230 18562 53282 18574
rect 53230 18498 53282 18510
rect 58942 18562 58994 18574
rect 65662 18562 65714 18574
rect 59154 18510 59166 18562
rect 59218 18510 59230 18562
rect 58942 18498 58994 18510
rect 65662 18498 65714 18510
rect 68910 18562 68962 18574
rect 68910 18498 68962 18510
rect 70030 18562 70082 18574
rect 70030 18498 70082 18510
rect 73838 18562 73890 18574
rect 73838 18498 73890 18510
rect 77534 18562 77586 18574
rect 77534 18498 77586 18510
rect 77758 18562 77810 18574
rect 77758 18498 77810 18510
rect 3950 18450 4002 18462
rect 6414 18450 6466 18462
rect 5394 18398 5406 18450
rect 5458 18398 5470 18450
rect 3950 18386 4002 18398
rect 6414 18386 6466 18398
rect 8318 18450 8370 18462
rect 8318 18386 8370 18398
rect 8654 18450 8706 18462
rect 8654 18386 8706 18398
rect 8990 18450 9042 18462
rect 8990 18386 9042 18398
rect 10110 18450 10162 18462
rect 10110 18386 10162 18398
rect 14030 18450 14082 18462
rect 18398 18450 18450 18462
rect 14466 18398 14478 18450
rect 14530 18398 14542 18450
rect 14030 18386 14082 18398
rect 18398 18386 18450 18398
rect 18734 18450 18786 18462
rect 18734 18386 18786 18398
rect 19406 18450 19458 18462
rect 19406 18386 19458 18398
rect 20638 18450 20690 18462
rect 22878 18450 22930 18462
rect 21858 18398 21870 18450
rect 21922 18398 21934 18450
rect 20638 18386 20690 18398
rect 22878 18386 22930 18398
rect 23326 18450 23378 18462
rect 23326 18386 23378 18398
rect 24894 18450 24946 18462
rect 24894 18386 24946 18398
rect 26686 18450 26738 18462
rect 26686 18386 26738 18398
rect 27134 18450 27186 18462
rect 27134 18386 27186 18398
rect 27694 18450 27746 18462
rect 27694 18386 27746 18398
rect 28030 18450 28082 18462
rect 34862 18450 34914 18462
rect 30146 18398 30158 18450
rect 30210 18398 30222 18450
rect 28030 18386 28082 18398
rect 34862 18386 34914 18398
rect 35198 18450 35250 18462
rect 35198 18386 35250 18398
rect 38670 18450 38722 18462
rect 45502 18450 45554 18462
rect 50206 18450 50258 18462
rect 40562 18398 40574 18450
rect 40626 18398 40638 18450
rect 42242 18398 42254 18450
rect 42306 18398 42318 18450
rect 46946 18398 46958 18450
rect 47010 18398 47022 18450
rect 38670 18386 38722 18398
rect 45502 18386 45554 18398
rect 50206 18386 50258 18398
rect 50654 18450 50706 18462
rect 50654 18386 50706 18398
rect 51438 18450 51490 18462
rect 51438 18386 51490 18398
rect 52334 18450 52386 18462
rect 54798 18450 54850 18462
rect 53778 18398 53790 18450
rect 53842 18398 53854 18450
rect 52334 18386 52386 18398
rect 54798 18386 54850 18398
rect 58046 18450 58098 18462
rect 58046 18386 58098 18398
rect 58158 18450 58210 18462
rect 58158 18386 58210 18398
rect 58270 18450 58322 18462
rect 61294 18450 61346 18462
rect 64094 18450 64146 18462
rect 59714 18398 59726 18450
rect 59778 18398 59790 18450
rect 62066 18398 62078 18450
rect 62130 18398 62142 18450
rect 58270 18386 58322 18398
rect 61294 18386 61346 18398
rect 64094 18386 64146 18398
rect 64654 18450 64706 18462
rect 64654 18386 64706 18398
rect 65774 18450 65826 18462
rect 67118 18450 67170 18462
rect 71598 18450 71650 18462
rect 65874 18398 65886 18450
rect 65938 18398 65950 18450
rect 70690 18398 70702 18450
rect 70754 18398 70766 18450
rect 65774 18386 65826 18398
rect 67118 18386 67170 18398
rect 71598 18386 71650 18398
rect 71822 18450 71874 18462
rect 74622 18450 74674 18462
rect 76078 18450 76130 18462
rect 72146 18398 72158 18450
rect 72210 18398 72222 18450
rect 75170 18398 75182 18450
rect 75234 18398 75246 18450
rect 76738 18398 76750 18450
rect 76802 18398 76814 18450
rect 78082 18398 78094 18450
rect 78146 18398 78158 18450
rect 71822 18386 71874 18398
rect 74622 18386 74674 18398
rect 76078 18386 76130 18398
rect 7870 18338 7922 18350
rect 4946 18286 4958 18338
rect 5010 18286 5022 18338
rect 7870 18274 7922 18286
rect 10446 18338 10498 18350
rect 13470 18338 13522 18350
rect 11330 18286 11342 18338
rect 11394 18286 11406 18338
rect 10446 18274 10498 18286
rect 13470 18274 13522 18286
rect 15262 18338 15314 18350
rect 15262 18274 15314 18286
rect 16158 18338 16210 18350
rect 16158 18274 16210 18286
rect 21422 18338 21474 18350
rect 26238 18338 26290 18350
rect 22194 18286 22206 18338
rect 22258 18286 22270 18338
rect 21422 18274 21474 18286
rect 26238 18274 26290 18286
rect 28590 18338 28642 18350
rect 28590 18274 28642 18286
rect 32062 18338 32114 18350
rect 32062 18274 32114 18286
rect 32286 18338 32338 18350
rect 32286 18274 32338 18286
rect 35758 18338 35810 18350
rect 35758 18274 35810 18286
rect 37998 18338 38050 18350
rect 43486 18338 43538 18350
rect 44942 18338 44994 18350
rect 51550 18338 51602 18350
rect 55022 18338 55074 18350
rect 66670 18338 66722 18350
rect 38882 18286 38894 18338
rect 38946 18286 38958 18338
rect 40450 18286 40462 18338
rect 40514 18286 40526 18338
rect 42578 18286 42590 18338
rect 42642 18286 42654 18338
rect 43810 18286 43822 18338
rect 43874 18286 43886 18338
rect 47170 18286 47182 18338
rect 47234 18286 47246 18338
rect 54114 18286 54126 18338
rect 54178 18286 54190 18338
rect 61730 18286 61742 18338
rect 61794 18286 61806 18338
rect 37998 18274 38050 18286
rect 43486 18274 43538 18286
rect 44942 18274 44994 18286
rect 51550 18274 51602 18286
rect 55022 18274 55074 18286
rect 66670 18274 66722 18286
rect 68350 18338 68402 18350
rect 69346 18286 69358 18338
rect 69410 18286 69422 18338
rect 70914 18286 70926 18338
rect 70978 18286 70990 18338
rect 73714 18286 73726 18338
rect 73778 18286 73790 18338
rect 68350 18274 68402 18286
rect 3838 18226 3890 18238
rect 3838 18162 3890 18174
rect 6526 18226 6578 18238
rect 6526 18162 6578 18174
rect 24446 18226 24498 18238
rect 36654 18226 36706 18238
rect 66222 18226 66274 18238
rect 32610 18174 32622 18226
rect 32674 18174 32686 18226
rect 39778 18174 39790 18226
rect 39842 18174 39854 18226
rect 42354 18174 42366 18226
rect 42418 18174 42430 18226
rect 59490 18174 59502 18226
rect 59554 18174 59566 18226
rect 24446 18162 24498 18174
rect 36654 18162 36706 18174
rect 66222 18162 66274 18174
rect 74062 18226 74114 18238
rect 74062 18162 74114 18174
rect 1344 18058 78624 18092
rect 1344 18006 10874 18058
rect 10926 18006 10978 18058
rect 11030 18006 11082 18058
rect 11134 18006 30194 18058
rect 30246 18006 30298 18058
rect 30350 18006 30402 18058
rect 30454 18006 49514 18058
rect 49566 18006 49618 18058
rect 49670 18006 49722 18058
rect 49774 18006 68834 18058
rect 68886 18006 68938 18058
rect 68990 18006 69042 18058
rect 69094 18006 78624 18058
rect 1344 17972 78624 18006
rect 5854 17890 5906 17902
rect 3938 17838 3950 17890
rect 4002 17838 4014 17890
rect 5854 17826 5906 17838
rect 10110 17890 10162 17902
rect 10110 17826 10162 17838
rect 12462 17890 12514 17902
rect 19182 17890 19234 17902
rect 74510 17890 74562 17902
rect 16258 17838 16270 17890
rect 16322 17838 16334 17890
rect 63858 17838 63870 17890
rect 63922 17887 63934 17890
rect 64194 17887 64206 17890
rect 63922 17841 64206 17887
rect 63922 17838 63934 17841
rect 64194 17838 64206 17841
rect 64258 17887 64270 17890
rect 64866 17887 64878 17890
rect 64258 17841 64878 17887
rect 64258 17838 64270 17841
rect 64866 17838 64878 17841
rect 64930 17838 64942 17890
rect 65538 17838 65550 17890
rect 65602 17887 65614 17890
rect 65762 17887 65774 17890
rect 65602 17841 65774 17887
rect 65602 17838 65614 17841
rect 65762 17838 65774 17841
rect 65826 17838 65838 17890
rect 12462 17826 12514 17838
rect 19182 17826 19234 17838
rect 74510 17826 74562 17838
rect 4622 17778 4674 17790
rect 3826 17726 3838 17778
rect 3890 17726 3902 17778
rect 4622 17714 4674 17726
rect 5742 17778 5794 17790
rect 5742 17714 5794 17726
rect 7982 17778 8034 17790
rect 7982 17714 8034 17726
rect 9550 17778 9602 17790
rect 9550 17714 9602 17726
rect 10558 17778 10610 17790
rect 10558 17714 10610 17726
rect 19742 17778 19794 17790
rect 19742 17714 19794 17726
rect 20414 17778 20466 17790
rect 20414 17714 20466 17726
rect 20974 17778 21026 17790
rect 20974 17714 21026 17726
rect 22766 17778 22818 17790
rect 33630 17778 33682 17790
rect 31154 17726 31166 17778
rect 31218 17726 31230 17778
rect 32162 17726 32174 17778
rect 32226 17726 32238 17778
rect 22766 17714 22818 17726
rect 33630 17714 33682 17726
rect 34190 17778 34242 17790
rect 34190 17714 34242 17726
rect 34526 17778 34578 17790
rect 39678 17778 39730 17790
rect 47630 17778 47682 17790
rect 37762 17726 37774 17778
rect 37826 17726 37838 17778
rect 41682 17726 41694 17778
rect 41746 17726 41758 17778
rect 45826 17726 45838 17778
rect 45890 17726 45902 17778
rect 34526 17714 34578 17726
rect 39678 17714 39730 17726
rect 47630 17714 47682 17726
rect 53342 17778 53394 17790
rect 53342 17714 53394 17726
rect 58494 17778 58546 17790
rect 58494 17714 58546 17726
rect 61854 17778 61906 17790
rect 61854 17714 61906 17726
rect 63422 17778 63474 17790
rect 63422 17714 63474 17726
rect 64878 17778 64930 17790
rect 64878 17714 64930 17726
rect 65774 17778 65826 17790
rect 71150 17778 71202 17790
rect 70130 17726 70142 17778
rect 70194 17726 70206 17778
rect 65774 17714 65826 17726
rect 71150 17714 71202 17726
rect 75182 17778 75234 17790
rect 75182 17714 75234 17726
rect 6974 17666 7026 17678
rect 2258 17614 2270 17666
rect 2322 17614 2334 17666
rect 3602 17614 3614 17666
rect 3666 17614 3678 17666
rect 6974 17602 7026 17614
rect 7534 17666 7586 17678
rect 7534 17602 7586 17614
rect 8878 17666 8930 17678
rect 8878 17602 8930 17614
rect 9662 17666 9714 17678
rect 13582 17666 13634 17678
rect 17614 17666 17666 17678
rect 19070 17666 19122 17678
rect 9762 17614 9774 17666
rect 9826 17614 9838 17666
rect 16930 17614 16942 17666
rect 16994 17614 17006 17666
rect 18274 17614 18286 17666
rect 18338 17614 18350 17666
rect 9662 17602 9714 17614
rect 13582 17602 13634 17614
rect 17614 17602 17666 17614
rect 19070 17602 19122 17614
rect 22206 17666 22258 17678
rect 28814 17666 28866 17678
rect 26786 17614 26798 17666
rect 26850 17614 26862 17666
rect 22206 17602 22258 17614
rect 28814 17602 28866 17614
rect 30494 17666 30546 17678
rect 35310 17666 35362 17678
rect 31602 17614 31614 17666
rect 31666 17614 31678 17666
rect 32498 17614 32510 17666
rect 32562 17614 32574 17666
rect 30494 17602 30546 17614
rect 35310 17602 35362 17614
rect 36430 17666 36482 17678
rect 36430 17602 36482 17614
rect 36766 17666 36818 17678
rect 46622 17666 46674 17678
rect 37874 17614 37886 17666
rect 37938 17614 37950 17666
rect 39330 17614 39342 17666
rect 39394 17614 39406 17666
rect 45714 17614 45726 17666
rect 45778 17614 45790 17666
rect 36766 17602 36818 17614
rect 46622 17602 46674 17614
rect 47518 17666 47570 17678
rect 47518 17602 47570 17614
rect 51326 17666 51378 17678
rect 69358 17666 69410 17678
rect 71262 17666 71314 17678
rect 62066 17614 62078 17666
rect 62130 17614 62142 17666
rect 69794 17614 69806 17666
rect 69858 17614 69870 17666
rect 51326 17602 51378 17614
rect 69358 17602 69410 17614
rect 71262 17602 71314 17614
rect 71486 17666 71538 17678
rect 71486 17602 71538 17614
rect 74622 17666 74674 17678
rect 76078 17666 76130 17678
rect 75618 17614 75630 17666
rect 75682 17614 75694 17666
rect 74622 17602 74674 17614
rect 76078 17602 76130 17614
rect 77310 17666 77362 17678
rect 77310 17602 77362 17614
rect 77646 17666 77698 17678
rect 77646 17602 77698 17614
rect 8542 17554 8594 17566
rect 8542 17490 8594 17502
rect 11790 17554 11842 17566
rect 11790 17490 11842 17502
rect 12574 17554 12626 17566
rect 12574 17490 12626 17502
rect 13918 17554 13970 17566
rect 13918 17490 13970 17502
rect 21870 17554 21922 17566
rect 21870 17490 21922 17502
rect 26350 17554 26402 17566
rect 26350 17490 26402 17502
rect 30158 17554 30210 17566
rect 35198 17554 35250 17566
rect 31714 17502 31726 17554
rect 31778 17502 31790 17554
rect 30158 17490 30210 17502
rect 35198 17490 35250 17502
rect 35982 17554 36034 17566
rect 35982 17490 36034 17502
rect 36542 17554 36594 17566
rect 36542 17490 36594 17502
rect 38558 17554 38610 17566
rect 38558 17490 38610 17502
rect 40238 17554 40290 17566
rect 40238 17490 40290 17502
rect 41806 17554 41858 17566
rect 41806 17490 41858 17502
rect 42030 17554 42082 17566
rect 42030 17490 42082 17502
rect 50766 17554 50818 17566
rect 50766 17490 50818 17502
rect 51438 17554 51490 17566
rect 51438 17490 51490 17502
rect 52446 17554 52498 17566
rect 52446 17490 52498 17502
rect 58046 17554 58098 17566
rect 58046 17490 58098 17502
rect 58270 17554 58322 17566
rect 58270 17490 58322 17502
rect 58606 17554 58658 17566
rect 58606 17490 58658 17502
rect 61742 17554 61794 17566
rect 61742 17490 61794 17502
rect 71038 17554 71090 17566
rect 71038 17490 71090 17502
rect 73950 17554 74002 17566
rect 73950 17490 74002 17502
rect 74510 17554 74562 17566
rect 74510 17490 74562 17502
rect 77422 17554 77474 17566
rect 77422 17490 77474 17502
rect 2046 17442 2098 17454
rect 2046 17378 2098 17390
rect 4958 17442 5010 17454
rect 4958 17378 5010 17390
rect 6862 17442 6914 17454
rect 6862 17378 6914 17390
rect 7086 17442 7138 17454
rect 7086 17378 7138 17390
rect 8654 17442 8706 17454
rect 8654 17378 8706 17390
rect 9438 17442 9490 17454
rect 9438 17378 9490 17390
rect 12462 17442 12514 17454
rect 12462 17378 12514 17390
rect 13806 17442 13858 17454
rect 13806 17378 13858 17390
rect 14366 17442 14418 17454
rect 14366 17378 14418 17390
rect 14814 17442 14866 17454
rect 14814 17378 14866 17390
rect 19182 17442 19234 17454
rect 19182 17378 19234 17390
rect 21982 17442 22034 17454
rect 21982 17378 22034 17390
rect 25790 17442 25842 17454
rect 25790 17378 25842 17390
rect 26238 17442 26290 17454
rect 26238 17378 26290 17390
rect 26462 17442 26514 17454
rect 26462 17378 26514 17390
rect 28142 17442 28194 17454
rect 28142 17378 28194 17390
rect 29598 17442 29650 17454
rect 29598 17378 29650 17390
rect 30270 17442 30322 17454
rect 30270 17378 30322 17390
rect 33294 17442 33346 17454
rect 33294 17378 33346 17390
rect 34974 17442 35026 17454
rect 34974 17378 35026 17390
rect 39566 17442 39618 17454
rect 39566 17378 39618 17390
rect 40350 17442 40402 17454
rect 40350 17378 40402 17390
rect 40574 17442 40626 17454
rect 40574 17378 40626 17390
rect 40910 17442 40962 17454
rect 40910 17378 40962 17390
rect 44718 17442 44770 17454
rect 44718 17378 44770 17390
rect 47294 17442 47346 17454
rect 47294 17378 47346 17390
rect 47742 17442 47794 17454
rect 47742 17378 47794 17390
rect 48974 17442 49026 17454
rect 48974 17378 49026 17390
rect 49422 17442 49474 17454
rect 49422 17378 49474 17390
rect 50318 17442 50370 17454
rect 50318 17378 50370 17390
rect 51662 17442 51714 17454
rect 51662 17378 51714 17390
rect 52222 17442 52274 17454
rect 52222 17378 52274 17390
rect 52334 17442 52386 17454
rect 52334 17378 52386 17390
rect 63086 17442 63138 17454
rect 63086 17378 63138 17390
rect 63870 17442 63922 17454
rect 63870 17378 63922 17390
rect 64430 17442 64482 17454
rect 64430 17378 64482 17390
rect 65326 17442 65378 17454
rect 65326 17378 65378 17390
rect 73502 17442 73554 17454
rect 73502 17378 73554 17390
rect 77982 17442 78034 17454
rect 77982 17378 78034 17390
rect 1344 17274 78784 17308
rect 1344 17222 20534 17274
rect 20586 17222 20638 17274
rect 20690 17222 20742 17274
rect 20794 17222 39854 17274
rect 39906 17222 39958 17274
rect 40010 17222 40062 17274
rect 40114 17222 59174 17274
rect 59226 17222 59278 17274
rect 59330 17222 59382 17274
rect 59434 17222 78494 17274
rect 78546 17222 78598 17274
rect 78650 17222 78702 17274
rect 78754 17222 78784 17274
rect 1344 17188 78784 17222
rect 11902 17106 11954 17118
rect 9762 17054 9774 17106
rect 9826 17054 9838 17106
rect 11902 17042 11954 17054
rect 12350 17106 12402 17118
rect 12350 17042 12402 17054
rect 12798 17106 12850 17118
rect 12798 17042 12850 17054
rect 13470 17106 13522 17118
rect 13470 17042 13522 17054
rect 14590 17106 14642 17118
rect 14590 17042 14642 17054
rect 17054 17106 17106 17118
rect 17054 17042 17106 17054
rect 18174 17106 18226 17118
rect 18174 17042 18226 17054
rect 19182 17106 19234 17118
rect 19182 17042 19234 17054
rect 19630 17106 19682 17118
rect 19630 17042 19682 17054
rect 20190 17106 20242 17118
rect 20190 17042 20242 17054
rect 29150 17106 29202 17118
rect 29150 17042 29202 17054
rect 30270 17106 30322 17118
rect 30270 17042 30322 17054
rect 30494 17106 30546 17118
rect 30494 17042 30546 17054
rect 32734 17106 32786 17118
rect 32734 17042 32786 17054
rect 33518 17106 33570 17118
rect 33518 17042 33570 17054
rect 38670 17106 38722 17118
rect 38670 17042 38722 17054
rect 39230 17106 39282 17118
rect 39230 17042 39282 17054
rect 40686 17106 40738 17118
rect 40686 17042 40738 17054
rect 40910 17106 40962 17118
rect 40910 17042 40962 17054
rect 47630 17106 47682 17118
rect 47630 17042 47682 17054
rect 48638 17106 48690 17118
rect 48638 17042 48690 17054
rect 50542 17106 50594 17118
rect 50542 17042 50594 17054
rect 52782 17106 52834 17118
rect 52782 17042 52834 17054
rect 52894 17106 52946 17118
rect 52894 17042 52946 17054
rect 53678 17106 53730 17118
rect 60286 17106 60338 17118
rect 58034 17054 58046 17106
rect 58098 17054 58110 17106
rect 53678 17042 53730 17054
rect 60286 17042 60338 17054
rect 60734 17106 60786 17118
rect 60734 17042 60786 17054
rect 63086 17106 63138 17118
rect 74062 17106 74114 17118
rect 70018 17054 70030 17106
rect 70082 17054 70094 17106
rect 63086 17042 63138 17054
rect 74062 17042 74114 17054
rect 3950 16994 4002 17006
rect 3950 16930 4002 16942
rect 4734 16994 4786 17006
rect 4734 16930 4786 16942
rect 13582 16994 13634 17006
rect 13582 16930 13634 16942
rect 16830 16994 16882 17006
rect 16830 16930 16882 16942
rect 32510 16994 32562 17006
rect 32510 16930 32562 16942
rect 32846 16994 32898 17006
rect 46174 16994 46226 17006
rect 42466 16942 42478 16994
rect 42530 16942 42542 16994
rect 43810 16942 43822 16994
rect 43874 16942 43886 16994
rect 32846 16930 32898 16942
rect 46174 16930 46226 16942
rect 46286 16994 46338 17006
rect 55470 16994 55522 17006
rect 64654 16994 64706 17006
rect 49970 16942 49982 16994
rect 50034 16942 50046 16994
rect 61394 16942 61406 16994
rect 61458 16942 61470 16994
rect 46286 16930 46338 16942
rect 55470 16930 55522 16942
rect 64654 16930 64706 16942
rect 67566 16994 67618 17006
rect 67566 16930 67618 16942
rect 73726 16994 73778 17006
rect 73726 16930 73778 16942
rect 76750 16994 76802 17006
rect 76750 16930 76802 16942
rect 5294 16882 5346 16894
rect 7870 16882 7922 16894
rect 2034 16830 2046 16882
rect 2098 16830 2110 16882
rect 3602 16830 3614 16882
rect 3666 16830 3678 16882
rect 6962 16830 6974 16882
rect 7026 16830 7038 16882
rect 5294 16818 5346 16830
rect 7870 16818 7922 16830
rect 10334 16882 10386 16894
rect 10334 16818 10386 16830
rect 13246 16882 13298 16894
rect 13246 16818 13298 16830
rect 14142 16882 14194 16894
rect 14142 16818 14194 16830
rect 15710 16882 15762 16894
rect 15710 16818 15762 16830
rect 16158 16882 16210 16894
rect 16158 16818 16210 16830
rect 16718 16882 16770 16894
rect 16718 16818 16770 16830
rect 17726 16882 17778 16894
rect 17726 16818 17778 16830
rect 18286 16882 18338 16894
rect 18286 16818 18338 16830
rect 18398 16882 18450 16894
rect 22206 16882 22258 16894
rect 24670 16882 24722 16894
rect 21522 16830 21534 16882
rect 21586 16830 21598 16882
rect 24322 16830 24334 16882
rect 24386 16830 24398 16882
rect 18398 16818 18450 16830
rect 22206 16818 22258 16830
rect 24670 16818 24722 16830
rect 24782 16882 24834 16894
rect 24782 16818 24834 16830
rect 24894 16882 24946 16894
rect 30158 16882 30210 16894
rect 31838 16882 31890 16894
rect 25890 16830 25902 16882
rect 25954 16830 25966 16882
rect 27234 16830 27246 16882
rect 27298 16830 27310 16882
rect 31154 16830 31166 16882
rect 31218 16830 31230 16882
rect 24894 16818 24946 16830
rect 30158 16818 30210 16830
rect 31838 16818 31890 16830
rect 32062 16882 32114 16894
rect 35870 16882 35922 16894
rect 34962 16830 34974 16882
rect 35026 16830 35038 16882
rect 32062 16818 32114 16830
rect 35870 16818 35922 16830
rect 36542 16882 36594 16894
rect 40126 16882 40178 16894
rect 36866 16830 36878 16882
rect 36930 16830 36942 16882
rect 37538 16830 37550 16882
rect 37602 16830 37614 16882
rect 37762 16830 37774 16882
rect 37826 16830 37838 16882
rect 36542 16818 36594 16830
rect 40126 16818 40178 16830
rect 40574 16882 40626 16894
rect 40574 16818 40626 16830
rect 46510 16882 46562 16894
rect 46510 16818 46562 16830
rect 46958 16882 47010 16894
rect 46958 16818 47010 16830
rect 48190 16882 48242 16894
rect 48190 16818 48242 16830
rect 49534 16882 49586 16894
rect 49534 16818 49586 16830
rect 49758 16882 49810 16894
rect 49758 16818 49810 16830
rect 50318 16882 50370 16894
rect 50318 16818 50370 16830
rect 50990 16882 51042 16894
rect 54238 16882 54290 16894
rect 57486 16882 57538 16894
rect 51650 16830 51662 16882
rect 51714 16830 51726 16882
rect 55906 16830 55918 16882
rect 55970 16830 55982 16882
rect 50990 16818 51042 16830
rect 54238 16818 54290 16830
rect 57486 16818 57538 16830
rect 61294 16882 61346 16894
rect 61294 16818 61346 16830
rect 61630 16882 61682 16894
rect 64094 16882 64146 16894
rect 61842 16830 61854 16882
rect 61906 16830 61918 16882
rect 61630 16818 61682 16830
rect 64094 16818 64146 16830
rect 64206 16882 64258 16894
rect 64206 16818 64258 16830
rect 64430 16882 64482 16894
rect 66894 16882 66946 16894
rect 65762 16830 65774 16882
rect 65826 16830 65838 16882
rect 64430 16818 64482 16830
rect 66894 16818 66946 16830
rect 67342 16882 67394 16894
rect 67342 16818 67394 16830
rect 67454 16882 67506 16894
rect 67454 16818 67506 16830
rect 69470 16882 69522 16894
rect 69470 16818 69522 16830
rect 69694 16882 69746 16894
rect 69694 16818 69746 16830
rect 73950 16882 74002 16894
rect 73950 16818 74002 16830
rect 74174 16882 74226 16894
rect 76078 16882 76130 16894
rect 75170 16830 75182 16882
rect 75234 16830 75246 16882
rect 77410 16830 77422 16882
rect 77474 16830 77486 16882
rect 74174 16818 74226 16830
rect 76078 16818 76130 16830
rect 3838 16770 3890 16782
rect 2482 16718 2494 16770
rect 2546 16718 2558 16770
rect 3838 16706 3890 16718
rect 4510 16770 4562 16782
rect 8990 16770 9042 16782
rect 4834 16718 4846 16770
rect 4898 16718 4910 16770
rect 7074 16718 7086 16770
rect 7138 16718 7150 16770
rect 4510 16706 4562 16718
rect 8990 16706 9042 16718
rect 17950 16770 18002 16782
rect 22878 16770 22930 16782
rect 20626 16718 20638 16770
rect 20690 16718 20702 16770
rect 17950 16706 18002 16718
rect 22878 16706 22930 16718
rect 23774 16770 23826 16782
rect 29598 16770 29650 16782
rect 39566 16770 39618 16782
rect 25778 16718 25790 16770
rect 25842 16718 25854 16770
rect 28018 16718 28030 16770
rect 28082 16718 28094 16770
rect 35074 16718 35086 16770
rect 35138 16718 35150 16770
rect 23774 16706 23826 16718
rect 29598 16706 29650 16718
rect 39566 16706 39618 16718
rect 42030 16770 42082 16782
rect 42030 16706 42082 16718
rect 44046 16770 44098 16782
rect 44046 16706 44098 16718
rect 45614 16770 45666 16782
rect 45614 16706 45666 16718
rect 47070 16770 47122 16782
rect 52670 16770 52722 16782
rect 51874 16718 51886 16770
rect 51938 16718 51950 16770
rect 47070 16706 47122 16718
rect 52670 16706 52722 16718
rect 54462 16770 54514 16782
rect 57710 16770 57762 16782
rect 56354 16718 56366 16770
rect 56418 16718 56430 16770
rect 54462 16706 54514 16718
rect 57710 16706 57762 16718
rect 62638 16770 62690 16782
rect 62638 16706 62690 16718
rect 64766 16770 64818 16782
rect 66446 16770 66498 16782
rect 65538 16718 65550 16770
rect 65602 16718 65614 16770
rect 77074 16718 77086 16770
rect 77138 16718 77150 16770
rect 64766 16706 64818 16718
rect 66446 16706 66498 16718
rect 10110 16658 10162 16670
rect 62302 16658 62354 16670
rect 12002 16606 12014 16658
rect 12066 16655 12078 16658
rect 13122 16655 13134 16658
rect 12066 16609 13134 16655
rect 12066 16606 12078 16609
rect 13122 16606 13134 16609
rect 13186 16606 13198 16658
rect 22082 16606 22094 16658
rect 22146 16606 22158 16658
rect 37874 16606 37886 16658
rect 37938 16606 37950 16658
rect 38770 16606 38782 16658
rect 38834 16655 38846 16658
rect 39666 16655 39678 16658
rect 38834 16609 39678 16655
rect 38834 16606 38846 16609
rect 39666 16606 39678 16609
rect 39730 16606 39742 16658
rect 54786 16606 54798 16658
rect 54850 16606 54862 16658
rect 10110 16594 10162 16606
rect 62302 16594 62354 16606
rect 1344 16490 78624 16524
rect 1344 16438 10874 16490
rect 10926 16438 10978 16490
rect 11030 16438 11082 16490
rect 11134 16438 30194 16490
rect 30246 16438 30298 16490
rect 30350 16438 30402 16490
rect 30454 16438 49514 16490
rect 49566 16438 49618 16490
rect 49670 16438 49722 16490
rect 49774 16438 68834 16490
rect 68886 16438 68938 16490
rect 68990 16438 69042 16490
rect 69094 16438 78624 16490
rect 1344 16404 78624 16438
rect 4734 16322 4786 16334
rect 7758 16322 7810 16334
rect 11902 16322 11954 16334
rect 3042 16270 3054 16322
rect 3106 16270 3118 16322
rect 6850 16270 6862 16322
rect 6914 16270 6926 16322
rect 10210 16270 10222 16322
rect 10274 16319 10286 16322
rect 10994 16319 11006 16322
rect 10274 16273 11006 16319
rect 10274 16270 10286 16273
rect 10994 16270 11006 16273
rect 11058 16270 11070 16322
rect 4734 16258 4786 16270
rect 7758 16258 7810 16270
rect 11902 16258 11954 16270
rect 41582 16322 41634 16334
rect 41582 16258 41634 16270
rect 51550 16322 51602 16334
rect 51550 16258 51602 16270
rect 51886 16322 51938 16334
rect 64990 16322 65042 16334
rect 59490 16270 59502 16322
rect 59554 16270 59566 16322
rect 51886 16258 51938 16270
rect 64990 16258 65042 16270
rect 77422 16322 77474 16334
rect 77422 16258 77474 16270
rect 2270 16210 2322 16222
rect 4398 16210 4450 16222
rect 14366 16210 14418 16222
rect 3154 16158 3166 16210
rect 3218 16158 3230 16210
rect 6178 16158 6190 16210
rect 6242 16158 6254 16210
rect 2270 16146 2322 16158
rect 4398 16146 4450 16158
rect 14366 16146 14418 16158
rect 14814 16210 14866 16222
rect 14814 16146 14866 16158
rect 16270 16210 16322 16222
rect 16270 16146 16322 16158
rect 16718 16210 16770 16222
rect 16718 16146 16770 16158
rect 17166 16210 17218 16222
rect 19182 16210 19234 16222
rect 30270 16210 30322 16222
rect 35870 16210 35922 16222
rect 40910 16210 40962 16222
rect 17938 16158 17950 16210
rect 18002 16158 18014 16210
rect 20290 16158 20302 16210
rect 20354 16158 20366 16210
rect 26226 16158 26238 16210
rect 26290 16158 26302 16210
rect 32162 16158 32174 16210
rect 32226 16158 32238 16210
rect 33842 16158 33854 16210
rect 33906 16158 33918 16210
rect 40226 16158 40238 16210
rect 40290 16158 40302 16210
rect 17166 16146 17218 16158
rect 19182 16146 19234 16158
rect 30270 16146 30322 16158
rect 35870 16146 35922 16158
rect 40910 16146 40962 16158
rect 42142 16210 42194 16222
rect 49870 16210 49922 16222
rect 48850 16158 48862 16210
rect 48914 16158 48926 16210
rect 42142 16146 42194 16158
rect 49870 16146 49922 16158
rect 50654 16210 50706 16222
rect 50654 16146 50706 16158
rect 51326 16210 51378 16222
rect 51326 16146 51378 16158
rect 55022 16210 55074 16222
rect 60622 16210 60674 16222
rect 62638 16210 62690 16222
rect 57474 16158 57486 16210
rect 57538 16158 57550 16210
rect 59826 16158 59838 16210
rect 59890 16158 59902 16210
rect 61954 16158 61966 16210
rect 62018 16158 62030 16210
rect 55022 16146 55074 16158
rect 60622 16146 60674 16158
rect 62638 16146 62690 16158
rect 62862 16210 62914 16222
rect 62862 16146 62914 16158
rect 63646 16210 63698 16222
rect 70366 16210 70418 16222
rect 75518 16210 75570 16222
rect 66434 16158 66446 16210
rect 66498 16158 66510 16210
rect 72482 16158 72494 16210
rect 72546 16158 72558 16210
rect 74386 16158 74398 16210
rect 74450 16158 74462 16210
rect 63646 16146 63698 16158
rect 70366 16146 70418 16158
rect 75518 16146 75570 16158
rect 77982 16210 78034 16222
rect 77982 16146 78034 16158
rect 7646 16098 7698 16110
rect 3602 16046 3614 16098
rect 3666 16046 3678 16098
rect 6626 16046 6638 16098
rect 6690 16046 6702 16098
rect 7646 16034 7698 16046
rect 9662 16098 9714 16110
rect 9662 16034 9714 16046
rect 11342 16098 11394 16110
rect 11342 16034 11394 16046
rect 11454 16098 11506 16110
rect 13918 16098 13970 16110
rect 11554 16046 11566 16098
rect 11618 16046 11630 16098
rect 11454 16034 11506 16046
rect 13918 16034 13970 16046
rect 18174 16098 18226 16110
rect 18174 16034 18226 16046
rect 20414 16098 20466 16110
rect 20414 16034 20466 16046
rect 21646 16098 21698 16110
rect 21646 16034 21698 16046
rect 22206 16098 22258 16110
rect 22206 16034 22258 16046
rect 22654 16098 22706 16110
rect 24782 16098 24834 16110
rect 24210 16046 24222 16098
rect 24274 16046 24286 16098
rect 22654 16034 22706 16046
rect 24782 16034 24834 16046
rect 24894 16098 24946 16110
rect 26910 16098 26962 16110
rect 26114 16046 26126 16098
rect 26178 16046 26190 16098
rect 24894 16034 24946 16046
rect 26910 16034 26962 16046
rect 27246 16098 27298 16110
rect 27246 16034 27298 16046
rect 30830 16098 30882 16110
rect 35086 16098 35138 16110
rect 31938 16046 31950 16098
rect 32002 16046 32014 16098
rect 30830 16034 30882 16046
rect 35086 16034 35138 16046
rect 35422 16098 35474 16110
rect 39006 16098 39058 16110
rect 38434 16046 38446 16098
rect 38498 16046 38510 16098
rect 35422 16034 35474 16046
rect 39006 16034 39058 16046
rect 39902 16098 39954 16110
rect 39902 16034 39954 16046
rect 40126 16098 40178 16110
rect 40126 16034 40178 16046
rect 46286 16098 46338 16110
rect 46286 16034 46338 16046
rect 46398 16098 46450 16110
rect 46398 16034 46450 16046
rect 47630 16098 47682 16110
rect 49422 16098 49474 16110
rect 48514 16046 48526 16098
rect 48578 16046 48590 16098
rect 47630 16034 47682 16046
rect 49422 16034 49474 16046
rect 54574 16098 54626 16110
rect 54574 16034 54626 16046
rect 55582 16098 55634 16110
rect 55582 16034 55634 16046
rect 55918 16098 55970 16110
rect 55918 16034 55970 16046
rect 56590 16098 56642 16110
rect 56590 16034 56642 16046
rect 56926 16098 56978 16110
rect 61854 16098 61906 16110
rect 64318 16098 64370 16110
rect 59938 16046 59950 16098
rect 60002 16046 60014 16098
rect 61394 16046 61406 16098
rect 61458 16046 61470 16098
rect 62066 16046 62078 16098
rect 62130 16046 62142 16098
rect 56926 16034 56978 16046
rect 61854 16034 61906 16046
rect 64318 16034 64370 16046
rect 65326 16098 65378 16110
rect 73278 16098 73330 16110
rect 74846 16098 74898 16110
rect 66210 16046 66222 16098
rect 66274 16046 66286 16098
rect 69906 16046 69918 16098
rect 69970 16046 69982 16098
rect 70130 16046 70142 16098
rect 70194 16046 70206 16098
rect 72370 16046 72382 16098
rect 72434 16046 72446 16098
rect 74162 16046 74174 16098
rect 74226 16046 74238 16098
rect 65326 16034 65378 16046
rect 73278 16034 73330 16046
rect 74846 16034 74898 16046
rect 75966 16098 76018 16110
rect 75966 16034 76018 16046
rect 76302 16098 76354 16110
rect 76302 16034 76354 16046
rect 4622 15986 4674 15998
rect 4622 15922 4674 15934
rect 7758 15986 7810 15998
rect 7758 15922 7810 15934
rect 9998 15986 10050 15998
rect 9998 15922 10050 15934
rect 12574 15986 12626 15998
rect 12574 15922 12626 15934
rect 12686 15986 12738 15998
rect 12686 15922 12738 15934
rect 13806 15986 13858 15998
rect 13806 15922 13858 15934
rect 17950 15986 18002 15998
rect 17950 15922 18002 15934
rect 18398 15986 18450 15998
rect 18398 15922 18450 15934
rect 19630 15986 19682 15998
rect 19630 15922 19682 15934
rect 20302 15986 20354 15998
rect 20302 15922 20354 15934
rect 20862 15986 20914 15998
rect 20862 15922 20914 15934
rect 26462 15986 26514 15998
rect 26462 15922 26514 15934
rect 27134 15986 27186 15998
rect 27134 15922 27186 15934
rect 29598 15986 29650 15998
rect 29598 15922 29650 15934
rect 32622 15986 32674 15998
rect 32622 15922 32674 15934
rect 33518 15986 33570 15998
rect 33518 15922 33570 15934
rect 34414 15986 34466 15998
rect 34414 15922 34466 15934
rect 39118 15986 39170 15998
rect 39118 15922 39170 15934
rect 39678 15986 39730 15998
rect 39678 15922 39730 15934
rect 41582 15986 41634 15998
rect 41582 15922 41634 15934
rect 41694 15986 41746 15998
rect 41694 15922 41746 15934
rect 46622 15986 46674 15998
rect 46622 15922 46674 15934
rect 47742 15986 47794 15998
rect 47742 15922 47794 15934
rect 56366 15986 56418 15998
rect 56366 15922 56418 15934
rect 57822 15986 57874 15998
rect 57822 15922 57874 15934
rect 64878 15986 64930 15998
rect 64878 15922 64930 15934
rect 66894 15986 66946 15998
rect 66894 15922 66946 15934
rect 76078 15986 76130 15998
rect 76078 15922 76130 15934
rect 77310 15986 77362 15998
rect 77310 15922 77362 15934
rect 9214 15874 9266 15886
rect 9214 15810 9266 15822
rect 9886 15874 9938 15886
rect 9886 15810 9938 15822
rect 10446 15874 10498 15886
rect 10446 15810 10498 15822
rect 11230 15874 11282 15886
rect 11230 15810 11282 15822
rect 12350 15874 12402 15886
rect 12350 15810 12402 15822
rect 13582 15874 13634 15886
rect 13582 15810 13634 15822
rect 15262 15874 15314 15886
rect 15262 15810 15314 15822
rect 15934 15874 15986 15886
rect 15934 15810 15986 15822
rect 17838 15874 17890 15886
rect 17838 15810 17890 15822
rect 20638 15874 20690 15886
rect 20638 15810 20690 15822
rect 23326 15874 23378 15886
rect 23326 15810 23378 15822
rect 25454 15874 25506 15886
rect 25454 15810 25506 15822
rect 28814 15874 28866 15886
rect 28814 15810 28866 15822
rect 29710 15874 29762 15886
rect 29710 15810 29762 15822
rect 29934 15874 29986 15886
rect 29934 15810 29986 15822
rect 30942 15874 30994 15886
rect 30942 15810 30994 15822
rect 31166 15874 31218 15886
rect 31166 15810 31218 15822
rect 33742 15874 33794 15886
rect 33742 15810 33794 15822
rect 34526 15874 34578 15886
rect 34526 15810 34578 15822
rect 34750 15874 34802 15886
rect 34750 15810 34802 15822
rect 35310 15874 35362 15886
rect 35310 15810 35362 15822
rect 37662 15874 37714 15886
rect 37662 15810 37714 15822
rect 40238 15874 40290 15886
rect 40238 15810 40290 15822
rect 42702 15874 42754 15886
rect 42702 15810 42754 15822
rect 46174 15874 46226 15886
rect 46174 15810 46226 15822
rect 47966 15874 48018 15886
rect 47966 15810 48018 15822
rect 55694 15874 55746 15886
rect 55694 15810 55746 15822
rect 56590 15874 56642 15886
rect 56590 15810 56642 15822
rect 57598 15874 57650 15886
rect 57598 15810 57650 15822
rect 61630 15874 61682 15886
rect 64654 15874 64706 15886
rect 63186 15822 63198 15874
rect 63250 15822 63262 15874
rect 61630 15810 61682 15822
rect 64654 15810 64706 15822
rect 70814 15874 70866 15886
rect 70814 15810 70866 15822
rect 71262 15874 71314 15886
rect 71262 15810 71314 15822
rect 77422 15874 77474 15886
rect 77422 15810 77474 15822
rect 1344 15706 78784 15740
rect 1344 15654 20534 15706
rect 20586 15654 20638 15706
rect 20690 15654 20742 15706
rect 20794 15654 39854 15706
rect 39906 15654 39958 15706
rect 40010 15654 40062 15706
rect 40114 15654 59174 15706
rect 59226 15654 59278 15706
rect 59330 15654 59382 15706
rect 59434 15654 78494 15706
rect 78546 15654 78598 15706
rect 78650 15654 78702 15706
rect 78754 15654 78784 15706
rect 1344 15620 78784 15654
rect 2382 15538 2434 15550
rect 2382 15474 2434 15486
rect 5854 15538 5906 15550
rect 15262 15538 15314 15550
rect 11554 15486 11566 15538
rect 11618 15486 11630 15538
rect 14466 15486 14478 15538
rect 14530 15486 14542 15538
rect 5854 15474 5906 15486
rect 15262 15474 15314 15486
rect 15710 15538 15762 15550
rect 15710 15474 15762 15486
rect 17054 15538 17106 15550
rect 17054 15474 17106 15486
rect 18510 15538 18562 15550
rect 18510 15474 18562 15486
rect 19182 15538 19234 15550
rect 19182 15474 19234 15486
rect 19406 15538 19458 15550
rect 19406 15474 19458 15486
rect 19966 15538 20018 15550
rect 19966 15474 20018 15486
rect 20638 15538 20690 15550
rect 20638 15474 20690 15486
rect 21534 15538 21586 15550
rect 21534 15474 21586 15486
rect 21646 15538 21698 15550
rect 21646 15474 21698 15486
rect 28142 15538 28194 15550
rect 28142 15474 28194 15486
rect 30494 15538 30546 15550
rect 30494 15474 30546 15486
rect 31726 15538 31778 15550
rect 31726 15474 31778 15486
rect 31950 15538 32002 15550
rect 31950 15474 32002 15486
rect 34190 15538 34242 15550
rect 34190 15474 34242 15486
rect 34302 15538 34354 15550
rect 34302 15474 34354 15486
rect 35198 15538 35250 15550
rect 35198 15474 35250 15486
rect 35646 15538 35698 15550
rect 35646 15474 35698 15486
rect 39678 15538 39730 15550
rect 39678 15474 39730 15486
rect 45502 15538 45554 15550
rect 45502 15474 45554 15486
rect 46174 15538 46226 15550
rect 46174 15474 46226 15486
rect 47294 15538 47346 15550
rect 47294 15474 47346 15486
rect 50878 15538 50930 15550
rect 50878 15474 50930 15486
rect 57374 15538 57426 15550
rect 57374 15474 57426 15486
rect 60286 15538 60338 15550
rect 60286 15474 60338 15486
rect 61294 15538 61346 15550
rect 61294 15474 61346 15486
rect 61966 15538 62018 15550
rect 61966 15474 62018 15486
rect 62302 15538 62354 15550
rect 62302 15474 62354 15486
rect 64318 15538 64370 15550
rect 64318 15474 64370 15486
rect 65886 15538 65938 15550
rect 65886 15474 65938 15486
rect 69470 15538 69522 15550
rect 69470 15474 69522 15486
rect 70254 15538 70306 15550
rect 70254 15474 70306 15486
rect 71038 15538 71090 15550
rect 71038 15474 71090 15486
rect 73726 15538 73778 15550
rect 73726 15474 73778 15486
rect 75406 15538 75458 15550
rect 75406 15474 75458 15486
rect 78094 15538 78146 15550
rect 78094 15474 78146 15486
rect 2830 15426 2882 15438
rect 16718 15426 16770 15438
rect 12674 15374 12686 15426
rect 12738 15374 12750 15426
rect 2830 15362 2882 15374
rect 16718 15362 16770 15374
rect 16830 15426 16882 15438
rect 16830 15362 16882 15374
rect 21086 15426 21138 15438
rect 21086 15362 21138 15374
rect 24558 15426 24610 15438
rect 24558 15362 24610 15374
rect 43374 15426 43426 15438
rect 43374 15362 43426 15374
rect 44046 15426 44098 15438
rect 44046 15362 44098 15374
rect 44158 15426 44210 15438
rect 50542 15426 50594 15438
rect 46386 15374 46398 15426
rect 46450 15423 46462 15426
rect 46722 15423 46734 15426
rect 46450 15377 46734 15423
rect 46450 15374 46462 15377
rect 46722 15374 46734 15377
rect 46786 15374 46798 15426
rect 44158 15362 44210 15374
rect 50542 15362 50594 15374
rect 50654 15426 50706 15438
rect 50654 15362 50706 15374
rect 51214 15426 51266 15438
rect 51214 15362 51266 15374
rect 70926 15426 70978 15438
rect 70926 15362 70978 15374
rect 71598 15426 71650 15438
rect 71598 15362 71650 15374
rect 73390 15426 73442 15438
rect 73390 15362 73442 15374
rect 73502 15426 73554 15438
rect 73502 15362 73554 15374
rect 74062 15426 74114 15438
rect 74062 15362 74114 15374
rect 74510 15426 74562 15438
rect 74510 15362 74562 15374
rect 76862 15426 76914 15438
rect 76862 15362 76914 15374
rect 77534 15426 77586 15438
rect 77534 15362 77586 15374
rect 3950 15314 4002 15326
rect 3042 15262 3054 15314
rect 3106 15262 3118 15314
rect 3950 15250 4002 15262
rect 5406 15314 5458 15326
rect 11006 15314 11058 15326
rect 18286 15314 18338 15326
rect 19518 15314 19570 15326
rect 8530 15262 8542 15314
rect 8594 15262 8606 15314
rect 13234 15262 13246 15314
rect 13298 15262 13310 15314
rect 13906 15262 13918 15314
rect 13970 15262 13982 15314
rect 18050 15262 18062 15314
rect 18114 15262 18126 15314
rect 18722 15262 18734 15314
rect 18786 15262 18798 15314
rect 5406 15250 5458 15262
rect 11006 15250 11058 15262
rect 18286 15250 18338 15262
rect 19518 15250 19570 15262
rect 21310 15314 21362 15326
rect 21310 15250 21362 15262
rect 22878 15314 22930 15326
rect 28030 15314 28082 15326
rect 23986 15262 23998 15314
rect 24050 15262 24062 15314
rect 22878 15250 22930 15262
rect 28030 15250 28082 15262
rect 28254 15314 28306 15326
rect 28254 15250 28306 15262
rect 28702 15314 28754 15326
rect 28702 15250 28754 15262
rect 31838 15314 31890 15326
rect 31838 15250 31890 15262
rect 32398 15314 32450 15326
rect 32398 15250 32450 15262
rect 34414 15314 34466 15326
rect 39118 15314 39170 15326
rect 34738 15262 34750 15314
rect 34802 15262 34814 15314
rect 38770 15262 38782 15314
rect 38834 15262 38846 15314
rect 34414 15250 34466 15262
rect 39118 15250 39170 15262
rect 42478 15314 42530 15326
rect 43822 15314 43874 15326
rect 43026 15262 43038 15314
rect 43090 15262 43102 15314
rect 42478 15250 42530 15262
rect 43822 15250 43874 15262
rect 44606 15314 44658 15326
rect 46286 15314 46338 15326
rect 45938 15262 45950 15314
rect 46002 15262 46014 15314
rect 44606 15250 44658 15262
rect 46286 15250 46338 15262
rect 46846 15314 46898 15326
rect 46846 15250 46898 15262
rect 47966 15314 48018 15326
rect 51662 15314 51714 15326
rect 53118 15314 53170 15326
rect 60062 15314 60114 15326
rect 48402 15262 48414 15314
rect 48466 15262 48478 15314
rect 52770 15262 52782 15314
rect 52834 15262 52846 15314
rect 54114 15262 54126 15314
rect 54178 15262 54190 15314
rect 47966 15250 48018 15262
rect 51662 15250 51714 15262
rect 53118 15250 53170 15262
rect 60062 15250 60114 15262
rect 60398 15314 60450 15326
rect 60398 15250 60450 15262
rect 60734 15314 60786 15326
rect 60734 15250 60786 15262
rect 62974 15314 63026 15326
rect 68910 15314 68962 15326
rect 71262 15314 71314 15326
rect 76750 15314 76802 15326
rect 63298 15262 63310 15314
rect 63362 15262 63374 15314
rect 70018 15262 70030 15314
rect 70082 15262 70094 15314
rect 76178 15262 76190 15314
rect 76242 15262 76254 15314
rect 62974 15250 63026 15262
rect 68910 15250 68962 15262
rect 71262 15250 71314 15262
rect 76750 15250 76802 15262
rect 77422 15314 77474 15326
rect 77422 15250 77474 15262
rect 4510 15202 4562 15214
rect 4510 15138 4562 15150
rect 4958 15202 5010 15214
rect 4958 15138 5010 15150
rect 8990 15202 9042 15214
rect 8990 15138 9042 15150
rect 9662 15202 9714 15214
rect 9662 15138 9714 15150
rect 11230 15202 11282 15214
rect 11230 15138 11282 15150
rect 16270 15202 16322 15214
rect 16270 15138 16322 15150
rect 18398 15202 18450 15214
rect 18398 15138 18450 15150
rect 21422 15202 21474 15214
rect 21422 15138 21474 15150
rect 22430 15202 22482 15214
rect 27470 15202 27522 15214
rect 23874 15150 23886 15202
rect 23938 15150 23950 15202
rect 22430 15138 22482 15150
rect 27470 15138 27522 15150
rect 30046 15202 30098 15214
rect 30046 15138 30098 15150
rect 32174 15202 32226 15214
rect 32174 15138 32226 15150
rect 38222 15202 38274 15214
rect 62862 15202 62914 15214
rect 43138 15150 43150 15202
rect 43202 15150 43214 15202
rect 38222 15138 38274 15150
rect 62862 15138 62914 15150
rect 65326 15202 65378 15214
rect 65326 15138 65378 15150
rect 70366 15202 70418 15214
rect 70366 15138 70418 15150
rect 72494 15202 72546 15214
rect 72494 15138 72546 15150
rect 72606 15090 72658 15102
rect 54002 15038 54014 15090
rect 54066 15038 54078 15090
rect 72606 15026 72658 15038
rect 77534 15090 77586 15102
rect 77534 15026 77586 15038
rect 1344 14922 78624 14956
rect 1344 14870 10874 14922
rect 10926 14870 10978 14922
rect 11030 14870 11082 14922
rect 11134 14870 30194 14922
rect 30246 14870 30298 14922
rect 30350 14870 30402 14922
rect 30454 14870 49514 14922
rect 49566 14870 49618 14922
rect 49670 14870 49722 14922
rect 49774 14870 68834 14922
rect 68886 14870 68938 14922
rect 68990 14870 69042 14922
rect 69094 14870 78624 14922
rect 1344 14836 78624 14870
rect 3726 14754 3778 14766
rect 3726 14690 3778 14702
rect 13806 14754 13858 14766
rect 13806 14690 13858 14702
rect 28030 14754 28082 14766
rect 28030 14690 28082 14702
rect 28702 14754 28754 14766
rect 28702 14690 28754 14702
rect 39790 14754 39842 14766
rect 58046 14754 58098 14766
rect 46722 14702 46734 14754
rect 46786 14702 46798 14754
rect 56690 14702 56702 14754
rect 56754 14702 56766 14754
rect 39790 14690 39842 14702
rect 58046 14690 58098 14702
rect 63870 14754 63922 14766
rect 63870 14690 63922 14702
rect 64206 14754 64258 14766
rect 64206 14690 64258 14702
rect 77422 14754 77474 14766
rect 77422 14690 77474 14702
rect 5630 14642 5682 14654
rect 5630 14578 5682 14590
rect 9438 14642 9490 14654
rect 9438 14578 9490 14590
rect 17054 14642 17106 14654
rect 20302 14642 20354 14654
rect 17602 14590 17614 14642
rect 17666 14590 17678 14642
rect 19842 14590 19854 14642
rect 19906 14590 19918 14642
rect 17054 14578 17106 14590
rect 20302 14578 20354 14590
rect 20862 14642 20914 14654
rect 20862 14578 20914 14590
rect 21646 14642 21698 14654
rect 21646 14578 21698 14590
rect 22542 14642 22594 14654
rect 22542 14578 22594 14590
rect 24670 14642 24722 14654
rect 24670 14578 24722 14590
rect 26126 14642 26178 14654
rect 36206 14642 36258 14654
rect 49422 14642 49474 14654
rect 32498 14590 32510 14642
rect 32562 14590 32574 14642
rect 38210 14590 38222 14642
rect 38274 14590 38286 14642
rect 42242 14590 42254 14642
rect 42306 14590 42318 14642
rect 46162 14590 46174 14642
rect 46226 14590 46238 14642
rect 26126 14578 26178 14590
rect 36206 14578 36258 14590
rect 49422 14578 49474 14590
rect 51998 14642 52050 14654
rect 59614 14642 59666 14654
rect 57026 14590 57038 14642
rect 57090 14590 57102 14642
rect 51998 14578 52050 14590
rect 59614 14578 59666 14590
rect 61518 14642 61570 14654
rect 61518 14578 61570 14590
rect 63646 14642 63698 14654
rect 67902 14642 67954 14654
rect 72382 14642 72434 14654
rect 73950 14642 74002 14654
rect 66994 14590 67006 14642
rect 67058 14590 67070 14642
rect 69682 14590 69694 14642
rect 69746 14590 69758 14642
rect 73042 14590 73054 14642
rect 73106 14590 73118 14642
rect 63646 14578 63698 14590
rect 67902 14578 67954 14590
rect 72382 14578 72434 14590
rect 73950 14578 74002 14590
rect 74510 14642 74562 14654
rect 74510 14578 74562 14590
rect 4622 14530 4674 14542
rect 8654 14530 8706 14542
rect 2818 14478 2830 14530
rect 2882 14478 2894 14530
rect 8082 14478 8094 14530
rect 8146 14478 8158 14530
rect 4622 14466 4674 14478
rect 8654 14466 8706 14478
rect 8766 14530 8818 14542
rect 8766 14466 8818 14478
rect 9998 14530 10050 14542
rect 9998 14466 10050 14478
rect 12462 14530 12514 14542
rect 12910 14530 12962 14542
rect 12562 14478 12574 14530
rect 12626 14478 12638 14530
rect 12462 14466 12514 14478
rect 12910 14466 12962 14478
rect 13694 14530 13746 14542
rect 24222 14530 24274 14542
rect 26014 14530 26066 14542
rect 34750 14530 34802 14542
rect 18050 14478 18062 14530
rect 18114 14478 18126 14530
rect 19170 14478 19182 14530
rect 19234 14478 19246 14530
rect 25442 14478 25454 14530
rect 25506 14478 25518 14530
rect 28018 14478 28030 14530
rect 28082 14478 28094 14530
rect 32386 14478 32398 14530
rect 32450 14478 32462 14530
rect 33506 14478 33518 14530
rect 33570 14478 33582 14530
rect 13694 14466 13746 14478
rect 24222 14466 24274 14478
rect 26014 14466 26066 14478
rect 34750 14466 34802 14478
rect 34974 14530 35026 14542
rect 40686 14530 40738 14542
rect 49310 14530 49362 14542
rect 38434 14478 38446 14530
rect 38498 14478 38510 14530
rect 45938 14478 45950 14530
rect 46002 14478 46014 14530
rect 48738 14478 48750 14530
rect 48802 14478 48814 14530
rect 34974 14466 35026 14478
rect 40686 14466 40738 14478
rect 49310 14466 49362 14478
rect 51102 14530 51154 14542
rect 54910 14530 54962 14542
rect 60510 14530 60562 14542
rect 54002 14478 54014 14530
rect 54066 14478 54078 14530
rect 54226 14478 54238 14530
rect 54290 14478 54302 14530
rect 57138 14478 57150 14530
rect 57202 14478 57214 14530
rect 60050 14478 60062 14530
rect 60114 14478 60126 14530
rect 51102 14466 51154 14478
rect 54910 14466 54962 14478
rect 60510 14466 60562 14478
rect 62078 14530 62130 14542
rect 62078 14466 62130 14478
rect 62414 14530 62466 14542
rect 67678 14530 67730 14542
rect 66882 14478 66894 14530
rect 66946 14478 66958 14530
rect 62414 14466 62466 14478
rect 67678 14466 67730 14478
rect 68014 14530 68066 14542
rect 70478 14530 70530 14542
rect 70018 14478 70030 14530
rect 70082 14478 70094 14530
rect 68014 14466 68066 14478
rect 70478 14466 70530 14478
rect 71486 14530 71538 14542
rect 77534 14530 77586 14542
rect 71698 14478 71710 14530
rect 71762 14478 71774 14530
rect 73490 14478 73502 14530
rect 73554 14478 73566 14530
rect 75058 14478 75070 14530
rect 75122 14478 75134 14530
rect 71486 14466 71538 14478
rect 77534 14466 77586 14478
rect 3838 14418 3890 14430
rect 1922 14366 1934 14418
rect 1986 14366 1998 14418
rect 3838 14354 3890 14366
rect 4510 14418 4562 14430
rect 4510 14354 4562 14366
rect 7086 14418 7138 14430
rect 7086 14354 7138 14366
rect 9326 14418 9378 14430
rect 9326 14354 9378 14366
rect 12238 14418 12290 14430
rect 12238 14354 12290 14366
rect 13806 14418 13858 14430
rect 13806 14354 13858 14366
rect 14366 14418 14418 14430
rect 14366 14354 14418 14366
rect 14590 14418 14642 14430
rect 14590 14354 14642 14366
rect 14702 14418 14754 14430
rect 14702 14354 14754 14366
rect 15598 14418 15650 14430
rect 15598 14354 15650 14366
rect 23886 14418 23938 14430
rect 23886 14354 23938 14366
rect 27694 14418 27746 14430
rect 27694 14354 27746 14366
rect 28814 14418 28866 14430
rect 39118 14418 39170 14430
rect 33954 14366 33966 14418
rect 34018 14366 34030 14418
rect 28814 14354 28866 14366
rect 39118 14354 39170 14366
rect 39902 14418 39954 14430
rect 39902 14354 39954 14366
rect 40350 14418 40402 14430
rect 40350 14354 40402 14366
rect 40574 14418 40626 14430
rect 44382 14418 44434 14430
rect 42466 14366 42478 14418
rect 42530 14366 42542 14418
rect 44146 14366 44158 14418
rect 44210 14366 44222 14418
rect 40574 14354 40626 14366
rect 44382 14354 44434 14366
rect 49982 14418 50034 14430
rect 49982 14354 50034 14366
rect 50318 14418 50370 14430
rect 50318 14354 50370 14366
rect 50766 14418 50818 14430
rect 50766 14354 50818 14366
rect 54462 14418 54514 14430
rect 54462 14354 54514 14366
rect 58158 14418 58210 14430
rect 58158 14354 58210 14366
rect 62750 14418 62802 14430
rect 62750 14354 62802 14366
rect 66110 14418 66162 14430
rect 66110 14354 66162 14366
rect 68350 14418 68402 14430
rect 76066 14366 76078 14418
rect 76130 14366 76142 14418
rect 68350 14354 68402 14366
rect 3726 14306 3778 14318
rect 3726 14242 3778 14254
rect 4286 14306 4338 14318
rect 4286 14242 4338 14254
rect 6078 14306 6130 14318
rect 6078 14242 6130 14254
rect 6638 14306 6690 14318
rect 6638 14242 6690 14254
rect 7198 14306 7250 14318
rect 7198 14242 7250 14254
rect 9550 14306 9602 14318
rect 9550 14242 9602 14254
rect 12350 14306 12402 14318
rect 12350 14242 12402 14254
rect 15150 14306 15202 14318
rect 15150 14242 15202 14254
rect 16158 14306 16210 14318
rect 16158 14242 16210 14254
rect 16494 14306 16546 14318
rect 16494 14242 16546 14254
rect 21982 14306 22034 14318
rect 21982 14242 22034 14254
rect 23998 14306 24050 14318
rect 23998 14242 24050 14254
rect 28702 14306 28754 14318
rect 35758 14306 35810 14318
rect 35298 14254 35310 14306
rect 35362 14254 35374 14306
rect 28702 14242 28754 14254
rect 35758 14242 35810 14254
rect 37662 14306 37714 14318
rect 37662 14242 37714 14254
rect 39790 14306 39842 14318
rect 39790 14242 39842 14254
rect 41582 14306 41634 14318
rect 41582 14242 41634 14254
rect 50094 14306 50146 14318
rect 50094 14242 50146 14254
rect 50878 14306 50930 14318
rect 50878 14242 50930 14254
rect 58046 14306 58098 14318
rect 58046 14242 58098 14254
rect 61406 14306 61458 14318
rect 61406 14242 61458 14254
rect 61630 14306 61682 14318
rect 61630 14242 61682 14254
rect 62638 14306 62690 14318
rect 62638 14242 62690 14254
rect 77422 14306 77474 14318
rect 77422 14242 77474 14254
rect 1344 14138 78784 14172
rect 1344 14086 20534 14138
rect 20586 14086 20638 14138
rect 20690 14086 20742 14138
rect 20794 14086 39854 14138
rect 39906 14086 39958 14138
rect 40010 14086 40062 14138
rect 40114 14086 59174 14138
rect 59226 14086 59278 14138
rect 59330 14086 59382 14138
rect 59434 14086 78494 14138
rect 78546 14086 78598 14138
rect 78650 14086 78702 14138
rect 78754 14086 78784 14138
rect 1344 14052 78784 14086
rect 4510 13970 4562 13982
rect 4510 13906 4562 13918
rect 9886 13970 9938 13982
rect 16830 13970 16882 13982
rect 12002 13918 12014 13970
rect 12066 13918 12078 13970
rect 9886 13906 9938 13918
rect 16830 13906 16882 13918
rect 17054 13970 17106 13982
rect 17054 13906 17106 13918
rect 18846 13970 18898 13982
rect 18846 13906 18898 13918
rect 18958 13970 19010 13982
rect 18958 13906 19010 13918
rect 19854 13970 19906 13982
rect 19854 13906 19906 13918
rect 26238 13970 26290 13982
rect 26238 13906 26290 13918
rect 35086 13970 35138 13982
rect 35086 13906 35138 13918
rect 37662 13970 37714 13982
rect 37662 13906 37714 13918
rect 40686 13970 40738 13982
rect 40686 13906 40738 13918
rect 43150 13970 43202 13982
rect 43150 13906 43202 13918
rect 43262 13970 43314 13982
rect 43262 13906 43314 13918
rect 43374 13970 43426 13982
rect 43374 13906 43426 13918
rect 46286 13970 46338 13982
rect 46286 13906 46338 13918
rect 46510 13970 46562 13982
rect 46510 13906 46562 13918
rect 48414 13970 48466 13982
rect 48414 13906 48466 13918
rect 55134 13970 55186 13982
rect 55134 13906 55186 13918
rect 64654 13970 64706 13982
rect 64654 13906 64706 13918
rect 67230 13970 67282 13982
rect 67230 13906 67282 13918
rect 67454 13970 67506 13982
rect 67454 13906 67506 13918
rect 67790 13970 67842 13982
rect 67790 13906 67842 13918
rect 72046 13970 72098 13982
rect 72046 13906 72098 13918
rect 72158 13970 72210 13982
rect 72158 13906 72210 13918
rect 2382 13858 2434 13870
rect 2382 13794 2434 13806
rect 4062 13858 4114 13870
rect 4062 13794 4114 13806
rect 4734 13858 4786 13870
rect 4734 13794 4786 13806
rect 8654 13858 8706 13870
rect 14814 13858 14866 13870
rect 12898 13806 12910 13858
rect 12962 13806 12974 13858
rect 8654 13794 8706 13806
rect 14814 13794 14866 13806
rect 23102 13858 23154 13870
rect 23102 13794 23154 13806
rect 24782 13858 24834 13870
rect 24782 13794 24834 13806
rect 26014 13858 26066 13870
rect 26014 13794 26066 13806
rect 26686 13858 26738 13870
rect 37886 13858 37938 13870
rect 30146 13806 30158 13858
rect 30210 13806 30222 13858
rect 26686 13794 26738 13806
rect 37886 13794 37938 13806
rect 37998 13858 38050 13870
rect 37998 13794 38050 13806
rect 45390 13858 45442 13870
rect 45390 13794 45442 13806
rect 46174 13858 46226 13870
rect 46174 13794 46226 13806
rect 48638 13858 48690 13870
rect 48638 13794 48690 13806
rect 49534 13858 49586 13870
rect 49534 13794 49586 13806
rect 53790 13858 53842 13870
rect 53790 13794 53842 13806
rect 61070 13858 61122 13870
rect 61070 13794 61122 13806
rect 62526 13858 62578 13870
rect 62526 13794 62578 13806
rect 65438 13858 65490 13870
rect 65438 13794 65490 13806
rect 65550 13858 65602 13870
rect 65550 13794 65602 13806
rect 67118 13858 67170 13870
rect 67118 13794 67170 13806
rect 68238 13858 68290 13870
rect 68238 13794 68290 13806
rect 73502 13858 73554 13870
rect 73502 13794 73554 13806
rect 73614 13858 73666 13870
rect 73614 13794 73666 13806
rect 75406 13858 75458 13870
rect 75406 13794 75458 13806
rect 2270 13746 2322 13758
rect 2270 13682 2322 13694
rect 2606 13746 2658 13758
rect 4846 13746 4898 13758
rect 3378 13694 3390 13746
rect 3442 13694 3454 13746
rect 2606 13682 2658 13694
rect 4846 13682 4898 13694
rect 5742 13746 5794 13758
rect 9774 13746 9826 13758
rect 8194 13694 8206 13746
rect 8258 13694 8270 13746
rect 5742 13682 5794 13694
rect 9774 13682 9826 13694
rect 11454 13746 11506 13758
rect 16718 13746 16770 13758
rect 14130 13694 14142 13746
rect 14194 13694 14206 13746
rect 11454 13682 11506 13694
rect 16718 13682 16770 13694
rect 17838 13746 17890 13758
rect 17838 13682 17890 13694
rect 18398 13746 18450 13758
rect 18398 13682 18450 13694
rect 18622 13746 18674 13758
rect 18622 13682 18674 13694
rect 19070 13746 19122 13758
rect 24670 13746 24722 13758
rect 20962 13694 20974 13746
rect 21026 13694 21038 13746
rect 22530 13694 22542 13746
rect 22594 13694 22606 13746
rect 19070 13682 19122 13694
rect 24670 13682 24722 13694
rect 25006 13746 25058 13758
rect 25006 13682 25058 13694
rect 25566 13746 25618 13758
rect 25566 13682 25618 13694
rect 27470 13746 27522 13758
rect 34750 13746 34802 13758
rect 28130 13694 28142 13746
rect 28194 13694 28206 13746
rect 29474 13694 29486 13746
rect 29538 13694 29550 13746
rect 27470 13682 27522 13694
rect 34750 13682 34802 13694
rect 34862 13746 34914 13758
rect 34862 13682 34914 13694
rect 35310 13746 35362 13758
rect 35310 13682 35362 13694
rect 35982 13746 36034 13758
rect 39678 13746 39730 13758
rect 40574 13746 40626 13758
rect 38882 13694 38894 13746
rect 38946 13694 38958 13746
rect 40226 13694 40238 13746
rect 40290 13694 40302 13746
rect 35982 13682 36034 13694
rect 39678 13682 39730 13694
rect 40574 13682 40626 13694
rect 40798 13746 40850 13758
rect 40798 13682 40850 13694
rect 43822 13746 43874 13758
rect 48750 13746 48802 13758
rect 54014 13746 54066 13758
rect 44930 13694 44942 13746
rect 44994 13694 45006 13746
rect 49970 13694 49982 13746
rect 50034 13694 50046 13746
rect 43822 13682 43874 13694
rect 48750 13682 48802 13694
rect 54014 13682 54066 13694
rect 54910 13746 54962 13758
rect 54910 13682 54962 13694
rect 55134 13746 55186 13758
rect 55134 13682 55186 13694
rect 55470 13746 55522 13758
rect 60286 13746 60338 13758
rect 59826 13694 59838 13746
rect 59890 13694 59902 13746
rect 55470 13682 55522 13694
rect 60286 13682 60338 13694
rect 62750 13746 62802 13758
rect 65774 13746 65826 13758
rect 62962 13694 62974 13746
rect 63026 13694 63038 13746
rect 62750 13682 62802 13694
rect 65774 13682 65826 13694
rect 66558 13746 66610 13758
rect 66558 13682 66610 13694
rect 71486 13746 71538 13758
rect 71486 13682 71538 13694
rect 72270 13746 72322 13758
rect 72270 13682 72322 13694
rect 72718 13746 72770 13758
rect 72718 13682 72770 13694
rect 73278 13746 73330 13758
rect 73278 13682 73330 13694
rect 75294 13746 75346 13758
rect 76850 13694 76862 13746
rect 76914 13694 76926 13746
rect 75294 13682 75346 13694
rect 1822 13634 1874 13646
rect 5294 13634 5346 13646
rect 12798 13634 12850 13646
rect 3602 13582 3614 13634
rect 3666 13582 3678 13634
rect 7746 13582 7758 13634
rect 7810 13582 7822 13634
rect 1822 13570 1874 13582
rect 5294 13570 5346 13582
rect 12798 13570 12850 13582
rect 15262 13634 15314 13646
rect 15262 13570 15314 13582
rect 15710 13634 15762 13646
rect 15710 13570 15762 13582
rect 16158 13634 16210 13646
rect 26126 13634 26178 13646
rect 34078 13634 34130 13646
rect 20850 13582 20862 13634
rect 20914 13582 20926 13634
rect 28018 13582 28030 13634
rect 28082 13582 28094 13634
rect 16158 13570 16210 13582
rect 26126 13570 26178 13582
rect 34078 13570 34130 13582
rect 35758 13634 35810 13646
rect 35758 13570 35810 13582
rect 36318 13634 36370 13646
rect 36318 13570 36370 13582
rect 37214 13634 37266 13646
rect 59390 13634 59442 13646
rect 61966 13634 62018 13646
rect 39106 13582 39118 13634
rect 39170 13582 39182 13634
rect 44482 13582 44494 13634
rect 44546 13582 44558 13634
rect 49858 13582 49870 13634
rect 49922 13582 49934 13634
rect 60946 13582 60958 13634
rect 61010 13582 61022 13634
rect 37214 13570 37266 13582
rect 59390 13570 59442 13582
rect 61966 13570 62018 13582
rect 66110 13634 66162 13646
rect 66110 13570 66162 13582
rect 69806 13634 69858 13646
rect 69806 13570 69858 13582
rect 70366 13634 70418 13646
rect 70366 13570 70418 13582
rect 70814 13634 70866 13646
rect 70814 13570 70866 13582
rect 71374 13634 71426 13646
rect 71374 13570 71426 13582
rect 76190 13634 76242 13646
rect 76962 13582 76974 13634
rect 77026 13582 77038 13634
rect 76190 13570 76242 13582
rect 9886 13522 9938 13534
rect 9886 13458 9938 13470
rect 11678 13522 11730 13534
rect 54350 13522 54402 13534
rect 17602 13470 17614 13522
rect 17666 13519 17678 13522
rect 18162 13519 18174 13522
rect 17666 13473 18174 13519
rect 17666 13470 17678 13473
rect 18162 13470 18174 13473
rect 18226 13470 18238 13522
rect 11678 13458 11730 13470
rect 54350 13458 54402 13470
rect 61294 13522 61346 13534
rect 61294 13458 61346 13470
rect 75406 13522 75458 13534
rect 75406 13458 75458 13470
rect 1344 13354 78624 13388
rect 1344 13302 10874 13354
rect 10926 13302 10978 13354
rect 11030 13302 11082 13354
rect 11134 13302 30194 13354
rect 30246 13302 30298 13354
rect 30350 13302 30402 13354
rect 30454 13302 49514 13354
rect 49566 13302 49618 13354
rect 49670 13302 49722 13354
rect 49774 13302 68834 13354
rect 68886 13302 68938 13354
rect 68990 13302 69042 13354
rect 69094 13302 78624 13354
rect 1344 13268 78624 13302
rect 3390 13186 3442 13198
rect 3390 13122 3442 13134
rect 13806 13186 13858 13198
rect 13806 13122 13858 13134
rect 36654 13186 36706 13198
rect 42590 13186 42642 13198
rect 55358 13186 55410 13198
rect 77310 13186 77362 13198
rect 38322 13134 38334 13186
rect 38386 13134 38398 13186
rect 44258 13134 44270 13186
rect 44322 13134 44334 13186
rect 55682 13134 55694 13186
rect 55746 13134 55758 13186
rect 68450 13134 68462 13186
rect 68514 13134 68526 13186
rect 76402 13134 76414 13186
rect 76466 13134 76478 13186
rect 36654 13122 36706 13134
rect 42590 13122 42642 13134
rect 55358 13122 55410 13134
rect 77310 13122 77362 13134
rect 2830 13074 2882 13086
rect 2830 13010 2882 13022
rect 3614 13074 3666 13086
rect 3614 13010 3666 13022
rect 3950 13074 4002 13086
rect 3950 13010 4002 13022
rect 8990 13074 9042 13086
rect 14366 13074 14418 13086
rect 12338 13022 12350 13074
rect 12402 13022 12414 13074
rect 8990 13010 9042 13022
rect 14366 13010 14418 13022
rect 15262 13074 15314 13086
rect 17838 13074 17890 13086
rect 45950 13074 46002 13086
rect 17154 13022 17166 13074
rect 17218 13022 17230 13074
rect 25218 13022 25230 13074
rect 25282 13022 25294 13074
rect 32162 13022 32174 13074
rect 32226 13022 32238 13074
rect 37874 13022 37886 13074
rect 37938 13022 37950 13074
rect 43586 13022 43598 13074
rect 43650 13022 43662 13074
rect 15262 13010 15314 13022
rect 17838 13010 17890 13022
rect 45950 13010 46002 13022
rect 48974 13074 49026 13086
rect 48974 13010 49026 13022
rect 50990 13074 51042 13086
rect 54462 13074 54514 13086
rect 54338 13022 54350 13074
rect 54402 13022 54414 13074
rect 50990 13010 51042 13022
rect 54462 13010 54514 13022
rect 59278 13074 59330 13086
rect 59278 13010 59330 13022
rect 61518 13074 61570 13086
rect 61518 13010 61570 13022
rect 64430 13074 64482 13086
rect 66334 13074 66386 13086
rect 71710 13074 71762 13086
rect 65426 13022 65438 13074
rect 65490 13022 65502 13074
rect 67218 13022 67230 13074
rect 67282 13022 67294 13074
rect 64430 13010 64482 13022
rect 66334 13010 66386 13022
rect 71710 13010 71762 13022
rect 77870 13074 77922 13086
rect 77870 13010 77922 13022
rect 3838 12962 3890 12974
rect 3838 12898 3890 12910
rect 4062 12962 4114 12974
rect 4062 12898 4114 12910
rect 18398 12962 18450 12974
rect 18398 12898 18450 12910
rect 19070 12962 19122 12974
rect 19070 12898 19122 12910
rect 19406 12962 19458 12974
rect 20750 12962 20802 12974
rect 25902 12962 25954 12974
rect 39902 12962 39954 12974
rect 40798 12962 40850 12974
rect 20402 12910 20414 12962
rect 20466 12910 20478 12962
rect 24994 12910 25006 12962
rect 25058 12910 25070 12962
rect 32610 12910 32622 12962
rect 32674 12910 32686 12962
rect 33954 12910 33966 12962
rect 34018 12910 34030 12962
rect 37762 12910 37774 12962
rect 37826 12910 37838 12962
rect 40338 12910 40350 12962
rect 40402 12910 40414 12962
rect 19406 12898 19458 12910
rect 20750 12898 20802 12910
rect 25902 12898 25954 12910
rect 39902 12898 39954 12910
rect 40798 12898 40850 12910
rect 42478 12962 42530 12974
rect 45838 12962 45890 12974
rect 49870 12962 49922 12974
rect 55134 12962 55186 12974
rect 43474 12910 43486 12962
rect 43538 12910 43550 12962
rect 49634 12910 49646 12962
rect 49698 12910 49710 12962
rect 53778 12910 53790 12962
rect 53842 12910 53854 12962
rect 42478 12898 42530 12910
rect 45838 12898 45890 12910
rect 49870 12898 49922 12910
rect 55134 12898 55186 12910
rect 56142 12962 56194 12974
rect 60174 12962 60226 12974
rect 59938 12910 59950 12962
rect 60002 12910 60014 12962
rect 56142 12898 56194 12910
rect 60174 12898 60226 12910
rect 61294 12962 61346 12974
rect 61294 12898 61346 12910
rect 61854 12962 61906 12974
rect 64990 12962 65042 12974
rect 67902 12962 67954 12974
rect 63970 12910 63982 12962
rect 64034 12910 64046 12962
rect 66770 12910 66782 12962
rect 66834 12910 66846 12962
rect 61854 12898 61906 12910
rect 64990 12898 65042 12910
rect 67902 12898 67954 12910
rect 68126 12962 68178 12974
rect 68126 12898 68178 12910
rect 71150 12962 71202 12974
rect 71150 12898 71202 12910
rect 71374 12962 71426 12974
rect 71374 12898 71426 12910
rect 71822 12962 71874 12974
rect 76302 12962 76354 12974
rect 76066 12910 76078 12962
rect 76130 12910 76142 12962
rect 71822 12898 71874 12910
rect 76302 12898 76354 12910
rect 4846 12850 4898 12862
rect 4846 12786 4898 12798
rect 4958 12850 5010 12862
rect 4958 12786 5010 12798
rect 8430 12850 8482 12862
rect 8430 12786 8482 12798
rect 8542 12850 8594 12862
rect 8542 12786 8594 12798
rect 13694 12850 13746 12862
rect 13694 12786 13746 12798
rect 13806 12850 13858 12862
rect 13806 12786 13858 12798
rect 18510 12850 18562 12862
rect 18510 12786 18562 12798
rect 18734 12850 18786 12862
rect 18734 12786 18786 12798
rect 20302 12850 20354 12862
rect 20302 12786 20354 12798
rect 21646 12850 21698 12862
rect 21646 12786 21698 12798
rect 22094 12850 22146 12862
rect 22094 12786 22146 12798
rect 29598 12850 29650 12862
rect 36542 12850 36594 12862
rect 34178 12798 34190 12850
rect 34242 12798 34254 12850
rect 29598 12786 29650 12798
rect 36542 12786 36594 12798
rect 46062 12850 46114 12862
rect 46062 12786 46114 12798
rect 51102 12850 51154 12862
rect 51102 12786 51154 12798
rect 61742 12850 61794 12862
rect 61742 12786 61794 12798
rect 70142 12850 70194 12862
rect 70142 12786 70194 12798
rect 70254 12850 70306 12862
rect 70254 12786 70306 12798
rect 77422 12850 77474 12862
rect 77422 12786 77474 12798
rect 2046 12738 2098 12750
rect 2046 12674 2098 12686
rect 2494 12738 2546 12750
rect 2494 12674 2546 12686
rect 4622 12738 4674 12750
rect 4622 12674 4674 12686
rect 7758 12738 7810 12750
rect 7758 12674 7810 12686
rect 8206 12738 8258 12750
rect 8206 12674 8258 12686
rect 11790 12738 11842 12750
rect 11790 12674 11842 12686
rect 12798 12738 12850 12750
rect 12798 12674 12850 12686
rect 14814 12738 14866 12750
rect 14814 12674 14866 12686
rect 16158 12738 16210 12750
rect 16158 12674 16210 12686
rect 16718 12738 16770 12750
rect 16718 12674 16770 12686
rect 19294 12738 19346 12750
rect 19294 12674 19346 12686
rect 20078 12738 20130 12750
rect 20078 12674 20130 12686
rect 20190 12738 20242 12750
rect 20190 12674 20242 12686
rect 27358 12738 27410 12750
rect 27358 12674 27410 12686
rect 28030 12738 28082 12750
rect 28030 12674 28082 12686
rect 29710 12738 29762 12750
rect 29710 12674 29762 12686
rect 29934 12738 29986 12750
rect 29934 12674 29986 12686
rect 30270 12738 30322 12750
rect 30270 12674 30322 12686
rect 31502 12738 31554 12750
rect 31502 12674 31554 12686
rect 35534 12738 35586 12750
rect 35534 12674 35586 12686
rect 35982 12738 36034 12750
rect 35982 12674 36034 12686
rect 36654 12738 36706 12750
rect 36654 12674 36706 12686
rect 41918 12738 41970 12750
rect 41918 12674 41970 12686
rect 42590 12738 42642 12750
rect 42590 12674 42642 12686
rect 45614 12738 45666 12750
rect 45614 12674 45666 12686
rect 50654 12738 50706 12750
rect 50654 12674 50706 12686
rect 50878 12738 50930 12750
rect 50878 12674 50930 12686
rect 52670 12738 52722 12750
rect 52670 12674 52722 12686
rect 56926 12738 56978 12750
rect 56926 12674 56978 12686
rect 62414 12738 62466 12750
rect 62414 12674 62466 12686
rect 62862 12738 62914 12750
rect 62862 12674 62914 12686
rect 69246 12738 69298 12750
rect 69246 12674 69298 12686
rect 70478 12738 70530 12750
rect 70478 12674 70530 12686
rect 71598 12738 71650 12750
rect 71598 12674 71650 12686
rect 72382 12738 72434 12750
rect 72382 12674 72434 12686
rect 1344 12570 78784 12604
rect 1344 12518 20534 12570
rect 20586 12518 20638 12570
rect 20690 12518 20742 12570
rect 20794 12518 39854 12570
rect 39906 12518 39958 12570
rect 40010 12518 40062 12570
rect 40114 12518 59174 12570
rect 59226 12518 59278 12570
rect 59330 12518 59382 12570
rect 59434 12518 78494 12570
rect 78546 12518 78598 12570
rect 78650 12518 78702 12570
rect 78754 12518 78784 12570
rect 1344 12484 78784 12518
rect 8878 12402 8930 12414
rect 8878 12338 8930 12350
rect 16158 12402 16210 12414
rect 16158 12338 16210 12350
rect 17054 12402 17106 12414
rect 17054 12338 17106 12350
rect 18286 12402 18338 12414
rect 18286 12338 18338 12350
rect 19070 12402 19122 12414
rect 19070 12338 19122 12350
rect 19294 12402 19346 12414
rect 19294 12338 19346 12350
rect 19854 12402 19906 12414
rect 19854 12338 19906 12350
rect 21086 12402 21138 12414
rect 21086 12338 21138 12350
rect 22542 12402 22594 12414
rect 22542 12338 22594 12350
rect 23326 12402 23378 12414
rect 23326 12338 23378 12350
rect 37214 12402 37266 12414
rect 37214 12338 37266 12350
rect 42926 12402 42978 12414
rect 42926 12338 42978 12350
rect 48862 12402 48914 12414
rect 48862 12338 48914 12350
rect 53118 12402 53170 12414
rect 53118 12338 53170 12350
rect 55918 12402 55970 12414
rect 55918 12338 55970 12350
rect 56590 12402 56642 12414
rect 56590 12338 56642 12350
rect 58046 12402 58098 12414
rect 58046 12338 58098 12350
rect 58494 12402 58546 12414
rect 64654 12402 64706 12414
rect 61282 12350 61294 12402
rect 61346 12350 61358 12402
rect 58494 12338 58546 12350
rect 64654 12338 64706 12350
rect 65998 12402 66050 12414
rect 65998 12338 66050 12350
rect 73502 12402 73554 12414
rect 73502 12338 73554 12350
rect 74062 12402 74114 12414
rect 74062 12338 74114 12350
rect 6078 12290 6130 12302
rect 4162 12238 4174 12290
rect 4226 12238 4238 12290
rect 5842 12238 5854 12290
rect 5906 12238 5918 12290
rect 6078 12226 6130 12238
rect 8542 12290 8594 12302
rect 8542 12226 8594 12238
rect 11790 12290 11842 12302
rect 11790 12226 11842 12238
rect 12350 12290 12402 12302
rect 12350 12226 12402 12238
rect 12462 12290 12514 12302
rect 18174 12290 18226 12302
rect 13458 12238 13470 12290
rect 13522 12238 13534 12290
rect 12462 12226 12514 12238
rect 18174 12226 18226 12238
rect 20526 12290 20578 12302
rect 20526 12226 20578 12238
rect 22206 12290 22258 12302
rect 22206 12226 22258 12238
rect 22318 12290 22370 12302
rect 22318 12226 22370 12238
rect 26686 12290 26738 12302
rect 26686 12226 26738 12238
rect 30830 12290 30882 12302
rect 30830 12226 30882 12238
rect 34750 12290 34802 12302
rect 34750 12226 34802 12238
rect 48638 12290 48690 12302
rect 48638 12226 48690 12238
rect 53566 12290 53618 12302
rect 53566 12226 53618 12238
rect 55246 12290 55298 12302
rect 55246 12226 55298 12238
rect 57486 12290 57538 12302
rect 57486 12226 57538 12238
rect 60174 12290 60226 12302
rect 60174 12226 60226 12238
rect 61966 12290 62018 12302
rect 61966 12226 62018 12238
rect 62078 12290 62130 12302
rect 62078 12226 62130 12238
rect 62526 12290 62578 12302
rect 62526 12226 62578 12238
rect 63422 12290 63474 12302
rect 63422 12226 63474 12238
rect 66670 12290 66722 12302
rect 66670 12226 66722 12238
rect 66782 12290 66834 12302
rect 66782 12226 66834 12238
rect 68798 12290 68850 12302
rect 68798 12226 68850 12238
rect 71262 12290 71314 12302
rect 71262 12226 71314 12238
rect 76750 12290 76802 12302
rect 76750 12226 76802 12238
rect 8766 12178 8818 12190
rect 2930 12126 2942 12178
rect 2994 12126 3006 12178
rect 4498 12126 4510 12178
rect 4562 12126 4574 12178
rect 8766 12114 8818 12126
rect 8990 12178 9042 12190
rect 12686 12178 12738 12190
rect 16494 12178 16546 12190
rect 9986 12126 9998 12178
rect 10050 12126 10062 12178
rect 13794 12126 13806 12178
rect 13858 12126 13870 12178
rect 14802 12126 14814 12178
rect 14866 12126 14878 12178
rect 8990 12114 9042 12126
rect 12686 12114 12738 12126
rect 16494 12114 16546 12126
rect 18958 12178 19010 12190
rect 18958 12114 19010 12126
rect 20638 12178 20690 12190
rect 48526 12178 48578 12190
rect 54462 12178 54514 12190
rect 26002 12126 26014 12178
rect 26066 12126 26078 12178
rect 27906 12126 27918 12178
rect 27970 12126 27982 12178
rect 28802 12126 28814 12178
rect 28866 12126 28878 12178
rect 30034 12126 30046 12178
rect 30098 12126 30110 12178
rect 34178 12126 34190 12178
rect 34242 12126 34254 12178
rect 39218 12126 39230 12178
rect 39282 12126 39294 12178
rect 43810 12126 43822 12178
rect 43874 12126 43886 12178
rect 49746 12126 49758 12178
rect 49810 12126 49822 12178
rect 54002 12126 54014 12178
rect 54066 12126 54078 12178
rect 20638 12114 20690 12126
rect 48526 12114 48578 12126
rect 54462 12114 54514 12126
rect 56478 12178 56530 12190
rect 56478 12114 56530 12126
rect 56814 12178 56866 12190
rect 63198 12178 63250 12190
rect 59490 12126 59502 12178
rect 59554 12126 59566 12178
rect 56814 12114 56866 12126
rect 63198 12114 63250 12126
rect 63534 12178 63586 12190
rect 63534 12114 63586 12126
rect 67006 12178 67058 12190
rect 67006 12114 67058 12126
rect 67678 12178 67730 12190
rect 67678 12114 67730 12126
rect 68238 12178 68290 12190
rect 73390 12178 73442 12190
rect 70466 12126 70478 12178
rect 70530 12126 70542 12178
rect 68238 12114 68290 12126
rect 73390 12114 73442 12126
rect 73726 12178 73778 12190
rect 76178 12126 76190 12178
rect 76242 12126 76254 12178
rect 77186 12126 77198 12178
rect 77250 12126 77262 12178
rect 73726 12114 73778 12126
rect 15374 12066 15426 12078
rect 1922 12014 1934 12066
rect 1986 12014 1998 12066
rect 10098 12014 10110 12066
rect 10162 12014 10174 12066
rect 15374 12002 15426 12014
rect 17614 12066 17666 12078
rect 17614 12002 17666 12014
rect 21534 12066 21586 12078
rect 21534 12002 21586 12014
rect 22878 12066 22930 12078
rect 22878 12002 22930 12014
rect 24894 12066 24946 12078
rect 35982 12066 36034 12078
rect 25778 12014 25790 12066
rect 25842 12014 25854 12066
rect 28578 12014 28590 12066
rect 28642 12014 28654 12066
rect 34402 12014 34414 12066
rect 34466 12014 34478 12066
rect 24894 12002 24946 12014
rect 35982 12002 36034 12014
rect 38558 12066 38610 12078
rect 42590 12066 42642 12078
rect 55134 12066 55186 12078
rect 60734 12066 60786 12078
rect 39554 12014 39566 12066
rect 39618 12014 39630 12066
rect 44146 12014 44158 12066
rect 44210 12014 44222 12066
rect 49858 12014 49870 12066
rect 49922 12014 49934 12066
rect 59714 12014 59726 12066
rect 59778 12014 59790 12066
rect 38558 12002 38610 12014
rect 42590 12002 42642 12014
rect 55134 12002 55186 12014
rect 60734 12002 60786 12014
rect 63982 12066 64034 12078
rect 69582 12066 69634 12078
rect 65538 12014 65550 12066
rect 65602 12014 65614 12066
rect 70354 12014 70366 12066
rect 70418 12014 70430 12066
rect 75506 12014 75518 12066
rect 75570 12014 75582 12066
rect 77522 12014 77534 12066
rect 77586 12014 77598 12066
rect 63982 12002 64034 12014
rect 69582 12002 69634 12014
rect 18286 11954 18338 11966
rect 10770 11902 10782 11954
rect 10834 11902 10846 11954
rect 18286 11890 18338 11902
rect 20526 11954 20578 11966
rect 20526 11890 20578 11902
rect 27582 11954 27634 11966
rect 27582 11890 27634 11902
rect 27918 11954 27970 11966
rect 60958 11954 61010 11966
rect 39666 11902 39678 11954
rect 39730 11902 39742 11954
rect 44482 11902 44494 11954
rect 44546 11902 44558 11954
rect 50082 11902 50094 11954
rect 50146 11902 50158 11954
rect 27918 11890 27970 11902
rect 60958 11890 61010 11902
rect 61966 11954 62018 11966
rect 61966 11890 62018 11902
rect 1344 11786 78624 11820
rect 1344 11734 10874 11786
rect 10926 11734 10978 11786
rect 11030 11734 11082 11786
rect 11134 11734 30194 11786
rect 30246 11734 30298 11786
rect 30350 11734 30402 11786
rect 30454 11734 49514 11786
rect 49566 11734 49618 11786
rect 49670 11734 49722 11786
rect 49774 11734 68834 11786
rect 68886 11734 68938 11786
rect 68990 11734 69042 11786
rect 69094 11734 78624 11786
rect 1344 11700 78624 11734
rect 13694 11618 13746 11630
rect 8978 11566 8990 11618
rect 9042 11566 9054 11618
rect 13694 11554 13746 11566
rect 44270 11618 44322 11630
rect 44270 11554 44322 11566
rect 70030 11618 70082 11630
rect 71250 11566 71262 11618
rect 71314 11566 71326 11618
rect 70030 11554 70082 11566
rect 2046 11506 2098 11518
rect 13022 11506 13074 11518
rect 3266 11454 3278 11506
rect 3330 11454 3342 11506
rect 5730 11454 5742 11506
rect 5794 11454 5806 11506
rect 8642 11454 8654 11506
rect 8706 11454 8718 11506
rect 2046 11442 2098 11454
rect 13022 11442 13074 11454
rect 16158 11506 16210 11518
rect 21646 11506 21698 11518
rect 18610 11454 18622 11506
rect 18674 11454 18686 11506
rect 20850 11454 20862 11506
rect 20914 11454 20926 11506
rect 16158 11442 16210 11454
rect 21646 11442 21698 11454
rect 21870 11506 21922 11518
rect 26798 11506 26850 11518
rect 24994 11454 25006 11506
rect 25058 11454 25070 11506
rect 21870 11442 21922 11454
rect 26798 11442 26850 11454
rect 29710 11506 29762 11518
rect 29710 11442 29762 11454
rect 34302 11506 34354 11518
rect 34302 11442 34354 11454
rect 36206 11506 36258 11518
rect 36206 11442 36258 11454
rect 43598 11506 43650 11518
rect 56366 11506 56418 11518
rect 57934 11506 57986 11518
rect 63310 11506 63362 11518
rect 66222 11506 66274 11518
rect 52322 11454 52334 11506
rect 52386 11454 52398 11506
rect 54226 11454 54238 11506
rect 54290 11454 54302 11506
rect 57250 11454 57262 11506
rect 57314 11454 57326 11506
rect 62290 11454 62302 11506
rect 62354 11454 62366 11506
rect 63746 11454 63758 11506
rect 63810 11454 63822 11506
rect 43598 11442 43650 11454
rect 56366 11442 56418 11454
rect 57934 11442 57986 11454
rect 63310 11442 63362 11454
rect 66222 11442 66274 11454
rect 66558 11506 66610 11518
rect 66558 11442 66610 11454
rect 67006 11506 67058 11518
rect 67006 11442 67058 11454
rect 67454 11506 67506 11518
rect 74846 11506 74898 11518
rect 71138 11454 71150 11506
rect 71202 11454 71214 11506
rect 67454 11442 67506 11454
rect 74846 11442 74898 11454
rect 76526 11506 76578 11518
rect 76526 11442 76578 11454
rect 77422 11506 77474 11518
rect 77422 11442 77474 11454
rect 3614 11394 3666 11406
rect 3154 11342 3166 11394
rect 3218 11342 3230 11394
rect 3614 11330 3666 11342
rect 4174 11394 4226 11406
rect 4174 11330 4226 11342
rect 4510 11394 4562 11406
rect 4510 11330 4562 11342
rect 4734 11394 4786 11406
rect 13918 11394 13970 11406
rect 8754 11342 8766 11394
rect 8818 11342 8830 11394
rect 4734 11330 4786 11342
rect 13918 11330 13970 11342
rect 14142 11394 14194 11406
rect 14142 11330 14194 11342
rect 14254 11394 14306 11406
rect 14254 11330 14306 11342
rect 15262 11394 15314 11406
rect 15262 11330 15314 11342
rect 18062 11394 18114 11406
rect 22094 11394 22146 11406
rect 18946 11342 18958 11394
rect 19010 11342 19022 11394
rect 20178 11342 20190 11394
rect 20242 11342 20254 11394
rect 18062 11330 18114 11342
rect 22094 11330 22146 11342
rect 22206 11394 22258 11406
rect 25790 11394 25842 11406
rect 24882 11342 24894 11394
rect 24946 11342 24958 11394
rect 22206 11330 22258 11342
rect 25790 11330 25842 11342
rect 26238 11394 26290 11406
rect 26238 11330 26290 11342
rect 26686 11394 26738 11406
rect 26686 11330 26738 11342
rect 26910 11394 26962 11406
rect 26910 11330 26962 11342
rect 29598 11394 29650 11406
rect 29598 11330 29650 11342
rect 33742 11394 33794 11406
rect 33742 11330 33794 11342
rect 34190 11394 34242 11406
rect 34190 11330 34242 11342
rect 34414 11394 34466 11406
rect 34414 11330 34466 11342
rect 35534 11394 35586 11406
rect 35534 11330 35586 11342
rect 40014 11394 40066 11406
rect 40014 11330 40066 11342
rect 44158 11394 44210 11406
rect 44158 11330 44210 11342
rect 48862 11394 48914 11406
rect 48862 11330 48914 11342
rect 49310 11394 49362 11406
rect 49310 11330 49362 11342
rect 51550 11394 51602 11406
rect 70142 11394 70194 11406
rect 73838 11394 73890 11406
rect 51986 11342 51998 11394
rect 52050 11342 52062 11394
rect 54114 11342 54126 11394
rect 54178 11342 54190 11394
rect 57026 11342 57038 11394
rect 57090 11342 57102 11394
rect 58258 11342 58270 11394
rect 58322 11342 58334 11394
rect 62178 11342 62190 11394
rect 62242 11342 62254 11394
rect 63858 11342 63870 11394
rect 63922 11342 63934 11394
rect 71362 11342 71374 11394
rect 71426 11342 71438 11394
rect 51550 11330 51602 11342
rect 70142 11330 70194 11342
rect 73838 11330 73890 11342
rect 74958 11394 75010 11406
rect 74958 11330 75010 11342
rect 75630 11394 75682 11406
rect 77758 11394 77810 11406
rect 75842 11342 75854 11394
rect 75906 11342 75918 11394
rect 75630 11330 75682 11342
rect 77758 11330 77810 11342
rect 5854 11282 5906 11294
rect 5854 11218 5906 11230
rect 6078 11282 6130 11294
rect 6078 11218 6130 11230
rect 16718 11282 16770 11294
rect 16718 11218 16770 11230
rect 17726 11282 17778 11294
rect 17726 11218 17778 11230
rect 30046 11282 30098 11294
rect 30046 11218 30098 11230
rect 39678 11282 39730 11294
rect 39678 11218 39730 11230
rect 40574 11282 40626 11294
rect 40574 11218 40626 11230
rect 48750 11282 48802 11294
rect 48750 11218 48802 11230
rect 53454 11282 53506 11294
rect 53454 11218 53506 11230
rect 58942 11282 58994 11294
rect 58942 11218 58994 11230
rect 60510 11282 60562 11294
rect 60510 11218 60562 11230
rect 61518 11282 61570 11294
rect 61518 11218 61570 11230
rect 77310 11282 77362 11294
rect 77310 11218 77362 11230
rect 77646 11282 77698 11294
rect 77646 11218 77698 11230
rect 4622 11170 4674 11182
rect 4622 11106 4674 11118
rect 12014 11170 12066 11182
rect 12014 11106 12066 11118
rect 12462 11170 12514 11182
rect 12462 11106 12514 11118
rect 14366 11170 14418 11182
rect 14366 11106 14418 11118
rect 14926 11170 14978 11182
rect 14926 11106 14978 11118
rect 15150 11170 15202 11182
rect 15150 11106 15202 11118
rect 15710 11170 15762 11182
rect 15710 11106 15762 11118
rect 17278 11170 17330 11182
rect 17278 11106 17330 11118
rect 17838 11170 17890 11182
rect 17838 11106 17890 11118
rect 22318 11170 22370 11182
rect 22318 11106 22370 11118
rect 28142 11170 28194 11182
rect 28142 11106 28194 11118
rect 28814 11170 28866 11182
rect 28814 11106 28866 11118
rect 29822 11170 29874 11182
rect 29822 11106 29874 11118
rect 31054 11170 31106 11182
rect 31054 11106 31106 11118
rect 34974 11170 35026 11182
rect 34974 11106 35026 11118
rect 35646 11170 35698 11182
rect 35646 11106 35698 11118
rect 35870 11170 35922 11182
rect 35870 11106 35922 11118
rect 39118 11170 39170 11182
rect 39118 11106 39170 11118
rect 39790 11170 39842 11182
rect 39790 11106 39842 11118
rect 40462 11170 40514 11182
rect 40462 11106 40514 11118
rect 41022 11170 41074 11182
rect 41022 11106 41074 11118
rect 44270 11170 44322 11182
rect 44270 11106 44322 11118
rect 48638 11170 48690 11182
rect 48638 11106 48690 11118
rect 50990 11170 51042 11182
rect 50990 11106 51042 11118
rect 55022 11170 55074 11182
rect 55022 11106 55074 11118
rect 58046 11170 58098 11182
rect 58046 11106 58098 11118
rect 64766 11170 64818 11182
rect 64766 11106 64818 11118
rect 69470 11170 69522 11182
rect 69470 11106 69522 11118
rect 70030 11170 70082 11182
rect 70030 11106 70082 11118
rect 72270 11170 72322 11182
rect 72270 11106 72322 11118
rect 74510 11170 74562 11182
rect 74510 11106 74562 11118
rect 74734 11170 74786 11182
rect 74734 11106 74786 11118
rect 1344 11002 78784 11036
rect 1344 10950 20534 11002
rect 20586 10950 20638 11002
rect 20690 10950 20742 11002
rect 20794 10950 39854 11002
rect 39906 10950 39958 11002
rect 40010 10950 40062 11002
rect 40114 10950 59174 11002
rect 59226 10950 59278 11002
rect 59330 10950 59382 11002
rect 59434 10950 78494 11002
rect 78546 10950 78598 11002
rect 78650 10950 78702 11002
rect 78754 10950 78784 11002
rect 1344 10916 78784 10950
rect 2830 10834 2882 10846
rect 8766 10834 8818 10846
rect 3826 10782 3838 10834
rect 3890 10782 3902 10834
rect 2830 10770 2882 10782
rect 8766 10770 8818 10782
rect 10558 10834 10610 10846
rect 10558 10770 10610 10782
rect 11342 10834 11394 10846
rect 11342 10770 11394 10782
rect 12798 10834 12850 10846
rect 12798 10770 12850 10782
rect 13358 10834 13410 10846
rect 13358 10770 13410 10782
rect 13582 10834 13634 10846
rect 13582 10770 13634 10782
rect 14926 10834 14978 10846
rect 14926 10770 14978 10782
rect 15934 10834 15986 10846
rect 15934 10770 15986 10782
rect 17614 10834 17666 10846
rect 17614 10770 17666 10782
rect 18622 10834 18674 10846
rect 18622 10770 18674 10782
rect 20638 10834 20690 10846
rect 20638 10770 20690 10782
rect 21310 10834 21362 10846
rect 21310 10770 21362 10782
rect 25790 10834 25842 10846
rect 25790 10770 25842 10782
rect 26014 10834 26066 10846
rect 26014 10770 26066 10782
rect 26462 10834 26514 10846
rect 26462 10770 26514 10782
rect 30830 10834 30882 10846
rect 30830 10770 30882 10782
rect 45390 10834 45442 10846
rect 45390 10770 45442 10782
rect 49422 10834 49474 10846
rect 49422 10770 49474 10782
rect 52446 10834 52498 10846
rect 52446 10770 52498 10782
rect 53006 10834 53058 10846
rect 53006 10770 53058 10782
rect 53118 10834 53170 10846
rect 53118 10770 53170 10782
rect 55806 10834 55858 10846
rect 55806 10770 55858 10782
rect 56478 10834 56530 10846
rect 56478 10770 56530 10782
rect 57710 10834 57762 10846
rect 57710 10770 57762 10782
rect 62302 10834 62354 10846
rect 62302 10770 62354 10782
rect 63086 10834 63138 10846
rect 63086 10770 63138 10782
rect 63534 10834 63586 10846
rect 63534 10770 63586 10782
rect 69358 10834 69410 10846
rect 69358 10770 69410 10782
rect 70478 10834 70530 10846
rect 70478 10770 70530 10782
rect 70814 10834 70866 10846
rect 70814 10770 70866 10782
rect 2606 10722 2658 10734
rect 2606 10658 2658 10670
rect 7870 10722 7922 10734
rect 7870 10658 7922 10670
rect 8654 10722 8706 10734
rect 8654 10658 8706 10670
rect 12462 10722 12514 10734
rect 12462 10658 12514 10670
rect 12574 10722 12626 10734
rect 12574 10658 12626 10670
rect 18174 10722 18226 10734
rect 18174 10658 18226 10670
rect 21534 10722 21586 10734
rect 21534 10658 21586 10670
rect 24334 10722 24386 10734
rect 24334 10658 24386 10670
rect 25678 10722 25730 10734
rect 25678 10658 25730 10670
rect 30494 10722 30546 10734
rect 30494 10658 30546 10670
rect 30606 10722 30658 10734
rect 30606 10658 30658 10670
rect 32958 10722 33010 10734
rect 32958 10658 33010 10670
rect 44382 10722 44434 10734
rect 44382 10658 44434 10670
rect 49646 10722 49698 10734
rect 49646 10658 49698 10670
rect 53230 10722 53282 10734
rect 53230 10658 53282 10670
rect 54238 10722 54290 10734
rect 54238 10658 54290 10670
rect 54350 10722 54402 10734
rect 54350 10658 54402 10670
rect 57822 10722 57874 10734
rect 57822 10658 57874 10670
rect 61966 10722 62018 10734
rect 61966 10658 62018 10670
rect 66670 10722 66722 10734
rect 66670 10658 66722 10670
rect 69470 10722 69522 10734
rect 69470 10658 69522 10670
rect 70142 10722 70194 10734
rect 70142 10658 70194 10670
rect 70254 10722 70306 10734
rect 70254 10658 70306 10670
rect 75742 10722 75794 10734
rect 75742 10658 75794 10670
rect 77982 10722 78034 10734
rect 77982 10658 78034 10670
rect 2494 10610 2546 10622
rect 2494 10546 2546 10558
rect 3278 10610 3330 10622
rect 3278 10546 3330 10558
rect 4398 10610 4450 10622
rect 6414 10610 6466 10622
rect 11118 10610 11170 10622
rect 6066 10558 6078 10610
rect 6130 10558 6142 10610
rect 7410 10558 7422 10610
rect 7474 10558 7486 10610
rect 4398 10546 4450 10558
rect 6414 10546 6466 10558
rect 11118 10546 11170 10558
rect 11230 10610 11282 10622
rect 13470 10610 13522 10622
rect 11666 10558 11678 10610
rect 11730 10558 11742 10610
rect 11230 10546 11282 10558
rect 13470 10546 13522 10558
rect 13694 10610 13746 10622
rect 14366 10610 14418 10622
rect 13906 10558 13918 10610
rect 13970 10558 13982 10610
rect 13694 10546 13746 10558
rect 14366 10546 14418 10558
rect 15486 10610 15538 10622
rect 15486 10546 15538 10558
rect 17054 10610 17106 10622
rect 17054 10546 17106 10558
rect 18398 10610 18450 10622
rect 18398 10546 18450 10558
rect 18734 10610 18786 10622
rect 19966 10610 20018 10622
rect 19506 10558 19518 10610
rect 19570 10558 19582 10610
rect 18734 10546 18786 10558
rect 19966 10546 20018 10558
rect 21198 10610 21250 10622
rect 28254 10610 28306 10622
rect 32398 10610 32450 10622
rect 35422 10610 35474 10622
rect 39230 10610 39282 10622
rect 40798 10610 40850 10622
rect 44830 10610 44882 10622
rect 22306 10558 22318 10610
rect 22370 10558 22382 10610
rect 23538 10558 23550 10610
rect 23602 10558 23614 10610
rect 29474 10558 29486 10610
rect 29538 10558 29550 10610
rect 31490 10558 31502 10610
rect 31554 10558 31566 10610
rect 33842 10558 33854 10610
rect 33906 10558 33918 10610
rect 35858 10558 35870 10610
rect 35922 10558 35934 10610
rect 38322 10558 38334 10610
rect 38386 10558 38398 10610
rect 40114 10558 40126 10610
rect 40178 10558 40190 10610
rect 42802 10558 42814 10610
rect 42866 10558 42878 10610
rect 43810 10558 43822 10610
rect 43874 10558 43886 10610
rect 21198 10546 21250 10558
rect 28254 10546 28306 10558
rect 32398 10546 32450 10558
rect 35422 10546 35474 10558
rect 39230 10546 39282 10558
rect 40798 10546 40850 10558
rect 44830 10546 44882 10558
rect 45278 10610 45330 10622
rect 45278 10546 45330 10558
rect 45502 10610 45554 10622
rect 47294 10610 47346 10622
rect 49758 10610 49810 10622
rect 46946 10558 46958 10610
rect 47010 10558 47022 10610
rect 48290 10558 48302 10610
rect 48354 10558 48366 10610
rect 45502 10546 45554 10558
rect 47294 10546 47346 10558
rect 49758 10546 49810 10558
rect 53678 10610 53730 10622
rect 53678 10546 53730 10558
rect 54014 10610 54066 10622
rect 54014 10546 54066 10558
rect 54798 10610 54850 10622
rect 54798 10546 54850 10558
rect 56590 10610 56642 10622
rect 62190 10610 62242 10622
rect 57474 10558 57486 10610
rect 57538 10558 57550 10610
rect 56590 10546 56642 10558
rect 62190 10546 62242 10558
rect 62414 10610 62466 10622
rect 62414 10546 62466 10558
rect 63310 10610 63362 10622
rect 63310 10546 63362 10558
rect 63422 10610 63474 10622
rect 63422 10546 63474 10558
rect 65550 10610 65602 10622
rect 76414 10610 76466 10622
rect 78094 10610 78146 10622
rect 65986 10558 65998 10610
rect 66050 10558 66062 10610
rect 67330 10558 67342 10610
rect 67394 10558 67406 10610
rect 68562 10558 68574 10610
rect 68626 10558 68638 10610
rect 72146 10558 72158 10610
rect 72210 10558 72222 10610
rect 73714 10558 73726 10610
rect 73778 10558 73790 10610
rect 74834 10558 74846 10610
rect 74898 10558 74910 10610
rect 76738 10558 76750 10610
rect 76802 10558 76814 10610
rect 65550 10546 65602 10558
rect 76414 10546 76466 10558
rect 78094 10546 78146 10558
rect 1934 10498 1986 10510
rect 1934 10434 1986 10446
rect 10446 10498 10498 10510
rect 10446 10434 10498 10446
rect 16606 10498 16658 10510
rect 16606 10434 16658 10446
rect 18510 10498 18562 10510
rect 29822 10498 29874 10510
rect 36318 10498 36370 10510
rect 22082 10446 22094 10498
rect 22146 10446 22158 10498
rect 27794 10446 27806 10498
rect 27858 10446 27870 10498
rect 29362 10446 29374 10498
rect 29426 10446 29438 10498
rect 31826 10446 31838 10498
rect 31890 10446 31902 10498
rect 33954 10446 33966 10498
rect 34018 10446 34030 10498
rect 18510 10434 18562 10446
rect 29822 10434 29874 10446
rect 36318 10434 36370 10446
rect 36878 10498 36930 10510
rect 41470 10498 41522 10510
rect 50318 10498 50370 10510
rect 38658 10446 38670 10498
rect 38722 10446 38734 10498
rect 40002 10446 40014 10498
rect 40066 10446 40078 10498
rect 44034 10446 44046 10498
rect 44098 10446 44110 10498
rect 36878 10434 36930 10446
rect 41470 10434 41522 10446
rect 50318 10434 50370 10446
rect 56702 10498 56754 10510
rect 56702 10434 56754 10446
rect 58382 10498 58434 10510
rect 58382 10434 58434 10446
rect 64654 10498 64706 10510
rect 72494 10498 72546 10510
rect 67554 10446 67566 10498
rect 67618 10446 67630 10498
rect 71810 10446 71822 10498
rect 71874 10446 71886 10498
rect 64654 10434 64706 10446
rect 72494 10434 72546 10446
rect 73390 10498 73442 10510
rect 73390 10434 73442 10446
rect 73502 10498 73554 10510
rect 76302 10498 76354 10510
rect 74946 10446 74958 10498
rect 75010 10446 75022 10498
rect 73502 10434 73554 10446
rect 76302 10434 76354 10446
rect 3502 10386 3554 10398
rect 3502 10322 3554 10334
rect 4622 10386 4674 10398
rect 8766 10386 8818 10398
rect 42478 10386 42530 10398
rect 4946 10334 4958 10386
rect 5010 10334 5022 10386
rect 14130 10334 14142 10386
rect 14194 10383 14206 10386
rect 14690 10383 14702 10386
rect 14194 10337 14702 10383
rect 14194 10334 14206 10337
rect 14690 10334 14702 10337
rect 14754 10334 14766 10386
rect 34402 10334 34414 10386
rect 34466 10334 34478 10386
rect 4622 10322 4674 10334
rect 8766 10322 8818 10334
rect 42478 10322 42530 10334
rect 42814 10386 42866 10398
rect 68238 10386 68290 10398
rect 48402 10334 48414 10386
rect 48466 10334 48478 10386
rect 42814 10322 42866 10334
rect 68238 10322 68290 10334
rect 68574 10386 68626 10398
rect 68574 10322 68626 10334
rect 69246 10386 69298 10398
rect 69246 10322 69298 10334
rect 77982 10386 78034 10398
rect 77982 10322 78034 10334
rect 1344 10218 78624 10252
rect 1344 10166 10874 10218
rect 10926 10166 10978 10218
rect 11030 10166 11082 10218
rect 11134 10166 30194 10218
rect 30246 10166 30298 10218
rect 30350 10166 30402 10218
rect 30454 10166 49514 10218
rect 49566 10166 49618 10218
rect 49670 10166 49722 10218
rect 49774 10166 68834 10218
rect 68886 10166 68938 10218
rect 68990 10166 69042 10218
rect 69094 10166 78624 10218
rect 1344 10132 78624 10166
rect 4510 10050 4562 10062
rect 4510 9986 4562 9998
rect 7646 10050 7698 10062
rect 7646 9986 7698 9998
rect 17390 10050 17442 10062
rect 17390 9986 17442 9998
rect 19518 10050 19570 10062
rect 19518 9986 19570 9998
rect 35534 10050 35586 10062
rect 35534 9986 35586 9998
rect 43150 10050 43202 10062
rect 43150 9986 43202 9998
rect 44606 10050 44658 10062
rect 62414 10050 62466 10062
rect 57250 9998 57262 10050
rect 57314 9998 57326 10050
rect 44606 9986 44658 9998
rect 62414 9986 62466 9998
rect 63422 10050 63474 10062
rect 72046 10050 72098 10062
rect 67554 9998 67566 10050
rect 67618 9998 67630 10050
rect 63422 9986 63474 9998
rect 72046 9986 72098 9998
rect 73278 10050 73330 10062
rect 73278 9986 73330 9998
rect 76526 10050 76578 10062
rect 77634 9998 77646 10050
rect 77698 10047 77710 10050
rect 77858 10047 77870 10050
rect 77698 10001 77870 10047
rect 77698 9998 77710 10001
rect 77858 9998 77870 10001
rect 77922 9998 77934 10050
rect 76526 9986 76578 9998
rect 7870 9938 7922 9950
rect 3714 9886 3726 9938
rect 3778 9886 3790 9938
rect 7870 9874 7922 9886
rect 8206 9938 8258 9950
rect 12574 9938 12626 9950
rect 15598 9938 15650 9950
rect 11330 9886 11342 9938
rect 11394 9886 11406 9938
rect 15026 9886 15038 9938
rect 15090 9886 15102 9938
rect 8206 9874 8258 9886
rect 12574 9874 12626 9886
rect 15598 9874 15650 9886
rect 18846 9938 18898 9950
rect 18846 9874 18898 9886
rect 20750 9938 20802 9950
rect 20750 9874 20802 9886
rect 21646 9938 21698 9950
rect 21646 9874 21698 9886
rect 22318 9938 22370 9950
rect 22318 9874 22370 9886
rect 26910 9938 26962 9950
rect 26910 9874 26962 9886
rect 30270 9938 30322 9950
rect 30270 9874 30322 9886
rect 30942 9938 30994 9950
rect 30942 9874 30994 9886
rect 32286 9938 32338 9950
rect 68350 9938 68402 9950
rect 74958 9938 75010 9950
rect 35746 9886 35758 9938
rect 35810 9886 35822 9938
rect 48514 9886 48526 9938
rect 48578 9886 48590 9938
rect 65538 9886 65550 9938
rect 65602 9886 65614 9938
rect 67218 9886 67230 9938
rect 67282 9886 67294 9938
rect 69458 9886 69470 9938
rect 69522 9886 69534 9938
rect 72370 9886 72382 9938
rect 72434 9886 72446 9938
rect 32286 9874 32338 9886
rect 68350 9874 68402 9886
rect 74958 9874 75010 9886
rect 76414 9938 76466 9950
rect 76414 9874 76466 9886
rect 77982 9938 78034 9950
rect 77982 9874 78034 9886
rect 4622 9826 4674 9838
rect 4622 9762 4674 9774
rect 5630 9826 5682 9838
rect 5630 9762 5682 9774
rect 8094 9826 8146 9838
rect 8094 9762 8146 9774
rect 8878 9826 8930 9838
rect 11678 9826 11730 9838
rect 10994 9774 11006 9826
rect 11058 9774 11070 9826
rect 8878 9762 8930 9774
rect 11678 9762 11730 9774
rect 13694 9826 13746 9838
rect 13694 9762 13746 9774
rect 18398 9826 18450 9838
rect 22878 9826 22930 9838
rect 18498 9774 18510 9826
rect 18562 9774 18574 9826
rect 18398 9762 18450 9774
rect 22878 9762 22930 9774
rect 25454 9826 25506 9838
rect 25454 9762 25506 9774
rect 26014 9826 26066 9838
rect 28478 9826 28530 9838
rect 26226 9774 26238 9826
rect 26290 9774 26302 9826
rect 26014 9762 26066 9774
rect 28478 9762 28530 9774
rect 29934 9826 29986 9838
rect 29934 9762 29986 9774
rect 33518 9826 33570 9838
rect 36430 9826 36482 9838
rect 35858 9774 35870 9826
rect 35922 9774 35934 9826
rect 33518 9762 33570 9774
rect 36430 9762 36482 9774
rect 38558 9826 38610 9838
rect 38558 9762 38610 9774
rect 38894 9826 38946 9838
rect 38894 9762 38946 9774
rect 39454 9826 39506 9838
rect 39454 9762 39506 9774
rect 39902 9826 39954 9838
rect 39902 9762 39954 9774
rect 40126 9826 40178 9838
rect 40126 9762 40178 9774
rect 41134 9826 41186 9838
rect 41134 9762 41186 9774
rect 41358 9826 41410 9838
rect 41358 9762 41410 9774
rect 44718 9826 44770 9838
rect 44718 9762 44770 9774
rect 45502 9826 45554 9838
rect 45502 9762 45554 9774
rect 45726 9826 45778 9838
rect 49758 9826 49810 9838
rect 45938 9774 45950 9826
rect 46002 9774 46014 9826
rect 48626 9774 48638 9826
rect 48690 9774 48702 9826
rect 45726 9762 45778 9774
rect 49758 9762 49810 9774
rect 49982 9826 50034 9838
rect 49982 9762 50034 9774
rect 51550 9826 51602 9838
rect 57374 9826 57426 9838
rect 69694 9826 69746 9838
rect 56690 9774 56702 9826
rect 56754 9774 56766 9826
rect 62402 9774 62414 9826
rect 62466 9774 62478 9826
rect 66994 9774 67006 9826
rect 67058 9774 67070 9826
rect 51550 9762 51602 9774
rect 57374 9762 57426 9774
rect 69694 9762 69746 9774
rect 70590 9826 70642 9838
rect 70590 9762 70642 9774
rect 71038 9826 71090 9838
rect 71038 9762 71090 9774
rect 71374 9826 71426 9838
rect 72930 9774 72942 9826
rect 72994 9774 73006 9826
rect 71374 9762 71426 9774
rect 2382 9714 2434 9726
rect 2382 9650 2434 9662
rect 5966 9714 6018 9726
rect 5966 9650 6018 9662
rect 17278 9714 17330 9726
rect 17278 9650 17330 9662
rect 18174 9714 18226 9726
rect 18174 9650 18226 9662
rect 19406 9714 19458 9726
rect 19406 9650 19458 9662
rect 19518 9714 19570 9726
rect 19518 9650 19570 9662
rect 23662 9714 23714 9726
rect 23662 9650 23714 9662
rect 29598 9714 29650 9726
rect 29598 9650 29650 9662
rect 33182 9714 33234 9726
rect 33182 9650 33234 9662
rect 34974 9714 35026 9726
rect 34974 9650 35026 9662
rect 36542 9714 36594 9726
rect 36542 9650 36594 9662
rect 43486 9714 43538 9726
rect 43486 9650 43538 9662
rect 44606 9714 44658 9726
rect 44606 9650 44658 9662
rect 48302 9714 48354 9726
rect 48302 9650 48354 9662
rect 50878 9714 50930 9726
rect 50878 9650 50930 9662
rect 50990 9714 51042 9726
rect 50990 9650 51042 9662
rect 59950 9714 60002 9726
rect 59950 9650 60002 9662
rect 62750 9714 62802 9726
rect 62750 9650 62802 9662
rect 63422 9714 63474 9726
rect 63422 9650 63474 9662
rect 63534 9714 63586 9726
rect 63534 9650 63586 9662
rect 70254 9714 70306 9726
rect 70254 9650 70306 9662
rect 71150 9714 71202 9726
rect 71150 9650 71202 9662
rect 72270 9714 72322 9726
rect 73166 9714 73218 9726
rect 73726 9714 73778 9726
rect 72482 9662 72494 9714
rect 72546 9711 72558 9714
rect 72818 9711 72830 9714
rect 72546 9665 72830 9711
rect 72546 9662 72558 9665
rect 72818 9662 72830 9665
rect 72882 9662 72894 9714
rect 73378 9662 73390 9714
rect 73442 9711 73454 9714
rect 73602 9711 73614 9714
rect 73442 9665 73614 9711
rect 73442 9662 73454 9665
rect 73602 9662 73614 9665
rect 73666 9662 73678 9714
rect 72270 9650 72322 9662
rect 73166 9650 73218 9662
rect 73726 9650 73778 9662
rect 1934 9602 1986 9614
rect 1934 9538 1986 9550
rect 2718 9602 2770 9614
rect 2718 9538 2770 9550
rect 3278 9602 3330 9614
rect 3278 9538 3330 9550
rect 4510 9602 4562 9614
rect 4510 9538 4562 9550
rect 5854 9602 5906 9614
rect 5854 9538 5906 9550
rect 6414 9602 6466 9614
rect 6414 9538 6466 9550
rect 7086 9602 7138 9614
rect 7086 9538 7138 9550
rect 8318 9602 8370 9614
rect 8318 9538 8370 9550
rect 9438 9602 9490 9614
rect 9438 9538 9490 9550
rect 9774 9602 9826 9614
rect 9774 9538 9826 9550
rect 12910 9602 12962 9614
rect 12910 9538 12962 9550
rect 13806 9602 13858 9614
rect 13806 9538 13858 9550
rect 14030 9602 14082 9614
rect 14030 9538 14082 9550
rect 14590 9602 14642 9614
rect 14590 9538 14642 9550
rect 16270 9602 16322 9614
rect 16270 9538 16322 9550
rect 16718 9602 16770 9614
rect 16718 9538 16770 9550
rect 17390 9602 17442 9614
rect 17390 9538 17442 9550
rect 18286 9602 18338 9614
rect 18286 9538 18338 9550
rect 20190 9602 20242 9614
rect 20190 9538 20242 9550
rect 22990 9602 23042 9614
rect 22990 9538 23042 9550
rect 23214 9602 23266 9614
rect 23214 9538 23266 9550
rect 23774 9602 23826 9614
rect 23774 9538 23826 9550
rect 23998 9602 24050 9614
rect 23998 9538 24050 9550
rect 24446 9602 24498 9614
rect 24446 9538 24498 9550
rect 28142 9602 28194 9614
rect 28142 9538 28194 9550
rect 29710 9602 29762 9614
rect 29710 9538 29762 9550
rect 33294 9602 33346 9614
rect 33294 9538 33346 9550
rect 33854 9602 33906 9614
rect 33854 9538 33906 9550
rect 36766 9602 36818 9614
rect 36766 9538 36818 9550
rect 37438 9602 37490 9614
rect 37438 9538 37490 9550
rect 38670 9602 38722 9614
rect 38670 9538 38722 9550
rect 40014 9602 40066 9614
rect 40014 9538 40066 9550
rect 40574 9602 40626 9614
rect 42142 9602 42194 9614
rect 41682 9550 41694 9602
rect 41746 9550 41758 9602
rect 40574 9538 40626 9550
rect 42142 9538 42194 9550
rect 42702 9602 42754 9614
rect 42702 9538 42754 9550
rect 43262 9602 43314 9614
rect 43262 9538 43314 9550
rect 43934 9602 43986 9614
rect 43934 9538 43986 9550
rect 49198 9602 49250 9614
rect 51214 9602 51266 9614
rect 50306 9550 50318 9602
rect 50370 9550 50382 9602
rect 49198 9538 49250 9550
rect 51214 9538 51266 9550
rect 52110 9602 52162 9614
rect 52110 9538 52162 9550
rect 52558 9602 52610 9614
rect 52558 9538 52610 9550
rect 53790 9602 53842 9614
rect 53790 9538 53842 9550
rect 54350 9602 54402 9614
rect 54350 9538 54402 9550
rect 54798 9602 54850 9614
rect 54798 9538 54850 9550
rect 55246 9602 55298 9614
rect 55246 9538 55298 9550
rect 55918 9602 55970 9614
rect 55918 9538 55970 9550
rect 58046 9602 58098 9614
rect 58046 9538 58098 9550
rect 58494 9602 58546 9614
rect 58494 9538 58546 9550
rect 59054 9602 59106 9614
rect 59054 9538 59106 9550
rect 59502 9602 59554 9614
rect 59502 9538 59554 9550
rect 65102 9602 65154 9614
rect 65102 9538 65154 9550
rect 66110 9602 66162 9614
rect 66110 9538 66162 9550
rect 69470 9602 69522 9614
rect 69470 9538 69522 9550
rect 70366 9602 70418 9614
rect 70366 9538 70418 9550
rect 74622 9602 74674 9614
rect 74622 9538 74674 9550
rect 75518 9602 75570 9614
rect 75518 9538 75570 9550
rect 75854 9602 75906 9614
rect 75854 9538 75906 9550
rect 77534 9602 77586 9614
rect 77534 9538 77586 9550
rect 1344 9434 78784 9468
rect 1344 9382 20534 9434
rect 20586 9382 20638 9434
rect 20690 9382 20742 9434
rect 20794 9382 39854 9434
rect 39906 9382 39958 9434
rect 40010 9382 40062 9434
rect 40114 9382 59174 9434
rect 59226 9382 59278 9434
rect 59330 9382 59382 9434
rect 59434 9382 78494 9434
rect 78546 9382 78598 9434
rect 78650 9382 78702 9434
rect 78754 9382 78784 9434
rect 1344 9348 78784 9382
rect 4734 9266 4786 9278
rect 4734 9202 4786 9214
rect 7870 9266 7922 9278
rect 7870 9202 7922 9214
rect 8094 9266 8146 9278
rect 8094 9202 8146 9214
rect 8654 9266 8706 9278
rect 8654 9202 8706 9214
rect 8878 9266 8930 9278
rect 8878 9202 8930 9214
rect 14702 9266 14754 9278
rect 14702 9202 14754 9214
rect 15150 9266 15202 9278
rect 15150 9202 15202 9214
rect 20078 9266 20130 9278
rect 20078 9202 20130 9214
rect 21646 9266 21698 9278
rect 21646 9202 21698 9214
rect 22654 9266 22706 9278
rect 22654 9202 22706 9214
rect 25006 9266 25058 9278
rect 25006 9202 25058 9214
rect 25902 9266 25954 9278
rect 25902 9202 25954 9214
rect 26126 9266 26178 9278
rect 26126 9202 26178 9214
rect 26238 9266 26290 9278
rect 26238 9202 26290 9214
rect 27022 9266 27074 9278
rect 27022 9202 27074 9214
rect 28814 9266 28866 9278
rect 28814 9202 28866 9214
rect 29486 9266 29538 9278
rect 29486 9202 29538 9214
rect 30830 9266 30882 9278
rect 30830 9202 30882 9214
rect 31390 9266 31442 9278
rect 31390 9202 31442 9214
rect 32734 9266 32786 9278
rect 32734 9202 32786 9214
rect 33854 9266 33906 9278
rect 33854 9202 33906 9214
rect 34302 9266 34354 9278
rect 34302 9202 34354 9214
rect 34974 9266 35026 9278
rect 34974 9202 35026 9214
rect 35758 9266 35810 9278
rect 35758 9202 35810 9214
rect 36542 9266 36594 9278
rect 36542 9202 36594 9214
rect 37886 9266 37938 9278
rect 37886 9202 37938 9214
rect 39566 9266 39618 9278
rect 39566 9202 39618 9214
rect 40686 9266 40738 9278
rect 40686 9202 40738 9214
rect 42142 9266 42194 9278
rect 42142 9202 42194 9214
rect 43038 9266 43090 9278
rect 43038 9202 43090 9214
rect 43598 9266 43650 9278
rect 43598 9202 43650 9214
rect 44046 9266 44098 9278
rect 44046 9202 44098 9214
rect 49982 9266 50034 9278
rect 49982 9202 50034 9214
rect 62750 9266 62802 9278
rect 62750 9202 62802 9214
rect 62862 9266 62914 9278
rect 62862 9202 62914 9214
rect 63534 9266 63586 9278
rect 63534 9202 63586 9214
rect 67230 9266 67282 9278
rect 67230 9202 67282 9214
rect 69022 9266 69074 9278
rect 69022 9202 69074 9214
rect 69582 9266 69634 9278
rect 69582 9202 69634 9214
rect 70030 9266 70082 9278
rect 70030 9202 70082 9214
rect 70926 9266 70978 9278
rect 70926 9202 70978 9214
rect 71710 9266 71762 9278
rect 71710 9202 71762 9214
rect 72270 9266 72322 9278
rect 72270 9202 72322 9214
rect 73502 9266 73554 9278
rect 73502 9202 73554 9214
rect 73614 9266 73666 9278
rect 73614 9202 73666 9214
rect 77086 9266 77138 9278
rect 77086 9202 77138 9214
rect 77422 9266 77474 9278
rect 77422 9202 77474 9214
rect 5742 9154 5794 9166
rect 5742 9090 5794 9102
rect 8990 9154 9042 9166
rect 8990 9090 9042 9102
rect 11342 9154 11394 9166
rect 11342 9090 11394 9102
rect 12014 9154 12066 9166
rect 12014 9090 12066 9102
rect 19294 9154 19346 9166
rect 19294 9090 19346 9102
rect 24334 9154 24386 9166
rect 24334 9090 24386 9102
rect 26350 9154 26402 9166
rect 26350 9090 26402 9102
rect 30606 9154 30658 9166
rect 30606 9090 30658 9102
rect 32846 9154 32898 9166
rect 32846 9090 32898 9102
rect 34862 9154 34914 9166
rect 34862 9090 34914 9102
rect 36430 9154 36482 9166
rect 36430 9090 36482 9102
rect 37326 9154 37378 9166
rect 37326 9090 37378 9102
rect 40014 9154 40066 9166
rect 40014 9090 40066 9102
rect 40574 9154 40626 9166
rect 40574 9090 40626 9102
rect 48750 9154 48802 9166
rect 48750 9090 48802 9102
rect 49422 9154 49474 9166
rect 54350 9154 54402 9166
rect 50866 9102 50878 9154
rect 50930 9102 50942 9154
rect 49422 9090 49474 9102
rect 54350 9090 54402 9102
rect 56142 9154 56194 9166
rect 56142 9090 56194 9102
rect 66782 9154 66834 9166
rect 66782 9090 66834 9102
rect 67454 9154 67506 9166
rect 67454 9090 67506 9102
rect 67566 9154 67618 9166
rect 67566 9090 67618 9102
rect 68238 9154 68290 9166
rect 68238 9090 68290 9102
rect 73390 9154 73442 9166
rect 73390 9090 73442 9102
rect 76862 9154 76914 9166
rect 76862 9090 76914 9102
rect 4286 9042 4338 9054
rect 4958 9042 5010 9054
rect 2818 8990 2830 9042
rect 2882 8990 2894 9042
rect 4610 8990 4622 9042
rect 4674 8990 4686 9042
rect 4286 8978 4338 8990
rect 4958 8978 5010 8990
rect 5518 9042 5570 9054
rect 5518 8978 5570 8990
rect 5854 9042 5906 9054
rect 7198 9042 7250 9054
rect 6738 8990 6750 9042
rect 6802 8990 6814 9042
rect 5854 8978 5906 8990
rect 7198 8978 7250 8990
rect 8206 9042 8258 9054
rect 11902 9042 11954 9054
rect 10882 8990 10894 9042
rect 10946 8990 10958 9042
rect 8206 8978 8258 8990
rect 11902 8978 11954 8990
rect 13246 9042 13298 9054
rect 13246 8978 13298 8990
rect 18062 9042 18114 9054
rect 18062 8978 18114 8990
rect 18622 9042 18674 9054
rect 18622 8978 18674 8990
rect 19182 9042 19234 9054
rect 19182 8978 19234 8990
rect 19518 9042 19570 9054
rect 19518 8978 19570 8990
rect 22094 9042 22146 9054
rect 28142 9042 28194 9054
rect 23538 8990 23550 9042
rect 23602 8990 23614 9042
rect 22094 8978 22146 8990
rect 28142 8978 28194 8990
rect 28702 9042 28754 9054
rect 28702 8978 28754 8990
rect 30494 9042 30546 9054
rect 30494 8978 30546 8990
rect 31502 9042 31554 9054
rect 31502 8978 31554 8990
rect 31614 9042 31666 9054
rect 32062 9042 32114 9054
rect 31714 8990 31726 9042
rect 31778 8990 31790 9042
rect 31614 8978 31666 8990
rect 32062 8978 32114 8990
rect 32510 9042 32562 9054
rect 32510 8978 32562 8990
rect 35198 9042 35250 9054
rect 35198 8978 35250 8990
rect 35646 9042 35698 9054
rect 35646 8978 35698 8990
rect 35982 9042 36034 9054
rect 35982 8978 36034 8990
rect 37214 9042 37266 9054
rect 37214 8978 37266 8990
rect 37550 9042 37602 9054
rect 37550 8978 37602 8990
rect 40910 9042 40962 9054
rect 40910 8978 40962 8990
rect 41582 9042 41634 9054
rect 41582 8978 41634 8990
rect 41806 9042 41858 9054
rect 41806 8978 41858 8990
rect 42030 9042 42082 9054
rect 42030 8978 42082 8990
rect 42254 9042 42306 9054
rect 42254 8978 42306 8990
rect 42926 9042 42978 9054
rect 42926 8978 42978 8990
rect 43262 9042 43314 9054
rect 55918 9042 55970 9054
rect 51202 8990 51214 9042
rect 51266 8990 51278 9042
rect 52098 8990 52110 9042
rect 52162 8990 52174 9042
rect 54786 8990 54798 9042
rect 54850 8990 54862 9042
rect 43262 8978 43314 8990
rect 55918 8978 55970 8990
rect 56590 9042 56642 9054
rect 56590 8978 56642 8990
rect 57486 9042 57538 9054
rect 57486 8978 57538 8990
rect 58046 9042 58098 9054
rect 58046 8978 58098 8990
rect 58494 9042 58546 9054
rect 60846 9042 60898 9054
rect 62302 9042 62354 9054
rect 60162 8990 60174 9042
rect 60226 8990 60238 9042
rect 61506 8990 61518 9042
rect 61570 8990 61582 9042
rect 58494 8978 58546 8990
rect 60846 8978 60898 8990
rect 62302 8978 62354 8990
rect 62974 9042 63026 9054
rect 62974 8978 63026 8990
rect 64094 9042 64146 9054
rect 64094 8978 64146 8990
rect 65438 9042 65490 9054
rect 65438 8978 65490 8990
rect 68350 9042 68402 9054
rect 68350 8978 68402 8990
rect 69134 9042 69186 9054
rect 69134 8978 69186 8990
rect 71598 9042 71650 9054
rect 71598 8978 71650 8990
rect 71934 9042 71986 9054
rect 76750 9042 76802 9054
rect 73938 8990 73950 9042
rect 74002 8990 74014 9042
rect 75954 8990 75966 9042
rect 76018 8990 76030 9042
rect 71934 8978 71986 8990
rect 76750 8978 76802 8990
rect 3726 8930 3778 8942
rect 1922 8878 1934 8930
rect 1986 8878 1998 8930
rect 3726 8866 3778 8878
rect 4846 8930 4898 8942
rect 4846 8866 4898 8878
rect 9662 8930 9714 8942
rect 15486 8930 15538 8942
rect 10434 8878 10446 8930
rect 10498 8878 10510 8930
rect 9662 8866 9714 8878
rect 15486 8866 15538 8878
rect 20526 8930 20578 8942
rect 20526 8866 20578 8878
rect 20974 8930 21026 8942
rect 29934 8930 29986 8942
rect 23762 8878 23774 8930
rect 23826 8878 23838 8930
rect 27682 8878 27694 8930
rect 27746 8878 27758 8930
rect 20974 8866 21026 8878
rect 29934 8866 29986 8878
rect 38334 8930 38386 8942
rect 38334 8866 38386 8878
rect 52782 8930 52834 8942
rect 52782 8866 52834 8878
rect 53566 8930 53618 8942
rect 56030 8930 56082 8942
rect 54674 8878 54686 8930
rect 54738 8878 54750 8930
rect 53566 8866 53618 8878
rect 56030 8866 56082 8878
rect 62526 8930 62578 8942
rect 62526 8866 62578 8878
rect 64542 8930 64594 8942
rect 64542 8866 64594 8878
rect 65774 8930 65826 8942
rect 65774 8866 65826 8878
rect 66334 8930 66386 8942
rect 66334 8866 66386 8878
rect 70478 8930 70530 8942
rect 70478 8866 70530 8878
rect 74510 8930 74562 8942
rect 77870 8930 77922 8942
rect 75506 8878 75518 8930
rect 75570 8878 75582 8930
rect 74510 8866 74562 8878
rect 77870 8866 77922 8878
rect 12014 8818 12066 8830
rect 12014 8754 12066 8766
rect 13470 8818 13522 8830
rect 28814 8818 28866 8830
rect 13794 8766 13806 8818
rect 13858 8766 13870 8818
rect 13470 8754 13522 8766
rect 28814 8754 28866 8766
rect 36542 8818 36594 8830
rect 68238 8818 68290 8830
rect 59714 8766 59726 8818
rect 59778 8766 59790 8818
rect 36542 8754 36594 8766
rect 68238 8754 68290 8766
rect 69022 8818 69074 8830
rect 69022 8754 69074 8766
rect 1344 8650 78624 8684
rect 1344 8598 10874 8650
rect 10926 8598 10978 8650
rect 11030 8598 11082 8650
rect 11134 8598 30194 8650
rect 30246 8598 30298 8650
rect 30350 8598 30402 8650
rect 30454 8598 49514 8650
rect 49566 8598 49618 8650
rect 49670 8598 49722 8650
rect 49774 8598 68834 8650
rect 68886 8598 68938 8650
rect 68990 8598 69042 8650
rect 69094 8598 78624 8650
rect 1344 8564 78624 8598
rect 36430 8482 36482 8494
rect 36430 8418 36482 8430
rect 51102 8482 51154 8494
rect 56590 8482 56642 8494
rect 54898 8430 54910 8482
rect 54962 8430 54974 8482
rect 51102 8418 51154 8430
rect 56590 8418 56642 8430
rect 57374 8482 57426 8494
rect 57374 8418 57426 8430
rect 2158 8370 2210 8382
rect 2158 8306 2210 8318
rect 7198 8370 7250 8382
rect 13918 8370 13970 8382
rect 7746 8318 7758 8370
rect 7810 8318 7822 8370
rect 7198 8306 7250 8318
rect 13918 8306 13970 8318
rect 20078 8370 20130 8382
rect 24222 8370 24274 8382
rect 30158 8370 30210 8382
rect 23426 8318 23438 8370
rect 23490 8318 23502 8370
rect 28578 8318 28590 8370
rect 28642 8318 28654 8370
rect 20078 8306 20130 8318
rect 24222 8306 24274 8318
rect 30158 8306 30210 8318
rect 34862 8370 34914 8382
rect 34862 8306 34914 8318
rect 35310 8370 35362 8382
rect 35310 8306 35362 8318
rect 35758 8370 35810 8382
rect 35758 8306 35810 8318
rect 38110 8370 38162 8382
rect 38110 8306 38162 8318
rect 41470 8370 41522 8382
rect 41470 8306 41522 8318
rect 45838 8370 45890 8382
rect 45838 8306 45890 8318
rect 47518 8370 47570 8382
rect 47518 8306 47570 8318
rect 50542 8370 50594 8382
rect 60398 8370 60450 8382
rect 63086 8370 63138 8382
rect 55570 8318 55582 8370
rect 55634 8318 55646 8370
rect 61618 8318 61630 8370
rect 61682 8318 61694 8370
rect 50542 8306 50594 8318
rect 60398 8306 60450 8318
rect 63086 8306 63138 8318
rect 65774 8370 65826 8382
rect 69246 8370 69298 8382
rect 67554 8318 67566 8370
rect 67618 8318 67630 8370
rect 65774 8306 65826 8318
rect 69246 8306 69298 8318
rect 70478 8370 70530 8382
rect 70478 8306 70530 8318
rect 75406 8370 75458 8382
rect 77858 8318 77870 8370
rect 77922 8318 77934 8370
rect 75406 8306 75458 8318
rect 3054 8258 3106 8270
rect 3054 8194 3106 8206
rect 3390 8258 3442 8270
rect 4846 8258 4898 8270
rect 9326 8258 9378 8270
rect 4274 8206 4286 8258
rect 4338 8206 4350 8258
rect 4610 8206 4622 8258
rect 4674 8206 4686 8258
rect 8866 8206 8878 8258
rect 8930 8206 8942 8258
rect 3390 8194 3442 8206
rect 4846 8194 4898 8206
rect 9326 8194 9378 8206
rect 9774 8258 9826 8270
rect 16606 8258 16658 8270
rect 15250 8206 15262 8258
rect 15314 8206 15326 8258
rect 9774 8194 9826 8206
rect 16606 8194 16658 8206
rect 17166 8258 17218 8270
rect 17166 8194 17218 8206
rect 17502 8258 17554 8270
rect 18846 8258 18898 8270
rect 18274 8206 18286 8258
rect 18338 8206 18350 8258
rect 17502 8194 17554 8206
rect 18846 8194 18898 8206
rect 19518 8258 19570 8270
rect 19518 8194 19570 8206
rect 22654 8258 22706 8270
rect 26910 8258 26962 8270
rect 28814 8258 28866 8270
rect 23538 8206 23550 8258
rect 23602 8206 23614 8258
rect 28354 8206 28366 8258
rect 28418 8206 28430 8258
rect 22654 8194 22706 8206
rect 26910 8194 26962 8206
rect 28814 8194 28866 8206
rect 31390 8258 31442 8270
rect 33182 8258 33234 8270
rect 31826 8206 31838 8258
rect 31890 8206 31902 8258
rect 31390 8194 31442 8206
rect 33182 8194 33234 8206
rect 36206 8258 36258 8270
rect 37550 8258 37602 8270
rect 36754 8206 36766 8258
rect 36818 8206 36830 8258
rect 36206 8194 36258 8206
rect 37550 8194 37602 8206
rect 37774 8258 37826 8270
rect 37774 8194 37826 8206
rect 43486 8258 43538 8270
rect 46734 8258 46786 8270
rect 46274 8206 46286 8258
rect 46338 8206 46350 8258
rect 43486 8194 43538 8206
rect 46734 8194 46786 8206
rect 47406 8258 47458 8270
rect 47406 8194 47458 8206
rect 48078 8258 48130 8270
rect 56702 8258 56754 8270
rect 50754 8206 50766 8258
rect 50818 8206 50830 8258
rect 55458 8206 55470 8258
rect 55522 8206 55534 8258
rect 48078 8194 48130 8206
rect 56702 8194 56754 8206
rect 57486 8258 57538 8270
rect 57486 8194 57538 8206
rect 58382 8258 58434 8270
rect 60286 8258 60338 8270
rect 64990 8258 65042 8270
rect 59602 8206 59614 8258
rect 59666 8206 59678 8258
rect 62066 8206 62078 8258
rect 62130 8206 62142 8258
rect 63298 8206 63310 8258
rect 63362 8206 63374 8258
rect 63522 8206 63534 8258
rect 63586 8206 63598 8258
rect 58382 8194 58434 8206
rect 60286 8194 60338 8206
rect 64990 8194 65042 8206
rect 66670 8258 66722 8270
rect 66670 8194 66722 8206
rect 71150 8258 71202 8270
rect 72046 8258 72098 8270
rect 71362 8206 71374 8258
rect 71426 8206 71438 8258
rect 71150 8194 71202 8206
rect 72046 8194 72098 8206
rect 72718 8258 72770 8270
rect 73614 8258 73666 8270
rect 73154 8206 73166 8258
rect 73218 8206 73230 8258
rect 72718 8194 72770 8206
rect 73614 8194 73666 8206
rect 74622 8258 74674 8270
rect 74622 8194 74674 8206
rect 74958 8258 75010 8270
rect 74958 8194 75010 8206
rect 75518 8258 75570 8270
rect 77310 8258 77362 8270
rect 75954 8206 75966 8258
rect 76018 8206 76030 8258
rect 75518 8194 75570 8206
rect 77310 8194 77362 8206
rect 77534 8258 77586 8270
rect 77534 8194 77586 8206
rect 5854 8146 5906 8158
rect 5854 8082 5906 8094
rect 10110 8146 10162 8158
rect 19070 8146 19122 8158
rect 14242 8094 14254 8146
rect 14306 8094 14318 8146
rect 10110 8082 10162 8094
rect 19070 8082 19122 8094
rect 20190 8146 20242 8158
rect 20190 8082 20242 8094
rect 26350 8146 26402 8158
rect 26350 8082 26402 8094
rect 27022 8146 27074 8158
rect 27022 8082 27074 8094
rect 27246 8146 27298 8158
rect 27246 8082 27298 8094
rect 32286 8146 32338 8158
rect 32286 8082 32338 8094
rect 38222 8146 38274 8158
rect 47630 8146 47682 8158
rect 41570 8094 41582 8146
rect 41634 8094 41646 8146
rect 43250 8094 43262 8146
rect 43314 8094 43326 8146
rect 38222 8082 38274 8094
rect 47630 8082 47682 8094
rect 48526 8146 48578 8158
rect 48526 8082 48578 8094
rect 51886 8146 51938 8158
rect 51886 8082 51938 8094
rect 62526 8146 62578 8158
rect 62526 8082 62578 8094
rect 65326 8146 65378 8158
rect 65326 8082 65378 8094
rect 66782 8146 66834 8158
rect 66782 8082 66834 8094
rect 69806 8146 69858 8158
rect 69806 8082 69858 8094
rect 70366 8146 70418 8158
rect 70366 8082 70418 8094
rect 2494 8034 2546 8046
rect 2494 7970 2546 7982
rect 3166 8034 3218 8046
rect 3166 7970 3218 7982
rect 6190 8034 6242 8046
rect 6190 7970 6242 7982
rect 6638 8034 6690 8046
rect 6638 7970 6690 7982
rect 8206 8034 8258 8046
rect 8206 7970 8258 7982
rect 9998 8034 10050 8046
rect 9998 7970 10050 7982
rect 10670 8034 10722 8046
rect 10670 7970 10722 7982
rect 11006 8034 11058 8046
rect 17278 8034 17330 8046
rect 15810 7982 15822 8034
rect 15874 7982 15886 8034
rect 11006 7970 11058 7982
rect 17278 7970 17330 7982
rect 19966 8034 20018 8046
rect 19966 7970 20018 7982
rect 21646 8034 21698 8046
rect 21646 7970 21698 7982
rect 22206 8034 22258 8046
rect 22206 7970 22258 7982
rect 22430 8034 22482 8046
rect 22430 7970 22482 7982
rect 22542 8034 22594 8046
rect 22542 7970 22594 7982
rect 24670 8034 24722 8046
rect 24670 7970 24722 7982
rect 25118 8034 25170 8046
rect 25118 7970 25170 7982
rect 29486 8034 29538 8046
rect 29486 7970 29538 7982
rect 30718 8034 30770 8046
rect 30718 7970 30770 7982
rect 37998 8034 38050 8046
rect 37998 7970 38050 7982
rect 40686 8034 40738 8046
rect 40686 7970 40738 7982
rect 48638 8034 48690 8046
rect 48638 7970 48690 7982
rect 48862 8034 48914 8046
rect 48862 7970 48914 7982
rect 49198 8034 49250 8046
rect 49198 7970 49250 7982
rect 49646 8034 49698 8046
rect 49646 7970 49698 7982
rect 50430 8034 50482 8046
rect 50430 7970 50482 7982
rect 50654 8034 50706 8046
rect 50654 7970 50706 7982
rect 51550 8034 51602 8046
rect 51550 7970 51602 7982
rect 51774 8034 51826 8046
rect 51774 7970 51826 7982
rect 52334 8034 52386 8046
rect 52334 7970 52386 7982
rect 53342 8034 53394 8046
rect 53342 7970 53394 7982
rect 53790 8034 53842 8046
rect 53790 7970 53842 7982
rect 54238 8034 54290 8046
rect 54238 7970 54290 7982
rect 56590 8034 56642 8046
rect 56590 7970 56642 7982
rect 57374 8034 57426 8046
rect 57374 7970 57426 7982
rect 57934 8034 57986 8046
rect 57934 7970 57986 7982
rect 58830 8034 58882 8046
rect 58830 7970 58882 7982
rect 64654 8034 64706 8046
rect 64654 7970 64706 7982
rect 65214 8034 65266 8046
rect 65214 7970 65266 7982
rect 67006 8034 67058 8046
rect 67006 7970 67058 7982
rect 68014 8034 68066 8046
rect 68014 7970 68066 7982
rect 68462 8034 68514 8046
rect 68462 7970 68514 7982
rect 74174 8034 74226 8046
rect 74174 7970 74226 7982
rect 74734 8034 74786 8046
rect 74734 7970 74786 7982
rect 1344 7866 78784 7900
rect 1344 7814 20534 7866
rect 20586 7814 20638 7866
rect 20690 7814 20742 7866
rect 20794 7814 39854 7866
rect 39906 7814 39958 7866
rect 40010 7814 40062 7866
rect 40114 7814 59174 7866
rect 59226 7814 59278 7866
rect 59330 7814 59382 7866
rect 59434 7814 78494 7866
rect 78546 7814 78598 7866
rect 78650 7814 78702 7866
rect 78754 7814 78784 7866
rect 1344 7780 78784 7814
rect 1822 7698 1874 7710
rect 1822 7634 1874 7646
rect 2270 7698 2322 7710
rect 2270 7634 2322 7646
rect 5518 7698 5570 7710
rect 5518 7634 5570 7646
rect 6302 7698 6354 7710
rect 6302 7634 6354 7646
rect 9886 7698 9938 7710
rect 9886 7634 9938 7646
rect 10446 7698 10498 7710
rect 10446 7634 10498 7646
rect 10894 7698 10946 7710
rect 10894 7634 10946 7646
rect 12798 7698 12850 7710
rect 12798 7634 12850 7646
rect 13582 7698 13634 7710
rect 13582 7634 13634 7646
rect 13694 7698 13746 7710
rect 13694 7634 13746 7646
rect 14590 7698 14642 7710
rect 14590 7634 14642 7646
rect 14814 7698 14866 7710
rect 14814 7634 14866 7646
rect 15374 7698 15426 7710
rect 15374 7634 15426 7646
rect 15822 7698 15874 7710
rect 15822 7634 15874 7646
rect 17614 7698 17666 7710
rect 17614 7634 17666 7646
rect 23662 7698 23714 7710
rect 23662 7634 23714 7646
rect 26686 7698 26738 7710
rect 26686 7634 26738 7646
rect 27134 7698 27186 7710
rect 27134 7634 27186 7646
rect 28702 7698 28754 7710
rect 28702 7634 28754 7646
rect 28926 7698 28978 7710
rect 28926 7634 28978 7646
rect 29598 7698 29650 7710
rect 29598 7634 29650 7646
rect 29934 7698 29986 7710
rect 29934 7634 29986 7646
rect 32734 7698 32786 7710
rect 32734 7634 32786 7646
rect 40014 7698 40066 7710
rect 40014 7634 40066 7646
rect 44382 7698 44434 7710
rect 44382 7634 44434 7646
rect 48078 7698 48130 7710
rect 48078 7634 48130 7646
rect 53566 7698 53618 7710
rect 53566 7634 53618 7646
rect 59166 7698 59218 7710
rect 59166 7634 59218 7646
rect 61070 7698 61122 7710
rect 61070 7634 61122 7646
rect 63086 7698 63138 7710
rect 63086 7634 63138 7646
rect 65550 7698 65602 7710
rect 65550 7634 65602 7646
rect 65774 7698 65826 7710
rect 65774 7634 65826 7646
rect 66558 7698 66610 7710
rect 66558 7634 66610 7646
rect 67454 7698 67506 7710
rect 67454 7634 67506 7646
rect 68462 7698 68514 7710
rect 68462 7634 68514 7646
rect 69806 7698 69858 7710
rect 69806 7634 69858 7646
rect 69918 7698 69970 7710
rect 69918 7634 69970 7646
rect 73278 7698 73330 7710
rect 73278 7634 73330 7646
rect 75518 7698 75570 7710
rect 75518 7634 75570 7646
rect 2718 7586 2770 7598
rect 2718 7522 2770 7534
rect 3054 7586 3106 7598
rect 3054 7522 3106 7534
rect 6414 7586 6466 7598
rect 6414 7522 6466 7534
rect 7870 7586 7922 7598
rect 7870 7522 7922 7534
rect 9774 7586 9826 7598
rect 9774 7522 9826 7534
rect 19182 7586 19234 7598
rect 19182 7522 19234 7534
rect 23886 7586 23938 7598
rect 23886 7522 23938 7534
rect 29038 7586 29090 7598
rect 29038 7522 29090 7534
rect 31614 7586 31666 7598
rect 48302 7586 48354 7598
rect 36530 7534 36542 7586
rect 36594 7534 36606 7586
rect 31614 7522 31666 7534
rect 48302 7522 48354 7534
rect 52446 7586 52498 7598
rect 52446 7522 52498 7534
rect 56702 7586 56754 7598
rect 56702 7522 56754 7534
rect 63310 7586 63362 7598
rect 63310 7522 63362 7534
rect 68126 7586 68178 7598
rect 68126 7522 68178 7534
rect 70590 7586 70642 7598
rect 70590 7522 70642 7534
rect 75294 7586 75346 7598
rect 75294 7522 75346 7534
rect 76974 7586 77026 7598
rect 76974 7522 77026 7534
rect 77534 7586 77586 7598
rect 77534 7522 77586 7534
rect 77870 7586 77922 7598
rect 77870 7522 77922 7534
rect 4510 7474 4562 7486
rect 4162 7422 4174 7474
rect 4226 7422 4238 7474
rect 4510 7410 4562 7422
rect 5070 7474 5122 7486
rect 5070 7410 5122 7422
rect 5630 7474 5682 7486
rect 5630 7410 5682 7422
rect 5742 7474 5794 7486
rect 13470 7474 13522 7486
rect 14142 7474 14194 7486
rect 8418 7422 8430 7474
rect 8482 7422 8494 7474
rect 13794 7422 13806 7474
rect 13858 7422 13870 7474
rect 5742 7410 5794 7422
rect 13470 7410 13522 7422
rect 14142 7410 14194 7422
rect 14926 7474 14978 7486
rect 19070 7474 19122 7486
rect 23998 7474 24050 7486
rect 18498 7422 18510 7474
rect 18562 7422 18574 7474
rect 22754 7422 22766 7474
rect 22818 7422 22830 7474
rect 14926 7410 14978 7422
rect 19070 7410 19122 7422
rect 23998 7410 24050 7422
rect 28030 7474 28082 7486
rect 28030 7410 28082 7422
rect 31502 7474 31554 7486
rect 31502 7410 31554 7422
rect 31838 7474 31890 7486
rect 31838 7410 31890 7422
rect 32174 7474 32226 7486
rect 32174 7410 32226 7422
rect 32622 7474 32674 7486
rect 32622 7410 32674 7422
rect 32846 7474 32898 7486
rect 39902 7474 39954 7486
rect 37762 7422 37774 7474
rect 37826 7422 37838 7474
rect 32846 7410 32898 7422
rect 39902 7410 39954 7422
rect 40126 7474 40178 7486
rect 40126 7410 40178 7422
rect 40574 7474 40626 7486
rect 40574 7410 40626 7422
rect 44270 7474 44322 7486
rect 44270 7410 44322 7422
rect 44494 7474 44546 7486
rect 44494 7410 44546 7422
rect 44942 7474 44994 7486
rect 48414 7474 48466 7486
rect 52670 7474 52722 7486
rect 47394 7422 47406 7474
rect 47458 7422 47470 7474
rect 49858 7422 49870 7474
rect 49922 7422 49934 7474
rect 51090 7422 51102 7474
rect 51154 7422 51166 7474
rect 44942 7410 44994 7422
rect 48414 7410 48466 7422
rect 52670 7410 52722 7422
rect 52894 7474 52946 7486
rect 52894 7410 52946 7422
rect 53006 7474 53058 7486
rect 62638 7474 62690 7486
rect 54562 7422 54574 7474
rect 54626 7422 54638 7474
rect 56130 7422 56142 7474
rect 56194 7422 56206 7474
rect 53006 7410 53058 7422
rect 62638 7410 62690 7422
rect 65438 7474 65490 7486
rect 65438 7410 65490 7422
rect 66110 7474 66162 7486
rect 66110 7410 66162 7422
rect 67342 7474 67394 7486
rect 67342 7410 67394 7422
rect 67678 7474 67730 7486
rect 67678 7410 67730 7422
rect 69358 7474 69410 7486
rect 69358 7410 69410 7422
rect 70030 7474 70082 7486
rect 75182 7474 75234 7486
rect 76862 7474 76914 7486
rect 71698 7422 71710 7474
rect 71762 7422 71774 7474
rect 76290 7422 76302 7474
rect 76354 7422 76366 7474
rect 70030 7410 70082 7422
rect 75182 7410 75234 7422
rect 76862 7410 76914 7422
rect 4622 7362 4674 7374
rect 16270 7362 16322 7374
rect 8642 7310 8654 7362
rect 8706 7310 8718 7362
rect 4622 7298 4674 7310
rect 16270 7298 16322 7310
rect 16830 7362 16882 7374
rect 24782 7362 24834 7374
rect 22306 7310 22318 7362
rect 22370 7310 22382 7362
rect 16830 7298 16882 7310
rect 24782 7298 24834 7310
rect 25566 7362 25618 7374
rect 25566 7298 25618 7310
rect 26014 7362 26066 7374
rect 26014 7298 26066 7310
rect 28254 7362 28306 7374
rect 28254 7298 28306 7310
rect 30942 7362 30994 7374
rect 38446 7362 38498 7374
rect 36306 7310 36318 7362
rect 36370 7310 36382 7362
rect 30942 7298 30994 7310
rect 38446 7298 38498 7310
rect 39342 7362 39394 7374
rect 39342 7298 39394 7310
rect 45390 7362 45442 7374
rect 45390 7298 45442 7310
rect 46622 7362 46674 7374
rect 52782 7362 52834 7374
rect 57374 7362 57426 7374
rect 47282 7310 47294 7362
rect 47346 7310 47358 7362
rect 50082 7310 50094 7362
rect 50146 7310 50158 7362
rect 54674 7310 54686 7362
rect 54738 7310 54750 7362
rect 46622 7298 46674 7310
rect 52782 7298 52834 7310
rect 57374 7298 57426 7310
rect 57822 7362 57874 7374
rect 57822 7298 57874 7310
rect 58382 7362 58434 7374
rect 58382 7298 58434 7310
rect 58718 7362 58770 7374
rect 58718 7298 58770 7310
rect 59726 7362 59778 7374
rect 59726 7298 59778 7310
rect 60062 7362 60114 7374
rect 60062 7298 60114 7310
rect 60510 7362 60562 7374
rect 60510 7298 60562 7310
rect 61406 7362 61458 7374
rect 61406 7298 61458 7310
rect 61854 7362 61906 7374
rect 61854 7298 61906 7310
rect 63198 7362 63250 7374
rect 63198 7298 63250 7310
rect 63870 7362 63922 7374
rect 63870 7298 63922 7310
rect 64318 7362 64370 7374
rect 64318 7298 64370 7310
rect 64654 7362 64706 7374
rect 64654 7298 64706 7310
rect 69582 7362 69634 7374
rect 73838 7362 73890 7374
rect 71810 7310 71822 7362
rect 71874 7310 71886 7362
rect 69582 7298 69634 7310
rect 73838 7298 73890 7310
rect 74174 7362 74226 7374
rect 74174 7298 74226 7310
rect 74734 7362 74786 7374
rect 74734 7298 74786 7310
rect 9886 7250 9938 7262
rect 22642 7198 22654 7250
rect 22706 7198 22718 7250
rect 27682 7198 27694 7250
rect 27746 7198 27758 7250
rect 51314 7198 51326 7250
rect 51378 7198 51390 7250
rect 57922 7198 57934 7250
rect 57986 7247 57998 7250
rect 58706 7247 58718 7250
rect 57986 7201 58718 7247
rect 57986 7198 57998 7201
rect 58706 7198 58718 7201
rect 58770 7198 58782 7250
rect 60498 7198 60510 7250
rect 60562 7247 60574 7250
rect 61842 7247 61854 7250
rect 60562 7201 61854 7247
rect 60562 7198 60574 7201
rect 61842 7198 61854 7201
rect 61906 7198 61918 7250
rect 63970 7198 63982 7250
rect 64034 7247 64046 7250
rect 64642 7247 64654 7250
rect 64034 7201 64654 7247
rect 64034 7198 64046 7201
rect 64642 7198 64654 7201
rect 64706 7198 64718 7250
rect 68002 7198 68014 7250
rect 68066 7247 68078 7250
rect 68450 7247 68462 7250
rect 68066 7201 68462 7247
rect 68066 7198 68078 7201
rect 68450 7198 68462 7201
rect 68514 7198 68526 7250
rect 72258 7198 72270 7250
rect 72322 7198 72334 7250
rect 73826 7198 73838 7250
rect 73890 7247 73902 7250
rect 74162 7247 74174 7250
rect 73890 7201 74174 7247
rect 73890 7198 73902 7201
rect 74162 7198 74174 7201
rect 74226 7198 74238 7250
rect 9886 7186 9938 7198
rect 1344 7082 78624 7116
rect 1344 7030 10874 7082
rect 10926 7030 10978 7082
rect 11030 7030 11082 7082
rect 11134 7030 30194 7082
rect 30246 7030 30298 7082
rect 30350 7030 30402 7082
rect 30454 7030 49514 7082
rect 49566 7030 49618 7082
rect 49670 7030 49722 7082
rect 49774 7030 68834 7082
rect 68886 7030 68938 7082
rect 68990 7030 69042 7082
rect 69094 7030 78624 7082
rect 1344 6996 78624 7030
rect 35534 6914 35586 6926
rect 50094 6914 50146 6926
rect 18946 6862 18958 6914
rect 19010 6862 19022 6914
rect 32498 6862 32510 6914
rect 32562 6862 32574 6914
rect 39890 6862 39902 6914
rect 39954 6862 39966 6914
rect 35534 6850 35586 6862
rect 50094 6850 50146 6862
rect 50878 6914 50930 6926
rect 50878 6850 50930 6862
rect 54686 6914 54738 6926
rect 54686 6850 54738 6862
rect 55358 6914 55410 6926
rect 66434 6862 66446 6914
rect 66498 6862 66510 6914
rect 55358 6850 55410 6862
rect 8430 6802 8482 6814
rect 8430 6738 8482 6750
rect 13694 6802 13746 6814
rect 13694 6738 13746 6750
rect 15038 6802 15090 6814
rect 27806 6802 27858 6814
rect 22194 6750 22206 6802
rect 22258 6750 22270 6802
rect 15038 6738 15090 6750
rect 27806 6738 27858 6750
rect 29486 6802 29538 6814
rect 49534 6802 49586 6814
rect 32050 6750 32062 6802
rect 32114 6750 32126 6802
rect 43474 6750 43486 6802
rect 43538 6750 43550 6802
rect 29486 6738 29538 6750
rect 49534 6738 49586 6750
rect 55918 6802 55970 6814
rect 55918 6738 55970 6750
rect 60622 6802 60674 6814
rect 62178 6750 62190 6802
rect 62242 6750 62254 6802
rect 65762 6750 65774 6802
rect 65826 6750 65838 6802
rect 60622 6738 60674 6750
rect 4734 6690 4786 6702
rect 3042 6638 3054 6690
rect 3106 6638 3118 6690
rect 4734 6626 4786 6638
rect 9326 6690 9378 6702
rect 9326 6626 9378 6638
rect 9662 6690 9714 6702
rect 9662 6626 9714 6638
rect 10446 6690 10498 6702
rect 10446 6626 10498 6638
rect 10894 6690 10946 6702
rect 10894 6626 10946 6638
rect 12574 6690 12626 6702
rect 12574 6626 12626 6638
rect 12910 6690 12962 6702
rect 12910 6626 12962 6638
rect 13918 6690 13970 6702
rect 13918 6626 13970 6638
rect 14142 6690 14194 6702
rect 14142 6626 14194 6638
rect 15598 6690 15650 6702
rect 15598 6626 15650 6638
rect 16606 6690 16658 6702
rect 18062 6690 18114 6702
rect 19966 6690 20018 6702
rect 22654 6690 22706 6702
rect 17714 6638 17726 6690
rect 17778 6638 17790 6690
rect 19058 6638 19070 6690
rect 19122 6638 19134 6690
rect 21970 6638 21982 6690
rect 22034 6638 22046 6690
rect 16606 6626 16658 6638
rect 18062 6626 18114 6638
rect 19966 6626 20018 6638
rect 22654 6626 22706 6638
rect 23998 6690 24050 6702
rect 26350 6690 26402 6702
rect 24322 6638 24334 6690
rect 24386 6638 24398 6690
rect 23998 6626 24050 6638
rect 26350 6626 26402 6638
rect 27134 6690 27186 6702
rect 27134 6626 27186 6638
rect 27582 6690 27634 6702
rect 27582 6626 27634 6638
rect 28254 6690 28306 6702
rect 28254 6626 28306 6638
rect 31166 6690 31218 6702
rect 34974 6690 35026 6702
rect 32386 6638 32398 6690
rect 32450 6638 32462 6690
rect 31166 6626 31218 6638
rect 34974 6626 35026 6638
rect 35310 6690 35362 6702
rect 35310 6626 35362 6638
rect 39678 6690 39730 6702
rect 41022 6690 41074 6702
rect 40338 6638 40350 6690
rect 40402 6638 40414 6690
rect 39678 6626 39730 6638
rect 41022 6626 41074 6638
rect 41358 6690 41410 6702
rect 41358 6626 41410 6638
rect 42590 6690 42642 6702
rect 45950 6690 46002 6702
rect 51550 6690 51602 6702
rect 43026 6638 43038 6690
rect 43090 6638 43102 6690
rect 51202 6638 51214 6690
rect 51266 6638 51278 6690
rect 42590 6626 42642 6638
rect 45950 6626 46002 6638
rect 51550 6626 51602 6638
rect 52558 6690 52610 6702
rect 52558 6626 52610 6638
rect 54574 6690 54626 6702
rect 54574 6626 54626 6638
rect 55582 6690 55634 6702
rect 55582 6626 55634 6638
rect 55806 6690 55858 6702
rect 55806 6626 55858 6638
rect 56030 6690 56082 6702
rect 56030 6626 56082 6638
rect 59726 6690 59778 6702
rect 59726 6626 59778 6638
rect 61294 6690 61346 6702
rect 62974 6690 63026 6702
rect 62066 6638 62078 6690
rect 62130 6638 62142 6690
rect 61294 6626 61346 6638
rect 62974 6626 63026 6638
rect 64766 6690 64818 6702
rect 67790 6690 67842 6702
rect 68350 6690 68402 6702
rect 72606 6690 72658 6702
rect 65650 6638 65662 6690
rect 65714 6638 65726 6690
rect 68002 6638 68014 6690
rect 68066 6638 68078 6690
rect 70018 6638 70030 6690
rect 70082 6638 70094 6690
rect 70914 6638 70926 6690
rect 70978 6638 70990 6690
rect 72146 6638 72158 6690
rect 72210 6638 72222 6690
rect 64766 6626 64818 6638
rect 67790 6626 67842 6638
rect 68350 6626 68402 6638
rect 72606 6626 72658 6638
rect 73166 6690 73218 6702
rect 77422 6690 77474 6702
rect 76066 6638 76078 6690
rect 76130 6638 76142 6690
rect 73166 6626 73218 6638
rect 77422 6626 77474 6638
rect 4398 6578 4450 6590
rect 1922 6526 1934 6578
rect 1986 6526 1998 6578
rect 4398 6514 4450 6526
rect 24110 6578 24162 6590
rect 24110 6514 24162 6526
rect 25230 6578 25282 6590
rect 25230 6514 25282 6526
rect 26798 6578 26850 6590
rect 26798 6514 26850 6526
rect 28142 6578 28194 6590
rect 28142 6514 28194 6526
rect 31054 6578 31106 6590
rect 31054 6514 31106 6526
rect 34862 6578 34914 6590
rect 34862 6514 34914 6526
rect 36094 6578 36146 6590
rect 36094 6514 36146 6526
rect 36430 6578 36482 6590
rect 36430 6514 36482 6526
rect 49982 6578 50034 6590
rect 49982 6514 50034 6526
rect 51438 6578 51490 6590
rect 51438 6514 51490 6526
rect 56702 6578 56754 6590
rect 56702 6514 56754 6526
rect 56814 6578 56866 6590
rect 56814 6514 56866 6526
rect 59166 6578 59218 6590
rect 59166 6514 59218 6526
rect 64430 6578 64482 6590
rect 77310 6578 77362 6590
rect 69682 6526 69694 6578
rect 69746 6526 69758 6578
rect 75058 6526 75070 6578
rect 75122 6526 75134 6578
rect 64430 6514 64482 6526
rect 77310 6514 77362 6526
rect 3726 6466 3778 6478
rect 3726 6402 3778 6414
rect 4510 6466 4562 6478
rect 4510 6402 4562 6414
rect 5630 6466 5682 6478
rect 5630 6402 5682 6414
rect 6078 6466 6130 6478
rect 6078 6402 6130 6414
rect 8878 6466 8930 6478
rect 8878 6402 8930 6414
rect 9550 6466 9602 6478
rect 9550 6402 9602 6414
rect 10110 6466 10162 6478
rect 10110 6402 10162 6414
rect 10334 6466 10386 6478
rect 10334 6402 10386 6414
rect 11342 6466 11394 6478
rect 11342 6402 11394 6414
rect 12014 6466 12066 6478
rect 12014 6402 12066 6414
rect 12686 6466 12738 6478
rect 12686 6402 12738 6414
rect 14254 6466 14306 6478
rect 14254 6402 14306 6414
rect 14366 6466 14418 6478
rect 14366 6402 14418 6414
rect 16270 6466 16322 6478
rect 16270 6402 16322 6414
rect 16494 6466 16546 6478
rect 16494 6402 16546 6414
rect 23214 6466 23266 6478
rect 23214 6402 23266 6414
rect 23774 6466 23826 6478
rect 23774 6402 23826 6414
rect 23886 6466 23938 6478
rect 23886 6402 23938 6414
rect 24894 6466 24946 6478
rect 24894 6402 24946 6414
rect 25118 6466 25170 6478
rect 25118 6402 25170 6414
rect 25790 6466 25842 6478
rect 25790 6402 25842 6414
rect 26910 6466 26962 6478
rect 26910 6402 26962 6414
rect 28030 6466 28082 6478
rect 28030 6402 28082 6414
rect 28814 6466 28866 6478
rect 28814 6402 28866 6414
rect 30046 6466 30098 6478
rect 30046 6402 30098 6414
rect 30606 6466 30658 6478
rect 30606 6402 30658 6414
rect 34190 6466 34242 6478
rect 34190 6402 34242 6414
rect 35086 6466 35138 6478
rect 35086 6402 35138 6414
rect 36206 6466 36258 6478
rect 36206 6402 36258 6414
rect 36766 6466 36818 6478
rect 36766 6402 36818 6414
rect 37438 6466 37490 6478
rect 37438 6402 37490 6414
rect 37886 6466 37938 6478
rect 37886 6402 37938 6414
rect 41246 6466 41298 6478
rect 41246 6402 41298 6414
rect 42142 6466 42194 6478
rect 42142 6402 42194 6414
rect 44382 6466 44434 6478
rect 44382 6402 44434 6414
rect 44718 6466 44770 6478
rect 44718 6402 44770 6414
rect 45390 6466 45442 6478
rect 45390 6402 45442 6414
rect 46510 6466 46562 6478
rect 46510 6402 46562 6414
rect 47070 6466 47122 6478
rect 47070 6402 47122 6414
rect 47406 6466 47458 6478
rect 47406 6402 47458 6414
rect 47854 6466 47906 6478
rect 47854 6402 47906 6414
rect 48302 6466 48354 6478
rect 48302 6402 48354 6414
rect 48750 6466 48802 6478
rect 48750 6402 48802 6414
rect 50094 6466 50146 6478
rect 50094 6402 50146 6414
rect 51326 6466 51378 6478
rect 51326 6402 51378 6414
rect 52110 6466 52162 6478
rect 52110 6402 52162 6414
rect 53342 6466 53394 6478
rect 53342 6402 53394 6414
rect 53902 6466 53954 6478
rect 53902 6402 53954 6414
rect 54686 6466 54738 6478
rect 54686 6402 54738 6414
rect 57038 6466 57090 6478
rect 57038 6402 57090 6414
rect 57374 6466 57426 6478
rect 57374 6402 57426 6414
rect 57822 6466 57874 6478
rect 57822 6402 57874 6414
rect 58382 6466 58434 6478
rect 58382 6402 58434 6414
rect 60174 6466 60226 6478
rect 60174 6402 60226 6414
rect 63422 6466 63474 6478
rect 63422 6402 63474 6414
rect 63870 6466 63922 6478
rect 63870 6402 63922 6414
rect 64542 6466 64594 6478
rect 64542 6402 64594 6414
rect 67006 6466 67058 6478
rect 67006 6402 67058 6414
rect 67678 6466 67730 6478
rect 67678 6402 67730 6414
rect 67902 6466 67954 6478
rect 72494 6466 72546 6478
rect 71474 6414 71486 6466
rect 71538 6414 71550 6466
rect 67902 6402 67954 6414
rect 72494 6402 72546 6414
rect 72718 6466 72770 6478
rect 72718 6402 72770 6414
rect 73614 6466 73666 6478
rect 73614 6402 73666 6414
rect 74062 6466 74114 6478
rect 74062 6402 74114 6414
rect 77534 6466 77586 6478
rect 77534 6402 77586 6414
rect 77758 6466 77810 6478
rect 77758 6402 77810 6414
rect 1344 6298 78784 6332
rect 1344 6246 20534 6298
rect 20586 6246 20638 6298
rect 20690 6246 20742 6298
rect 20794 6246 39854 6298
rect 39906 6246 39958 6298
rect 40010 6246 40062 6298
rect 40114 6246 59174 6298
rect 59226 6246 59278 6298
rect 59330 6246 59382 6298
rect 59434 6246 78494 6298
rect 78546 6246 78598 6298
rect 78650 6246 78702 6298
rect 78754 6246 78784 6298
rect 1344 6212 78784 6246
rect 2494 6130 2546 6142
rect 2494 6066 2546 6078
rect 10222 6130 10274 6142
rect 10222 6066 10274 6078
rect 10446 6130 10498 6142
rect 10446 6066 10498 6078
rect 11118 6130 11170 6142
rect 11118 6066 11170 6078
rect 15486 6130 15538 6142
rect 15486 6066 15538 6078
rect 16046 6130 16098 6142
rect 16046 6066 16098 6078
rect 16830 6130 16882 6142
rect 16830 6066 16882 6078
rect 22094 6130 22146 6142
rect 22094 6066 22146 6078
rect 23326 6130 23378 6142
rect 37326 6130 37378 6142
rect 35410 6078 35422 6130
rect 35474 6078 35486 6130
rect 23326 6066 23378 6078
rect 37326 6066 37378 6078
rect 45950 6130 46002 6142
rect 45950 6066 46002 6078
rect 46174 6130 46226 6142
rect 46174 6066 46226 6078
rect 48526 6130 48578 6142
rect 48526 6066 48578 6078
rect 48638 6130 48690 6142
rect 48638 6066 48690 6078
rect 51662 6130 51714 6142
rect 51662 6066 51714 6078
rect 52446 6130 52498 6142
rect 52446 6066 52498 6078
rect 53342 6130 53394 6142
rect 53342 6066 53394 6078
rect 55806 6130 55858 6142
rect 55806 6066 55858 6078
rect 56030 6130 56082 6142
rect 56030 6066 56082 6078
rect 58942 6130 58994 6142
rect 58942 6066 58994 6078
rect 59054 6130 59106 6142
rect 59054 6066 59106 6078
rect 62638 6130 62690 6142
rect 62638 6066 62690 6078
rect 62862 6130 62914 6142
rect 62862 6066 62914 6078
rect 66670 6130 66722 6142
rect 68574 6130 68626 6142
rect 67554 6078 67566 6130
rect 67618 6078 67630 6130
rect 66670 6066 66722 6078
rect 68574 6066 68626 6078
rect 69806 6130 69858 6142
rect 69806 6066 69858 6078
rect 70254 6130 70306 6142
rect 70254 6066 70306 6078
rect 70702 6130 70754 6142
rect 70702 6066 70754 6078
rect 73278 6130 73330 6142
rect 73278 6066 73330 6078
rect 74286 6130 74338 6142
rect 74286 6066 74338 6078
rect 74510 6130 74562 6142
rect 74510 6066 74562 6078
rect 77982 6130 78034 6142
rect 77982 6066 78034 6078
rect 4622 6018 4674 6030
rect 4622 5954 4674 5966
rect 7422 6018 7474 6030
rect 16158 6018 16210 6030
rect 12786 5966 12798 6018
rect 12850 5966 12862 6018
rect 7422 5954 7474 5966
rect 16158 5954 16210 5966
rect 18510 6018 18562 6030
rect 18510 5954 18562 5966
rect 21758 6018 21810 6030
rect 21758 5954 21810 5966
rect 36318 6018 36370 6030
rect 36318 5954 36370 5966
rect 36542 6018 36594 6030
rect 36542 5954 36594 5966
rect 39118 6018 39170 6030
rect 39118 5954 39170 5966
rect 49646 6018 49698 6030
rect 49646 5954 49698 5966
rect 49758 6018 49810 6030
rect 49758 5954 49810 5966
rect 51438 6018 51490 6030
rect 51438 5954 51490 5966
rect 57710 6018 57762 6030
rect 57710 5954 57762 5966
rect 57822 6018 57874 6030
rect 57822 5954 57874 5966
rect 62190 6018 62242 6030
rect 62190 5954 62242 5966
rect 62974 6018 63026 6030
rect 62974 5954 63026 5966
rect 63646 6018 63698 6030
rect 63646 5954 63698 5966
rect 63758 6018 63810 6030
rect 63758 5954 63810 5966
rect 66558 6018 66610 6030
rect 66558 5954 66610 5966
rect 68798 6018 68850 6030
rect 68798 5954 68850 5966
rect 68910 6018 68962 6030
rect 68910 5954 68962 5966
rect 75966 6018 76018 6030
rect 75966 5954 76018 5966
rect 76526 6018 76578 6030
rect 76526 5954 76578 5966
rect 3838 5906 3890 5918
rect 8430 5906 8482 5918
rect 3490 5854 3502 5906
rect 3554 5854 3566 5906
rect 5394 5854 5406 5906
rect 5458 5854 5470 5906
rect 6738 5854 6750 5906
rect 6802 5854 6814 5906
rect 3838 5842 3890 5854
rect 8430 5842 8482 5854
rect 8654 5906 8706 5918
rect 15822 5906 15874 5918
rect 13122 5854 13134 5906
rect 13186 5854 13198 5906
rect 14018 5854 14030 5906
rect 14082 5854 14094 5906
rect 8654 5842 8706 5854
rect 15822 5842 15874 5854
rect 18286 5906 18338 5918
rect 18286 5842 18338 5854
rect 18622 5906 18674 5918
rect 18622 5842 18674 5854
rect 21982 5906 22034 5918
rect 21982 5842 22034 5854
rect 22206 5906 22258 5918
rect 22206 5842 22258 5854
rect 22878 5906 22930 5918
rect 23550 5906 23602 5918
rect 23202 5854 23214 5906
rect 23266 5854 23278 5906
rect 22878 5842 22930 5854
rect 23550 5842 23602 5854
rect 24446 5906 24498 5918
rect 28142 5906 28194 5918
rect 30942 5906 30994 5918
rect 32734 5906 32786 5918
rect 27122 5854 27134 5906
rect 27186 5854 27198 5906
rect 28802 5854 28814 5906
rect 28866 5854 28878 5906
rect 30034 5854 30046 5906
rect 30098 5854 30110 5906
rect 32050 5854 32062 5906
rect 32114 5854 32126 5906
rect 32498 5854 32510 5906
rect 32562 5854 32574 5906
rect 24446 5842 24498 5854
rect 28142 5842 28194 5854
rect 30942 5842 30994 5854
rect 32734 5842 32786 5854
rect 35086 5906 35138 5918
rect 35086 5842 35138 5854
rect 36206 5906 36258 5918
rect 36206 5842 36258 5854
rect 38670 5906 38722 5918
rect 40798 5906 40850 5918
rect 39554 5854 39566 5906
rect 39618 5854 39630 5906
rect 38670 5842 38722 5854
rect 40798 5842 40850 5854
rect 42142 5906 42194 5918
rect 42142 5842 42194 5854
rect 42590 5906 42642 5918
rect 45838 5906 45890 5918
rect 44930 5854 44942 5906
rect 44994 5854 45006 5906
rect 42590 5842 42642 5854
rect 45838 5842 45890 5854
rect 46286 5906 46338 5918
rect 46286 5842 46338 5854
rect 48414 5906 48466 5918
rect 48414 5842 48466 5854
rect 51326 5906 51378 5918
rect 51326 5842 51378 5854
rect 51998 5906 52050 5918
rect 55918 5906 55970 5918
rect 54898 5854 54910 5906
rect 54962 5854 54974 5906
rect 55570 5854 55582 5906
rect 55634 5854 55646 5906
rect 51998 5842 52050 5854
rect 55918 5842 55970 5854
rect 56142 5906 56194 5918
rect 56142 5842 56194 5854
rect 58046 5906 58098 5918
rect 59166 5906 59218 5918
rect 66894 5906 66946 5918
rect 58818 5854 58830 5906
rect 58882 5854 58894 5906
rect 60050 5854 60062 5906
rect 60114 5854 60126 5906
rect 61506 5854 61518 5906
rect 61570 5854 61582 5906
rect 65874 5854 65886 5906
rect 65938 5854 65950 5906
rect 58046 5842 58098 5854
rect 59166 5842 59218 5854
rect 66894 5842 66946 5854
rect 67902 5906 67954 5918
rect 67902 5842 67954 5854
rect 68126 5906 68178 5918
rect 74174 5906 74226 5918
rect 72034 5854 72046 5906
rect 72098 5854 72110 5906
rect 72370 5854 72382 5906
rect 72434 5854 72446 5906
rect 75282 5854 75294 5906
rect 75346 5854 75358 5906
rect 76962 5854 76974 5906
rect 77026 5854 77038 5906
rect 68126 5842 68178 5854
rect 74174 5842 74226 5854
rect 9998 5794 10050 5806
rect 6626 5742 6638 5794
rect 6690 5742 6702 5794
rect 8978 5742 8990 5794
rect 9042 5742 9054 5794
rect 9998 5730 10050 5742
rect 10334 5794 10386 5806
rect 10334 5730 10386 5742
rect 11566 5794 11618 5806
rect 11566 5730 11618 5742
rect 12014 5794 12066 5806
rect 12014 5730 12066 5742
rect 14702 5794 14754 5806
rect 14702 5730 14754 5742
rect 17614 5794 17666 5806
rect 17614 5730 17666 5742
rect 19070 5794 19122 5806
rect 19070 5730 19122 5742
rect 19518 5794 19570 5806
rect 19518 5730 19570 5742
rect 19966 5794 20018 5806
rect 19966 5730 20018 5742
rect 23438 5794 23490 5806
rect 23438 5730 23490 5742
rect 24894 5794 24946 5806
rect 24894 5730 24946 5742
rect 25678 5794 25730 5806
rect 25678 5730 25730 5742
rect 26238 5794 26290 5806
rect 33854 5794 33906 5806
rect 26674 5742 26686 5794
rect 26738 5742 26750 5794
rect 30370 5742 30382 5794
rect 30434 5742 30446 5794
rect 26238 5730 26290 5742
rect 33854 5730 33906 5742
rect 34414 5794 34466 5806
rect 34414 5730 34466 5742
rect 34862 5794 34914 5806
rect 34862 5730 34914 5742
rect 36878 5794 36930 5806
rect 36878 5730 36930 5742
rect 37774 5794 37826 5806
rect 43150 5794 43202 5806
rect 39442 5742 39454 5794
rect 39506 5742 39518 5794
rect 41682 5742 41694 5794
rect 41746 5742 41758 5794
rect 37774 5730 37826 5742
rect 43150 5730 43202 5742
rect 43486 5794 43538 5806
rect 43486 5730 43538 5742
rect 44158 5794 44210 5806
rect 46062 5794 46114 5806
rect 44818 5742 44830 5794
rect 44882 5742 44894 5794
rect 44158 5730 44210 5742
rect 46062 5730 46114 5742
rect 46846 5794 46898 5806
rect 46846 5730 46898 5742
rect 47294 5794 47346 5806
rect 47294 5730 47346 5742
rect 48190 5794 48242 5806
rect 48190 5730 48242 5742
rect 50206 5794 50258 5806
rect 50206 5730 50258 5742
rect 50654 5794 50706 5806
rect 50654 5730 50706 5742
rect 52894 5794 52946 5806
rect 52894 5730 52946 5742
rect 53790 5794 53842 5806
rect 53790 5730 53842 5742
rect 54462 5794 54514 5806
rect 54462 5730 54514 5742
rect 56702 5794 56754 5806
rect 56702 5730 56754 5742
rect 58494 5794 58546 5806
rect 64206 5794 64258 5806
rect 59938 5742 59950 5794
rect 60002 5742 60014 5794
rect 58494 5730 58546 5742
rect 64206 5730 64258 5742
rect 64654 5794 64706 5806
rect 69358 5794 69410 5806
rect 65538 5742 65550 5794
rect 65602 5742 65614 5794
rect 64654 5730 64706 5742
rect 69358 5730 69410 5742
rect 72606 5794 72658 5806
rect 75058 5742 75070 5794
rect 75122 5742 75134 5794
rect 77298 5742 77310 5794
rect 77362 5742 77374 5794
rect 72606 5730 72658 5742
rect 9774 5682 9826 5694
rect 47966 5682 48018 5694
rect 3602 5630 3614 5682
rect 3666 5630 3678 5682
rect 25554 5630 25566 5682
rect 25618 5679 25630 5682
rect 26450 5679 26462 5682
rect 25618 5633 26462 5679
rect 25618 5630 25630 5633
rect 26450 5630 26462 5633
rect 26514 5630 26526 5682
rect 9774 5618 9826 5630
rect 47966 5618 48018 5630
rect 49646 5682 49698 5694
rect 49646 5618 49698 5630
rect 63646 5682 63698 5694
rect 63646 5618 63698 5630
rect 1344 5514 78624 5548
rect 1344 5462 10874 5514
rect 10926 5462 10978 5514
rect 11030 5462 11082 5514
rect 11134 5462 30194 5514
rect 30246 5462 30298 5514
rect 30350 5462 30402 5514
rect 30454 5462 49514 5514
rect 49566 5462 49618 5514
rect 49670 5462 49722 5514
rect 49774 5462 68834 5514
rect 68886 5462 68938 5514
rect 68990 5462 69042 5514
rect 69094 5462 78624 5514
rect 1344 5428 78624 5462
rect 8654 5346 8706 5358
rect 14030 5346 14082 5358
rect 39790 5346 39842 5358
rect 13682 5294 13694 5346
rect 13746 5294 13758 5346
rect 22194 5294 22206 5346
rect 22258 5294 22270 5346
rect 25442 5294 25454 5346
rect 25506 5294 25518 5346
rect 27458 5294 27470 5346
rect 27522 5343 27534 5346
rect 28802 5343 28814 5346
rect 27522 5297 28814 5343
rect 27522 5294 27534 5297
rect 28802 5294 28814 5297
rect 28866 5294 28878 5346
rect 8654 5282 8706 5294
rect 14030 5282 14082 5294
rect 39790 5282 39842 5294
rect 46398 5346 46450 5358
rect 53566 5346 53618 5358
rect 49186 5294 49198 5346
rect 49250 5294 49262 5346
rect 46398 5282 46450 5294
rect 53566 5282 53618 5294
rect 56590 5346 56642 5358
rect 59042 5294 59054 5346
rect 59106 5343 59118 5346
rect 59266 5343 59278 5346
rect 59106 5297 59278 5343
rect 59106 5294 59118 5297
rect 59266 5294 59278 5297
rect 59330 5343 59342 5346
rect 60162 5343 60174 5346
rect 59330 5297 60174 5343
rect 59330 5294 59342 5297
rect 60162 5294 60174 5297
rect 60226 5294 60238 5346
rect 72482 5294 72494 5346
rect 72546 5294 72558 5346
rect 76290 5294 76302 5346
rect 76354 5294 76366 5346
rect 56590 5282 56642 5294
rect 4510 5234 4562 5246
rect 4510 5170 4562 5182
rect 7646 5234 7698 5246
rect 7646 5170 7698 5182
rect 7982 5234 8034 5246
rect 7982 5170 8034 5182
rect 9326 5234 9378 5246
rect 9326 5170 9378 5182
rect 9886 5234 9938 5246
rect 13022 5234 13074 5246
rect 10546 5182 10558 5234
rect 10610 5182 10622 5234
rect 9886 5170 9938 5182
rect 13022 5170 13074 5182
rect 14254 5234 14306 5246
rect 14254 5170 14306 5182
rect 14926 5234 14978 5246
rect 27470 5234 27522 5246
rect 21970 5182 21982 5234
rect 22034 5182 22046 5234
rect 14926 5170 14978 5182
rect 27470 5170 27522 5182
rect 27918 5234 27970 5246
rect 27918 5170 27970 5182
rect 32286 5234 32338 5246
rect 32286 5170 32338 5182
rect 34078 5234 34130 5246
rect 34078 5170 34130 5182
rect 39118 5234 39170 5246
rect 39118 5170 39170 5182
rect 42478 5234 42530 5246
rect 42478 5170 42530 5182
rect 42926 5234 42978 5246
rect 57598 5234 57650 5246
rect 47730 5182 47742 5234
rect 47794 5182 47806 5234
rect 50418 5182 50430 5234
rect 50482 5182 50494 5234
rect 42926 5170 42978 5182
rect 57598 5170 57650 5182
rect 59278 5234 59330 5246
rect 59278 5170 59330 5182
rect 61966 5234 62018 5246
rect 64878 5234 64930 5246
rect 64306 5182 64318 5234
rect 64370 5182 64382 5234
rect 61966 5170 62018 5182
rect 64878 5170 64930 5182
rect 69246 5234 69298 5246
rect 69246 5170 69298 5182
rect 69694 5234 69746 5246
rect 69694 5170 69746 5182
rect 70590 5234 70642 5246
rect 73502 5234 73554 5246
rect 77198 5234 77250 5246
rect 71698 5182 71710 5234
rect 71762 5182 71774 5234
rect 75618 5182 75630 5234
rect 75682 5182 75694 5234
rect 70590 5170 70642 5182
rect 73502 5170 73554 5182
rect 77198 5170 77250 5182
rect 4846 5122 4898 5134
rect 12126 5122 12178 5134
rect 2930 5070 2942 5122
rect 2994 5070 3006 5122
rect 3826 5070 3838 5122
rect 3890 5070 3902 5122
rect 10658 5070 10670 5122
rect 10722 5070 10734 5122
rect 4846 5058 4898 5070
rect 12126 5058 12178 5070
rect 15150 5122 15202 5134
rect 15150 5058 15202 5070
rect 17054 5122 17106 5134
rect 17054 5058 17106 5070
rect 17502 5122 17554 5134
rect 17502 5058 17554 5070
rect 18846 5122 18898 5134
rect 18846 5058 18898 5070
rect 19182 5122 19234 5134
rect 19182 5058 19234 5070
rect 20526 5122 20578 5134
rect 24558 5122 24610 5134
rect 26462 5122 26514 5134
rect 22530 5070 22542 5122
rect 22594 5070 22606 5122
rect 23874 5070 23886 5122
rect 23938 5070 23950 5122
rect 25554 5070 25566 5122
rect 25618 5070 25630 5122
rect 20526 5058 20578 5070
rect 24558 5058 24610 5070
rect 26462 5058 26514 5070
rect 28366 5122 28418 5134
rect 28366 5058 28418 5070
rect 28926 5122 28978 5134
rect 28926 5058 28978 5070
rect 29710 5122 29762 5134
rect 29710 5058 29762 5070
rect 30046 5122 30098 5134
rect 30046 5058 30098 5070
rect 30494 5122 30546 5134
rect 30494 5058 30546 5070
rect 33518 5122 33570 5134
rect 38110 5122 38162 5134
rect 35186 5070 35198 5122
rect 35250 5070 35262 5122
rect 33518 5058 33570 5070
rect 38110 5058 38162 5070
rect 38558 5122 38610 5134
rect 41022 5122 41074 5134
rect 40114 5070 40126 5122
rect 40178 5070 40190 5122
rect 38558 5058 38610 5070
rect 41022 5058 41074 5070
rect 41470 5122 41522 5134
rect 41470 5058 41522 5070
rect 43374 5122 43426 5134
rect 43374 5058 43426 5070
rect 44494 5122 44546 5134
rect 44494 5058 44546 5070
rect 45390 5122 45442 5134
rect 51774 5122 51826 5134
rect 55358 5122 55410 5134
rect 47618 5070 47630 5122
rect 47682 5070 47694 5122
rect 49298 5070 49310 5122
rect 49362 5070 49374 5122
rect 51090 5070 51102 5122
rect 51154 5070 51166 5122
rect 52098 5070 52110 5122
rect 52162 5070 52174 5122
rect 45390 5058 45442 5070
rect 51774 5058 51826 5070
rect 55358 5058 55410 5070
rect 57150 5122 57202 5134
rect 57150 5058 57202 5070
rect 60734 5122 60786 5134
rect 60734 5058 60786 5070
rect 62526 5122 62578 5134
rect 62526 5058 62578 5070
rect 63422 5122 63474 5134
rect 63422 5058 63474 5070
rect 65774 5122 65826 5134
rect 65774 5058 65826 5070
rect 66558 5122 66610 5134
rect 66558 5058 66610 5070
rect 67678 5122 67730 5134
rect 67678 5058 67730 5070
rect 67902 5122 67954 5134
rect 67902 5058 67954 5070
rect 70254 5122 70306 5134
rect 73950 5122 74002 5134
rect 77646 5122 77698 5134
rect 72034 5070 72046 5122
rect 72098 5070 72110 5122
rect 75506 5070 75518 5122
rect 75570 5070 75582 5122
rect 70254 5058 70306 5070
rect 73950 5058 74002 5070
rect 77646 5058 77698 5070
rect 78094 5122 78146 5134
rect 78094 5058 78146 5070
rect 8654 5010 8706 5022
rect 1922 4958 1934 5010
rect 1986 4958 1998 5010
rect 8654 4946 8706 4958
rect 8766 5010 8818 5022
rect 8766 4946 8818 4958
rect 11342 5010 11394 5022
rect 11342 4946 11394 4958
rect 16494 5010 16546 5022
rect 16494 4946 16546 4958
rect 16606 5010 16658 5022
rect 16606 4946 16658 4958
rect 18510 5010 18562 5022
rect 18510 4946 18562 4958
rect 29822 5010 29874 5022
rect 29822 4946 29874 4958
rect 30830 5010 30882 5022
rect 30830 4946 30882 4958
rect 32958 5010 33010 5022
rect 36766 5010 36818 5022
rect 34850 4958 34862 5010
rect 34914 4958 34926 5010
rect 36530 4958 36542 5010
rect 36594 4958 36606 5010
rect 32958 4946 33010 4958
rect 36766 4946 36818 4958
rect 39006 5010 39058 5022
rect 39006 4946 39058 4958
rect 40462 5010 40514 5022
rect 40462 4946 40514 4958
rect 44718 5010 44770 5022
rect 44718 4946 44770 4958
rect 45614 5010 45666 5022
rect 45614 4946 45666 4958
rect 45726 5010 45778 5022
rect 45726 4946 45778 4958
rect 46510 5010 46562 5022
rect 46510 4946 46562 4958
rect 53678 5010 53730 5022
rect 53678 4946 53730 4958
rect 54798 5010 54850 5022
rect 54798 4946 54850 4958
rect 56590 5010 56642 5022
rect 56590 4946 56642 4958
rect 56702 5010 56754 5022
rect 56702 4946 56754 4958
rect 58606 5010 58658 5022
rect 58606 4946 58658 4958
rect 60398 5010 60450 5022
rect 60398 4946 60450 4958
rect 60510 5010 60562 5022
rect 60510 4946 60562 4958
rect 63086 5010 63138 5022
rect 63086 4946 63138 4958
rect 65438 5010 65490 5022
rect 65438 4946 65490 4958
rect 65550 5010 65602 5022
rect 65550 4946 65602 4958
rect 66222 5010 66274 5022
rect 66222 4946 66274 4958
rect 68238 5010 68290 5022
rect 68238 4946 68290 4958
rect 3614 4898 3666 4910
rect 3614 4834 3666 4846
rect 11790 4898 11842 4910
rect 11790 4834 11842 4846
rect 12014 4898 12066 4910
rect 16270 4898 16322 4910
rect 15474 4846 15486 4898
rect 15538 4846 15550 4898
rect 12014 4834 12066 4846
rect 16270 4834 16322 4846
rect 17950 4898 18002 4910
rect 17950 4834 18002 4846
rect 18622 4898 18674 4910
rect 18622 4834 18674 4846
rect 19854 4898 19906 4910
rect 19854 4834 19906 4846
rect 19966 4898 20018 4910
rect 19966 4834 20018 4846
rect 20078 4898 20130 4910
rect 20078 4834 20130 4846
rect 20974 4898 21026 4910
rect 20974 4834 21026 4846
rect 27022 4898 27074 4910
rect 27022 4834 27074 4846
rect 30718 4898 30770 4910
rect 30718 4834 30770 4846
rect 31278 4898 31330 4910
rect 31278 4834 31330 4846
rect 31950 4898 32002 4910
rect 31950 4834 32002 4846
rect 32846 4898 32898 4910
rect 32846 4834 32898 4846
rect 33070 4898 33122 4910
rect 33070 4834 33122 4846
rect 37774 4898 37826 4910
rect 37774 4834 37826 4846
rect 39230 4898 39282 4910
rect 39230 4834 39282 4846
rect 40238 4898 40290 4910
rect 40238 4834 40290 4846
rect 40350 4898 40402 4910
rect 40350 4834 40402 4846
rect 41918 4898 41970 4910
rect 41918 4834 41970 4846
rect 44158 4898 44210 4910
rect 44158 4834 44210 4846
rect 44270 4898 44322 4910
rect 44270 4834 44322 4846
rect 44382 4898 44434 4910
rect 44382 4834 44434 4846
rect 46398 4898 46450 4910
rect 46398 4834 46450 4846
rect 53566 4898 53618 4910
rect 53566 4834 53618 4846
rect 54462 4898 54514 4910
rect 54462 4834 54514 4846
rect 54686 4898 54738 4910
rect 54686 4834 54738 4846
rect 55918 4898 55970 4910
rect 55918 4834 55970 4846
rect 58046 4898 58098 4910
rect 58046 4834 58098 4846
rect 58718 4898 58770 4910
rect 58718 4834 58770 4846
rect 58942 4898 58994 4910
rect 58942 4834 58994 4846
rect 59726 4898 59778 4910
rect 59726 4834 59778 4846
rect 61294 4898 61346 4910
rect 61294 4834 61346 4846
rect 63198 4898 63250 4910
rect 63198 4834 63250 4846
rect 63870 4898 63922 4910
rect 63870 4834 63922 4846
rect 66334 4898 66386 4910
rect 66334 4834 66386 4846
rect 66894 4898 66946 4910
rect 66894 4834 66946 4846
rect 68126 4898 68178 4910
rect 68126 4834 68178 4846
rect 68350 4898 68402 4910
rect 68350 4834 68402 4846
rect 73054 4898 73106 4910
rect 73054 4834 73106 4846
rect 74398 4898 74450 4910
rect 74398 4834 74450 4846
rect 1344 4730 78784 4764
rect 1344 4678 20534 4730
rect 20586 4678 20638 4730
rect 20690 4678 20742 4730
rect 20794 4678 39854 4730
rect 39906 4678 39958 4730
rect 40010 4678 40062 4730
rect 40114 4678 59174 4730
rect 59226 4678 59278 4730
rect 59330 4678 59382 4730
rect 59434 4678 78494 4730
rect 78546 4678 78598 4730
rect 78650 4678 78702 4730
rect 78754 4678 78784 4730
rect 1344 4644 78784 4678
rect 3614 4562 3666 4574
rect 3614 4498 3666 4510
rect 13806 4562 13858 4574
rect 17054 4562 17106 4574
rect 16370 4510 16382 4562
rect 16434 4510 16446 4562
rect 13806 4498 13858 4510
rect 17054 4498 17106 4510
rect 21086 4562 21138 4574
rect 21086 4498 21138 4510
rect 22094 4562 22146 4574
rect 22094 4498 22146 4510
rect 23438 4562 23490 4574
rect 23438 4498 23490 4510
rect 23774 4562 23826 4574
rect 23774 4498 23826 4510
rect 24558 4562 24610 4574
rect 24558 4498 24610 4510
rect 26126 4562 26178 4574
rect 26126 4498 26178 4510
rect 26350 4562 26402 4574
rect 26350 4498 26402 4510
rect 27246 4562 27298 4574
rect 27246 4498 27298 4510
rect 31278 4562 31330 4574
rect 31278 4498 31330 4510
rect 35534 4562 35586 4574
rect 35534 4498 35586 4510
rect 37886 4562 37938 4574
rect 37886 4498 37938 4510
rect 38110 4562 38162 4574
rect 38110 4498 38162 4510
rect 41694 4562 41746 4574
rect 41694 4498 41746 4510
rect 41918 4562 41970 4574
rect 41918 4498 41970 4510
rect 42702 4562 42754 4574
rect 42702 4498 42754 4510
rect 46958 4562 47010 4574
rect 46958 4498 47010 4510
rect 47518 4562 47570 4574
rect 47518 4498 47570 4510
rect 48414 4562 48466 4574
rect 48414 4498 48466 4510
rect 48638 4562 48690 4574
rect 48638 4498 48690 4510
rect 50542 4562 50594 4574
rect 50542 4498 50594 4510
rect 53006 4562 53058 4574
rect 53006 4498 53058 4510
rect 53678 4562 53730 4574
rect 57934 4562 57986 4574
rect 56466 4510 56478 4562
rect 56530 4510 56542 4562
rect 53678 4498 53730 4510
rect 57934 4498 57986 4510
rect 59614 4562 59666 4574
rect 59614 4498 59666 4510
rect 61518 4562 61570 4574
rect 61518 4498 61570 4510
rect 64430 4562 64482 4574
rect 72606 4562 72658 4574
rect 64430 4498 64482 4510
rect 71934 4506 71986 4518
rect 3950 4450 4002 4462
rect 3950 4386 4002 4398
rect 4510 4450 4562 4462
rect 4510 4386 4562 4398
rect 9886 4450 9938 4462
rect 9886 4386 9938 4398
rect 10558 4450 10610 4462
rect 10558 4386 10610 4398
rect 12798 4450 12850 4462
rect 21310 4450 21362 4462
rect 14802 4398 14814 4450
rect 14866 4398 14878 4450
rect 16258 4398 16270 4450
rect 16322 4398 16334 4450
rect 12798 4386 12850 4398
rect 21310 4386 21362 4398
rect 21982 4450 22034 4462
rect 21982 4386 22034 4398
rect 23998 4450 24050 4462
rect 23998 4386 24050 4398
rect 24110 4450 24162 4462
rect 24110 4386 24162 4398
rect 24782 4450 24834 4462
rect 24782 4386 24834 4398
rect 24894 4450 24946 4462
rect 24894 4386 24946 4398
rect 27694 4450 27746 4462
rect 27694 4386 27746 4398
rect 32846 4450 32898 4462
rect 32846 4386 32898 4398
rect 35646 4450 35698 4462
rect 35646 4386 35698 4398
rect 40350 4450 40402 4462
rect 40350 4386 40402 4398
rect 40462 4450 40514 4462
rect 40462 4386 40514 4398
rect 42030 4450 42082 4462
rect 42030 4386 42082 4398
rect 42254 4450 42306 4462
rect 47406 4450 47458 4462
rect 43474 4398 43486 4450
rect 43538 4398 43550 4450
rect 42254 4386 42306 4398
rect 47406 4386 47458 4398
rect 49758 4450 49810 4462
rect 49758 4386 49810 4398
rect 50094 4450 50146 4462
rect 50094 4386 50146 4398
rect 50766 4450 50818 4462
rect 50766 4386 50818 4398
rect 51550 4450 51602 4462
rect 51550 4386 51602 4398
rect 51662 4450 51714 4462
rect 57710 4450 57762 4462
rect 54786 4398 54798 4450
rect 54850 4398 54862 4450
rect 51662 4386 51714 4398
rect 57710 4386 57762 4398
rect 58942 4450 58994 4462
rect 58942 4386 58994 4398
rect 59054 4450 59106 4462
rect 59054 4386 59106 4398
rect 59838 4450 59890 4462
rect 59838 4386 59890 4398
rect 59950 4450 60002 4462
rect 59950 4386 60002 4398
rect 60398 4450 60450 4462
rect 68238 4450 68290 4462
rect 63522 4398 63534 4450
rect 63586 4398 63598 4450
rect 60398 4386 60450 4398
rect 68238 4386 68290 4398
rect 71374 4450 71426 4462
rect 72606 4498 72658 4510
rect 73278 4562 73330 4574
rect 73278 4498 73330 4510
rect 74062 4562 74114 4574
rect 74062 4498 74114 4510
rect 71934 4442 71986 4454
rect 72046 4450 72098 4462
rect 71374 4386 71426 4398
rect 72046 4386 72098 4398
rect 76750 4450 76802 4462
rect 76750 4386 76802 4398
rect 77086 4450 77138 4462
rect 77086 4386 77138 4398
rect 77646 4450 77698 4462
rect 77646 4386 77698 4398
rect 77982 4450 78034 4462
rect 77982 4386 78034 4398
rect 8654 4338 8706 4350
rect 12238 4338 12290 4350
rect 21422 4338 21474 4350
rect 3042 4286 3054 4338
rect 3106 4286 3118 4338
rect 11442 4286 11454 4338
rect 11506 4286 11518 4338
rect 14914 4286 14926 4338
rect 14978 4286 14990 4338
rect 17938 4286 17950 4338
rect 18002 4286 18014 4338
rect 20402 4286 20414 4338
rect 20466 4286 20478 4338
rect 8654 4274 8706 4286
rect 12238 4274 12290 4286
rect 21422 4274 21474 4286
rect 25678 4338 25730 4350
rect 27358 4338 27410 4350
rect 26002 4286 26014 4338
rect 26066 4286 26078 4338
rect 27010 4286 27022 4338
rect 27074 4286 27086 4338
rect 25678 4274 25730 4286
rect 27358 4274 27410 4286
rect 27470 4338 27522 4350
rect 32734 4338 32786 4350
rect 29138 4286 29150 4338
rect 29202 4286 29214 4338
rect 30146 4286 30158 4338
rect 30210 4286 30222 4338
rect 32162 4286 32174 4338
rect 32226 4286 32238 4338
rect 27470 4274 27522 4286
rect 32734 4274 32786 4286
rect 33630 4338 33682 4350
rect 35310 4338 35362 4350
rect 37774 4338 37826 4350
rect 41806 4338 41858 4350
rect 34066 4286 34078 4338
rect 34130 4286 34142 4338
rect 36754 4286 36766 4338
rect 36818 4286 36830 4338
rect 39442 4286 39454 4338
rect 39506 4286 39518 4338
rect 33630 4274 33682 4286
rect 35310 4274 35362 4286
rect 37774 4274 37826 4286
rect 41806 4274 41858 4286
rect 48750 4338 48802 4350
rect 48750 4274 48802 4286
rect 50878 4338 50930 4350
rect 50878 4274 50930 4286
rect 51326 4338 51378 4350
rect 51326 4274 51378 4286
rect 52446 4338 52498 4350
rect 52446 4274 52498 4286
rect 55134 4338 55186 4350
rect 55134 4274 55186 4286
rect 56142 4338 56194 4350
rect 56142 4274 56194 4286
rect 58046 4338 58098 4350
rect 58046 4274 58098 4286
rect 58158 4338 58210 4350
rect 61294 4338 61346 4350
rect 61966 4338 62018 4350
rect 74398 4338 74450 4350
rect 58370 4286 58382 4338
rect 58434 4286 58446 4338
rect 61618 4286 61630 4338
rect 61682 4286 61694 4338
rect 65650 4286 65662 4338
rect 65714 4286 65726 4338
rect 66994 4286 67006 4338
rect 67058 4286 67070 4338
rect 69570 4286 69582 4338
rect 69634 4286 69646 4338
rect 70914 4286 70926 4338
rect 70978 4286 70990 4338
rect 76178 4286 76190 4338
rect 76242 4286 76254 4338
rect 58158 4274 58210 4286
rect 61294 4274 61346 4286
rect 61966 4274 62018 4286
rect 74398 4274 74450 4286
rect 9102 4226 9154 4238
rect 13358 4226 13410 4238
rect 18958 4226 19010 4238
rect 22878 4226 22930 4238
rect 1922 4174 1934 4226
rect 1986 4174 1998 4226
rect 11106 4174 11118 4226
rect 11170 4174 11182 4226
rect 18274 4174 18286 4226
rect 18338 4174 18350 4226
rect 20290 4174 20302 4226
rect 20354 4174 20366 4226
rect 9102 4162 9154 4174
rect 13358 4162 13410 4174
rect 18958 4162 19010 4174
rect 22878 4162 22930 4174
rect 26238 4226 26290 4238
rect 36206 4226 36258 4238
rect 38670 4226 38722 4238
rect 55582 4226 55634 4238
rect 30594 4174 30606 4226
rect 30658 4174 30670 4226
rect 34402 4174 34414 4226
rect 34466 4174 34478 4226
rect 37090 4174 37102 4226
rect 37154 4174 37166 4226
rect 38882 4174 38894 4226
rect 38946 4174 38958 4226
rect 54114 4174 54126 4226
rect 54178 4174 54190 4226
rect 26238 4162 26290 4174
rect 36206 4162 36258 4174
rect 38670 4162 38722 4174
rect 55582 4162 55634 4174
rect 61406 4226 61458 4238
rect 62514 4174 62526 4226
rect 62578 4174 62590 4226
rect 65874 4174 65886 4226
rect 65938 4174 65950 4226
rect 69122 4174 69134 4226
rect 69186 4174 69198 4226
rect 75506 4174 75518 4226
rect 75570 4174 75582 4226
rect 61406 4162 61458 4174
rect 9998 4114 10050 4126
rect 22094 4114 22146 4126
rect 40350 4114 40402 4126
rect 20066 4062 20078 4114
rect 20130 4062 20142 4114
rect 28466 4062 28478 4114
rect 28530 4062 28542 4114
rect 9998 4050 10050 4062
rect 22094 4050 22146 4062
rect 40350 4050 40402 4062
rect 47518 4114 47570 4126
rect 47518 4050 47570 4062
rect 59054 4114 59106 4126
rect 72046 4114 72098 4126
rect 67666 4062 67678 4114
rect 67730 4062 67742 4114
rect 59054 4050 59106 4062
rect 72046 4050 72098 4062
rect 1344 3946 78624 3980
rect 1344 3894 10874 3946
rect 10926 3894 10978 3946
rect 11030 3894 11082 3946
rect 11134 3894 30194 3946
rect 30246 3894 30298 3946
rect 30350 3894 30402 3946
rect 30454 3894 49514 3946
rect 49566 3894 49618 3946
rect 49670 3894 49722 3946
rect 49774 3894 68834 3946
rect 68886 3894 68938 3946
rect 68990 3894 69042 3946
rect 69094 3894 78624 3946
rect 1344 3860 78624 3894
rect 34190 3778 34242 3790
rect 34190 3714 34242 3726
rect 42926 3778 42978 3790
rect 42926 3714 42978 3726
rect 59614 3778 59666 3790
rect 59614 3714 59666 3726
rect 67342 3778 67394 3790
rect 67666 3726 67678 3778
rect 67730 3726 67742 3778
rect 67342 3714 67394 3726
rect 15486 3666 15538 3678
rect 20526 3666 20578 3678
rect 4946 3614 4958 3666
rect 5010 3614 5022 3666
rect 7186 3614 7198 3666
rect 7250 3614 7262 3666
rect 10322 3614 10334 3666
rect 10386 3614 10398 3666
rect 14018 3614 14030 3666
rect 14082 3614 14094 3666
rect 18498 3614 18510 3666
rect 18562 3614 18574 3666
rect 20066 3614 20078 3666
rect 20130 3614 20142 3666
rect 15486 3602 15538 3614
rect 20526 3602 20578 3614
rect 21646 3666 21698 3678
rect 21646 3602 21698 3614
rect 22654 3666 22706 3678
rect 25454 3666 25506 3678
rect 24098 3614 24110 3666
rect 24162 3614 24174 3666
rect 22654 3602 22706 3614
rect 25454 3602 25506 3614
rect 27246 3666 27298 3678
rect 27246 3602 27298 3614
rect 27694 3666 27746 3678
rect 27694 3602 27746 3614
rect 28142 3666 28194 3678
rect 28142 3602 28194 3614
rect 30158 3666 30210 3678
rect 30158 3602 30210 3614
rect 31950 3666 32002 3678
rect 31950 3602 32002 3614
rect 38670 3666 38722 3678
rect 38670 3602 38722 3614
rect 45166 3666 45218 3678
rect 45166 3602 45218 3614
rect 45502 3666 45554 3678
rect 45502 3602 45554 3614
rect 46846 3666 46898 3678
rect 46846 3602 46898 3614
rect 47406 3666 47458 3678
rect 47406 3602 47458 3614
rect 53342 3666 53394 3678
rect 53342 3602 53394 3614
rect 53902 3666 53954 3678
rect 53902 3602 53954 3614
rect 55022 3666 55074 3678
rect 55022 3602 55074 3614
rect 63534 3666 63586 3678
rect 67118 3666 67170 3678
rect 72382 3666 72434 3678
rect 76302 3666 76354 3678
rect 65090 3614 65102 3666
rect 65154 3614 65166 3666
rect 68898 3614 68910 3666
rect 68962 3614 68974 3666
rect 74834 3614 74846 3666
rect 74898 3614 74910 3666
rect 63534 3602 63586 3614
rect 67118 3602 67170 3614
rect 72382 3602 72434 3614
rect 76302 3602 76354 3614
rect 77310 3666 77362 3678
rect 77310 3602 77362 3614
rect 5630 3554 5682 3566
rect 11454 3554 11506 3566
rect 2146 3502 2158 3554
rect 2210 3502 2222 3554
rect 9650 3502 9662 3554
rect 9714 3502 9726 3554
rect 5630 3490 5682 3502
rect 11454 3490 11506 3502
rect 11678 3554 11730 3566
rect 11678 3490 11730 3502
rect 13582 3554 13634 3566
rect 13582 3490 13634 3502
rect 15262 3554 15314 3566
rect 15262 3490 15314 3502
rect 15710 3554 15762 3566
rect 15710 3490 15762 3502
rect 16606 3554 16658 3566
rect 16606 3490 16658 3502
rect 17502 3554 17554 3566
rect 17502 3490 17554 3502
rect 17950 3554 18002 3566
rect 22094 3554 22146 3566
rect 18834 3502 18846 3554
rect 18898 3502 18910 3554
rect 19842 3502 19854 3554
rect 19906 3502 19918 3554
rect 17950 3490 18002 3502
rect 22094 3490 22146 3502
rect 24558 3554 24610 3566
rect 24558 3490 24610 3502
rect 25902 3554 25954 3566
rect 25902 3490 25954 3502
rect 29262 3554 29314 3566
rect 29262 3490 29314 3502
rect 32510 3554 32562 3566
rect 32510 3490 32562 3502
rect 34302 3554 34354 3566
rect 34302 3490 34354 3502
rect 34862 3554 34914 3566
rect 34862 3490 34914 3502
rect 35982 3554 36034 3566
rect 35982 3490 36034 3502
rect 37102 3554 37154 3566
rect 37102 3490 37154 3502
rect 38222 3554 38274 3566
rect 38222 3490 38274 3502
rect 39118 3554 39170 3566
rect 39118 3490 39170 3502
rect 39902 3554 39954 3566
rect 39902 3490 39954 3502
rect 40238 3554 40290 3566
rect 40238 3490 40290 3502
rect 42814 3554 42866 3566
rect 42814 3490 42866 3502
rect 43598 3554 43650 3566
rect 44942 3554 44994 3566
rect 44034 3502 44046 3554
rect 44098 3502 44110 3554
rect 43598 3490 43650 3502
rect 44942 3490 44994 3502
rect 45390 3554 45442 3566
rect 45390 3490 45442 3502
rect 52782 3554 52834 3566
rect 52782 3490 52834 3502
rect 54462 3554 54514 3566
rect 56926 3554 56978 3566
rect 55458 3502 55470 3554
rect 55522 3502 55534 3554
rect 54462 3490 54514 3502
rect 56926 3490 56978 3502
rect 57486 3554 57538 3566
rect 57486 3490 57538 3502
rect 59502 3554 59554 3566
rect 66558 3554 66610 3566
rect 64754 3502 64766 3554
rect 64818 3502 64830 3554
rect 59502 3490 59554 3502
rect 66558 3490 66610 3502
rect 68350 3554 68402 3566
rect 73378 3502 73390 3554
rect 73442 3502 73454 3554
rect 75506 3502 75518 3554
rect 75570 3502 75582 3554
rect 76738 3502 76750 3554
rect 76802 3502 76814 3554
rect 68350 3490 68402 3502
rect 6750 3442 6802 3454
rect 11566 3442 11618 3454
rect 2818 3390 2830 3442
rect 2882 3390 2894 3442
rect 8194 3390 8206 3442
rect 8258 3390 8270 3442
rect 6750 3378 6802 3390
rect 11566 3378 11618 3390
rect 11902 3442 11954 3454
rect 11902 3378 11954 3390
rect 12910 3442 12962 3454
rect 12910 3378 12962 3390
rect 15038 3442 15090 3454
rect 15038 3378 15090 3390
rect 23550 3442 23602 3454
rect 23550 3378 23602 3390
rect 26350 3442 26402 3454
rect 26350 3378 26402 3390
rect 28590 3442 28642 3454
rect 28590 3378 28642 3390
rect 30606 3442 30658 3454
rect 31614 3442 31666 3454
rect 30930 3390 30942 3442
rect 30994 3390 31006 3442
rect 30606 3378 30658 3390
rect 31614 3378 31666 3390
rect 33182 3442 33234 3454
rect 33182 3378 33234 3390
rect 34190 3442 34242 3454
rect 34190 3378 34242 3390
rect 36430 3442 36482 3454
rect 36430 3378 36482 3390
rect 39454 3442 39506 3454
rect 39454 3378 39506 3390
rect 41246 3442 41298 3454
rect 41246 3378 41298 3390
rect 42030 3442 42082 3454
rect 42030 3378 42082 3390
rect 46286 3442 46338 3454
rect 46286 3378 46338 3390
rect 47966 3442 48018 3454
rect 47966 3378 48018 3390
rect 48750 3442 48802 3454
rect 51774 3442 51826 3454
rect 50978 3390 50990 3442
rect 51042 3390 51054 3442
rect 48750 3378 48802 3390
rect 51774 3378 51826 3390
rect 58046 3442 58098 3454
rect 58942 3442 58994 3454
rect 65662 3442 65714 3454
rect 71374 3442 71426 3454
rect 58594 3390 58606 3442
rect 58658 3390 58670 3442
rect 62962 3390 62974 3442
rect 63026 3390 63038 3442
rect 66210 3390 66222 3442
rect 66274 3390 66286 3442
rect 70242 3390 70254 3442
rect 70306 3390 70318 3442
rect 58046 3378 58098 3390
rect 58942 3378 58994 3390
rect 65662 3378 65714 3390
rect 71374 3378 71426 3390
rect 77758 3442 77810 3454
rect 77758 3378 77810 3390
rect 15150 3330 15202 3342
rect 26686 3330 26738 3342
rect 33518 3330 33570 3342
rect 16258 3278 16270 3330
rect 16322 3278 16334 3330
rect 29586 3278 29598 3330
rect 29650 3278 29662 3330
rect 15150 3266 15202 3278
rect 26686 3266 26738 3278
rect 33518 3266 33570 3278
rect 35198 3330 35250 3342
rect 40126 3330 40178 3342
rect 37426 3278 37438 3330
rect 37490 3278 37502 3330
rect 35198 3266 35250 3278
rect 40126 3266 40178 3278
rect 41582 3330 41634 3342
rect 41582 3266 41634 3278
rect 42926 3330 42978 3342
rect 42926 3266 42978 3278
rect 45614 3330 45666 3342
rect 45614 3266 45666 3278
rect 56590 3330 56642 3342
rect 56590 3266 56642 3278
rect 56814 3330 56866 3342
rect 56814 3266 56866 3278
rect 59614 3330 59666 3342
rect 59614 3266 59666 3278
rect 60510 3330 60562 3342
rect 73166 3330 73218 3342
rect 71026 3278 71038 3330
rect 71090 3278 71102 3330
rect 60510 3266 60562 3278
rect 73166 3266 73218 3278
rect 1344 3162 78784 3196
rect 1344 3110 20534 3162
rect 20586 3110 20638 3162
rect 20690 3110 20742 3162
rect 20794 3110 39854 3162
rect 39906 3110 39958 3162
rect 40010 3110 40062 3162
rect 40114 3110 59174 3162
rect 59226 3110 59278 3162
rect 59330 3110 59382 3162
rect 59434 3110 78494 3162
rect 78546 3110 78598 3162
rect 78650 3110 78702 3162
rect 78754 3110 78784 3162
rect 1344 3076 78784 3110
<< via1 >>
rect 10874 36822 10926 36874
rect 10978 36822 11030 36874
rect 11082 36822 11134 36874
rect 30194 36822 30246 36874
rect 30298 36822 30350 36874
rect 30402 36822 30454 36874
rect 49514 36822 49566 36874
rect 49618 36822 49670 36874
rect 49722 36822 49774 36874
rect 68834 36822 68886 36874
rect 68938 36822 68990 36874
rect 69042 36822 69094 36874
rect 2046 36542 2098 36594
rect 4174 36542 4226 36594
rect 6974 36542 7026 36594
rect 9774 36542 9826 36594
rect 11790 36542 11842 36594
rect 14366 36542 14418 36594
rect 19294 36542 19346 36594
rect 21646 36542 21698 36594
rect 23886 36542 23938 36594
rect 26686 36542 26738 36594
rect 29374 36542 29426 36594
rect 31278 36542 31330 36594
rect 33518 36542 33570 36594
rect 34078 36542 34130 36594
rect 37214 36542 37266 36594
rect 41470 36542 41522 36594
rect 46398 36542 46450 36594
rect 48974 36542 49026 36594
rect 50990 36542 51042 36594
rect 54350 36542 54402 36594
rect 56814 36542 56866 36594
rect 58830 36542 58882 36594
rect 61742 36542 61794 36594
rect 64654 36542 64706 36594
rect 66446 36542 66498 36594
rect 68574 36542 68626 36594
rect 70702 36542 70754 36594
rect 74062 36542 74114 36594
rect 76974 36542 77026 36594
rect 77982 36542 78034 36594
rect 3166 36430 3218 36482
rect 4958 36430 5010 36482
rect 8094 36430 8146 36482
rect 10670 36430 10722 36482
rect 12574 36430 12626 36482
rect 13694 36430 13746 36482
rect 15486 36430 15538 36482
rect 17502 36430 17554 36482
rect 17726 36430 17778 36482
rect 17950 36430 18002 36482
rect 20414 36430 20466 36482
rect 22766 36430 22818 36482
rect 24558 36430 24610 36482
rect 27806 36430 27858 36482
rect 30494 36430 30546 36482
rect 32398 36430 32450 36482
rect 35198 36430 35250 36482
rect 35646 36430 35698 36482
rect 35870 36430 35922 36482
rect 36206 36430 36258 36482
rect 37438 36430 37490 36482
rect 38670 36430 38722 36482
rect 42590 36430 42642 36482
rect 47518 36430 47570 36482
rect 49870 36430 49922 36482
rect 51886 36430 51938 36482
rect 53678 36430 53730 36482
rect 57710 36430 57762 36482
rect 59838 36430 59890 36482
rect 61294 36430 61346 36482
rect 65774 36430 65826 36482
rect 67566 36430 67618 36482
rect 69470 36430 69522 36482
rect 71374 36430 71426 36482
rect 73390 36430 73442 36482
rect 75406 36430 75458 36482
rect 76302 36430 76354 36482
rect 16718 36318 16770 36370
rect 18062 36318 18114 36370
rect 25790 36318 25842 36370
rect 28590 36318 28642 36370
rect 36094 36318 36146 36370
rect 39454 36318 39506 36370
rect 43822 36318 43874 36370
rect 44158 36318 44210 36370
rect 52782 36318 52834 36370
rect 62862 36318 62914 36370
rect 63198 36318 63250 36370
rect 72494 36318 72546 36370
rect 5630 36206 5682 36258
rect 6078 36206 6130 36258
rect 8542 36206 8594 36258
rect 16382 36206 16434 36258
rect 18734 36206 18786 36258
rect 25230 36206 25282 36258
rect 25902 36206 25954 36258
rect 26126 36206 26178 36258
rect 43038 36206 43090 36258
rect 45054 36206 45106 36258
rect 45278 36206 45330 36258
rect 45390 36206 45442 36258
rect 45502 36206 45554 36258
rect 47966 36206 48018 36258
rect 53118 36206 53170 36258
rect 60510 36206 60562 36258
rect 63870 36206 63922 36258
rect 72830 36206 72882 36258
rect 75182 36206 75234 36258
rect 20534 36038 20586 36090
rect 20638 36038 20690 36090
rect 20742 36038 20794 36090
rect 39854 36038 39906 36090
rect 39958 36038 40010 36090
rect 40062 36038 40114 36090
rect 59174 36038 59226 36090
rect 59278 36038 59330 36090
rect 59382 36038 59434 36090
rect 78494 36038 78546 36090
rect 78598 36038 78650 36090
rect 78702 36038 78754 36090
rect 5294 35870 5346 35922
rect 14366 35870 14418 35922
rect 24894 35870 24946 35922
rect 26798 35870 26850 35922
rect 27470 35870 27522 35922
rect 28478 35870 28530 35922
rect 31166 35870 31218 35922
rect 33966 35870 34018 35922
rect 40574 35870 40626 35922
rect 49758 35870 49810 35922
rect 53342 35870 53394 35922
rect 60062 35870 60114 35922
rect 67454 35870 67506 35922
rect 67902 35870 67954 35922
rect 70478 35870 70530 35922
rect 71710 35870 71762 35922
rect 73278 35870 73330 35922
rect 1934 35758 1986 35810
rect 3614 35758 3666 35810
rect 4510 35758 4562 35810
rect 4846 35758 4898 35810
rect 12014 35758 12066 35810
rect 15038 35758 15090 35810
rect 17838 35758 17890 35810
rect 28590 35758 28642 35810
rect 34862 35758 34914 35810
rect 34974 35758 35026 35810
rect 36542 35758 36594 35810
rect 39006 35758 39058 35810
rect 42702 35758 42754 35810
rect 43934 35758 43986 35810
rect 52110 35758 52162 35810
rect 62974 35758 63026 35810
rect 72270 35758 72322 35810
rect 72606 35758 72658 35810
rect 74398 35758 74450 35810
rect 76078 35758 76130 35810
rect 77870 35758 77922 35810
rect 3054 35646 3106 35698
rect 3950 35646 4002 35698
rect 11006 35646 11058 35698
rect 11454 35646 11506 35698
rect 11902 35646 11954 35698
rect 12238 35646 12290 35698
rect 12686 35646 12738 35698
rect 12910 35646 12962 35698
rect 13582 35646 13634 35698
rect 16382 35646 16434 35698
rect 18846 35646 18898 35698
rect 19742 35646 19794 35698
rect 19966 35646 20018 35698
rect 21982 35646 22034 35698
rect 22430 35646 22482 35698
rect 23326 35646 23378 35698
rect 23998 35646 24050 35698
rect 24558 35646 24610 35698
rect 26462 35646 26514 35698
rect 27358 35646 27410 35698
rect 28478 35646 28530 35698
rect 29374 35646 29426 35698
rect 29598 35646 29650 35698
rect 29822 35646 29874 35698
rect 31054 35646 31106 35698
rect 31390 35646 31442 35698
rect 32398 35646 32450 35698
rect 32734 35646 32786 35698
rect 32846 35646 32898 35698
rect 33630 35646 33682 35698
rect 35086 35646 35138 35698
rect 37662 35646 37714 35698
rect 40126 35646 40178 35698
rect 41806 35646 41858 35698
rect 44942 35646 44994 35698
rect 45614 35646 45666 35698
rect 46062 35646 46114 35698
rect 47854 35646 47906 35698
rect 48078 35646 48130 35698
rect 51438 35646 51490 35698
rect 51998 35646 52050 35698
rect 55358 35646 55410 35698
rect 55918 35646 55970 35698
rect 56030 35646 56082 35698
rect 56142 35646 56194 35698
rect 59166 35646 59218 35698
rect 61406 35646 61458 35698
rect 61854 35646 61906 35698
rect 64206 35646 64258 35698
rect 64430 35646 64482 35698
rect 64766 35646 64818 35698
rect 65662 35646 65714 35698
rect 66558 35646 66610 35698
rect 67118 35646 67170 35698
rect 70814 35646 70866 35698
rect 74174 35646 74226 35698
rect 74958 35646 75010 35698
rect 76750 35646 76802 35698
rect 10446 35534 10498 35586
rect 15150 35534 15202 35586
rect 16046 35534 16098 35586
rect 16718 35534 16770 35586
rect 19518 35534 19570 35586
rect 21534 35534 21586 35586
rect 23102 35534 23154 35586
rect 26238 35534 26290 35586
rect 38110 35534 38162 35586
rect 42030 35534 42082 35586
rect 46510 35534 46562 35586
rect 48750 35534 48802 35586
rect 50542 35534 50594 35586
rect 52558 35534 52610 35586
rect 56590 35534 56642 35586
rect 57486 35534 57538 35586
rect 58046 35534 58098 35586
rect 58942 35534 58994 35586
rect 60510 35534 60562 35586
rect 62302 35534 62354 35586
rect 62862 35534 62914 35586
rect 64542 35534 64594 35586
rect 65774 35534 65826 35586
rect 68350 35534 68402 35586
rect 69022 35534 69074 35586
rect 69694 35534 69746 35586
rect 71262 35534 71314 35586
rect 14814 35422 14866 35474
rect 35534 35422 35586 35474
rect 49534 35422 49586 35474
rect 49870 35422 49922 35474
rect 57710 35422 57762 35474
rect 59390 35422 59442 35474
rect 59614 35422 59666 35474
rect 60622 35422 60674 35474
rect 63198 35422 63250 35474
rect 69582 35422 69634 35474
rect 10874 35254 10926 35306
rect 10978 35254 11030 35306
rect 11082 35254 11134 35306
rect 30194 35254 30246 35306
rect 30298 35254 30350 35306
rect 30402 35254 30454 35306
rect 49514 35254 49566 35306
rect 49618 35254 49670 35306
rect 49722 35254 49774 35306
rect 68834 35254 68886 35306
rect 68938 35254 68990 35306
rect 69042 35254 69094 35306
rect 15038 35086 15090 35138
rect 19742 35086 19794 35138
rect 20078 35086 20130 35138
rect 22654 35086 22706 35138
rect 22990 35086 23042 35138
rect 26014 35086 26066 35138
rect 32062 35086 32114 35138
rect 47182 35086 47234 35138
rect 48190 35086 48242 35138
rect 48302 35086 48354 35138
rect 48526 35086 48578 35138
rect 57374 35086 57426 35138
rect 58158 35086 58210 35138
rect 59166 35086 59218 35138
rect 64990 35086 65042 35138
rect 2158 34974 2210 35026
rect 4398 34974 4450 35026
rect 4846 34974 4898 35026
rect 11678 34974 11730 35026
rect 12014 34974 12066 35026
rect 13918 34974 13970 35026
rect 14142 34974 14194 35026
rect 17278 34974 17330 35026
rect 19518 34974 19570 35026
rect 21870 34974 21922 35026
rect 27470 34974 27522 35026
rect 27918 34974 27970 35026
rect 31390 34974 31442 35026
rect 42590 34974 42642 35026
rect 44718 34974 44770 35026
rect 46174 34974 46226 35026
rect 55694 34974 55746 35026
rect 57038 34974 57090 35026
rect 58158 34974 58210 35026
rect 62750 34974 62802 35026
rect 66222 34974 66274 35026
rect 69470 34974 69522 35026
rect 74062 34974 74114 35026
rect 76078 34974 76130 35026
rect 3054 34862 3106 34914
rect 3950 34862 4002 34914
rect 11342 34862 11394 34914
rect 12686 34862 12738 34914
rect 14366 34862 14418 34914
rect 14590 34862 14642 34914
rect 16382 34862 16434 34914
rect 16830 34862 16882 34914
rect 18958 34862 19010 34914
rect 20526 34862 20578 34914
rect 23550 34862 23602 34914
rect 23886 34862 23938 34914
rect 25342 34862 25394 34914
rect 26574 34862 26626 34914
rect 26798 34862 26850 34914
rect 28814 34862 28866 34914
rect 31278 34862 31330 34914
rect 34750 34862 34802 34914
rect 35198 34862 35250 34914
rect 35646 34862 35698 34914
rect 36542 34862 36594 34914
rect 39790 34862 39842 34914
rect 40350 34862 40402 34914
rect 40462 34862 40514 34914
rect 41358 34862 41410 34914
rect 44046 34862 44098 34914
rect 47182 34862 47234 34914
rect 49982 34862 50034 34914
rect 50878 34862 50930 34914
rect 55246 34862 55298 34914
rect 56030 34862 56082 34914
rect 56590 34862 56642 34914
rect 57262 34862 57314 34914
rect 59054 34862 59106 34914
rect 59726 34862 59778 34914
rect 62526 34862 62578 34914
rect 64990 34862 65042 34914
rect 65326 34862 65378 34914
rect 65550 34862 65602 34914
rect 65998 34862 66050 34914
rect 66670 34862 66722 34914
rect 73278 34862 73330 34914
rect 74958 34862 75010 34914
rect 12910 34750 12962 34802
rect 15822 34750 15874 34802
rect 18622 34750 18674 34802
rect 22430 34750 22482 34802
rect 23662 34750 23714 34802
rect 28478 34750 28530 34802
rect 30494 34750 30546 34802
rect 36206 34750 36258 34802
rect 36654 34750 36706 34802
rect 36766 34750 36818 34802
rect 37550 34750 37602 34802
rect 42814 34750 42866 34802
rect 46622 34750 46674 34802
rect 47518 34750 47570 34802
rect 48638 34750 48690 34802
rect 49758 34750 49810 34802
rect 51774 34750 51826 34802
rect 52110 34750 52162 34802
rect 56814 34750 56866 34802
rect 63198 34750 63250 34802
rect 63982 34750 64034 34802
rect 66446 34750 66498 34802
rect 69694 34750 69746 34802
rect 71374 34750 71426 34802
rect 72158 34750 72210 34802
rect 72270 34750 72322 34802
rect 72494 34750 72546 34802
rect 77310 34750 77362 34802
rect 78094 34750 78146 34802
rect 3614 34638 3666 34690
rect 18174 34638 18226 34690
rect 25006 34638 25058 34690
rect 25678 34638 25730 34690
rect 25902 34638 25954 34690
rect 29598 34638 29650 34690
rect 30270 34638 30322 34690
rect 30382 34638 30434 34690
rect 32622 34638 32674 34690
rect 37662 34638 37714 34690
rect 37774 34638 37826 34690
rect 41470 34638 41522 34690
rect 41694 34638 41746 34690
rect 45390 34638 45442 34690
rect 49198 34638 49250 34690
rect 50318 34638 50370 34690
rect 51214 34638 51266 34690
rect 57598 34638 57650 34690
rect 61294 34638 61346 34690
rect 64094 34638 64146 34690
rect 64766 34638 64818 34690
rect 67118 34638 67170 34690
rect 71262 34638 71314 34690
rect 73614 34638 73666 34690
rect 77646 34638 77698 34690
rect 20534 34470 20586 34522
rect 20638 34470 20690 34522
rect 20742 34470 20794 34522
rect 39854 34470 39906 34522
rect 39958 34470 40010 34522
rect 40062 34470 40114 34522
rect 59174 34470 59226 34522
rect 59278 34470 59330 34522
rect 59382 34470 59434 34522
rect 78494 34470 78546 34522
rect 78598 34470 78650 34522
rect 78702 34470 78754 34522
rect 12350 34302 12402 34354
rect 15598 34302 15650 34354
rect 16494 34302 16546 34354
rect 17838 34302 17890 34354
rect 18622 34302 18674 34354
rect 18846 34302 18898 34354
rect 26238 34302 26290 34354
rect 27470 34302 27522 34354
rect 30718 34302 30770 34354
rect 31502 34302 31554 34354
rect 33854 34302 33906 34354
rect 37438 34302 37490 34354
rect 39790 34302 39842 34354
rect 40462 34302 40514 34354
rect 40686 34302 40738 34354
rect 42478 34302 42530 34354
rect 43486 34302 43538 34354
rect 58270 34302 58322 34354
rect 59726 34302 59778 34354
rect 62750 34302 62802 34354
rect 65774 34302 65826 34354
rect 70142 34302 70194 34354
rect 72382 34302 72434 34354
rect 73614 34302 73666 34354
rect 8990 34190 9042 34242
rect 13470 34190 13522 34242
rect 13806 34190 13858 34242
rect 14590 34190 14642 34242
rect 16942 34190 16994 34242
rect 17726 34190 17778 34242
rect 17950 34190 18002 34242
rect 21982 34190 22034 34242
rect 24894 34190 24946 34242
rect 26014 34190 26066 34242
rect 27134 34190 27186 34242
rect 27246 34190 27298 34242
rect 31278 34190 31330 34242
rect 35758 34190 35810 34242
rect 39454 34190 39506 34242
rect 40350 34190 40402 34242
rect 43934 34190 43986 34242
rect 51550 34190 51602 34242
rect 51774 34190 51826 34242
rect 52446 34190 52498 34242
rect 52558 34190 52610 34242
rect 53902 34190 53954 34242
rect 55134 34190 55186 34242
rect 59390 34190 59442 34242
rect 59502 34190 59554 34242
rect 60174 34190 60226 34242
rect 62974 34190 63026 34242
rect 65662 34190 65714 34242
rect 71150 34190 71202 34242
rect 74062 34190 74114 34242
rect 74398 34190 74450 34242
rect 76750 34190 76802 34242
rect 77086 34190 77138 34242
rect 77646 34190 77698 34242
rect 3054 34078 3106 34130
rect 7198 34078 7250 34130
rect 8206 34078 8258 34130
rect 13022 34078 13074 34130
rect 13246 34078 13298 34130
rect 13694 34078 13746 34130
rect 18958 34078 19010 34130
rect 20078 34078 20130 34130
rect 21198 34078 21250 34130
rect 23326 34078 23378 34130
rect 23886 34078 23938 34130
rect 26238 34078 26290 34130
rect 26462 34078 26514 34130
rect 32846 34078 32898 34130
rect 33742 34078 33794 34130
rect 33966 34078 34018 34130
rect 34302 34078 34354 34130
rect 35422 34078 35474 34130
rect 43150 34078 43202 34130
rect 43598 34078 43650 34130
rect 50654 34078 50706 34130
rect 51886 34078 51938 34130
rect 52782 34078 52834 34130
rect 53790 34078 53842 34130
rect 57710 34078 57762 34130
rect 57934 34078 57986 34130
rect 58158 34078 58210 34130
rect 58382 34078 58434 34130
rect 60286 34078 60338 34130
rect 60510 34078 60562 34130
rect 60622 34078 60674 34130
rect 63086 34078 63138 34130
rect 65998 34078 66050 34130
rect 70254 34078 70306 34130
rect 70926 34078 70978 34130
rect 74958 34078 75010 34130
rect 77982 34078 78034 34130
rect 1934 33966 1986 34018
rect 6750 33966 6802 34018
rect 9662 33966 9714 34018
rect 14702 33966 14754 34018
rect 15150 33966 15202 34018
rect 20190 33966 20242 34018
rect 22990 33966 23042 34018
rect 24334 33966 24386 34018
rect 35198 33966 35250 34018
rect 37550 33966 37602 34018
rect 42590 33966 42642 34018
rect 50318 33966 50370 34018
rect 51102 33966 51154 34018
rect 53118 33966 53170 34018
rect 55246 33966 55298 34018
rect 57486 33966 57538 34018
rect 71822 33966 71874 34018
rect 76078 33966 76130 34018
rect 14366 33854 14418 33906
rect 31614 33854 31666 33906
rect 37214 33854 37266 33906
rect 42254 33854 42306 33906
rect 43486 33854 43538 33906
rect 53902 33854 53954 33906
rect 54910 33854 54962 33906
rect 70142 33854 70194 33906
rect 10874 33686 10926 33738
rect 10978 33686 11030 33738
rect 11082 33686 11134 33738
rect 30194 33686 30246 33738
rect 30298 33686 30350 33738
rect 30402 33686 30454 33738
rect 49514 33686 49566 33738
rect 49618 33686 49670 33738
rect 49722 33686 49774 33738
rect 68834 33686 68886 33738
rect 68938 33686 68990 33738
rect 69042 33686 69094 33738
rect 13806 33518 13858 33570
rect 23550 33518 23602 33570
rect 23886 33518 23938 33570
rect 30606 33518 30658 33570
rect 42814 33518 42866 33570
rect 61518 33518 61570 33570
rect 63198 33518 63250 33570
rect 65102 33518 65154 33570
rect 72270 33518 72322 33570
rect 73950 33518 74002 33570
rect 74398 33518 74450 33570
rect 3614 33406 3666 33458
rect 6750 33406 6802 33458
rect 8766 33406 8818 33458
rect 9774 33406 9826 33458
rect 14366 33406 14418 33458
rect 17278 33406 17330 33458
rect 21982 33406 22034 33458
rect 22430 33406 22482 33458
rect 22766 33406 22818 33458
rect 23326 33406 23378 33458
rect 28366 33406 28418 33458
rect 29934 33406 29986 33458
rect 32062 33406 32114 33458
rect 34974 33406 35026 33458
rect 37886 33406 37938 33458
rect 40126 33406 40178 33458
rect 42590 33406 42642 33458
rect 43934 33406 43986 33458
rect 47294 33406 47346 33458
rect 47742 33406 47794 33458
rect 49310 33406 49362 33458
rect 53790 33406 53842 33458
rect 55694 33406 55746 33458
rect 71150 33406 71202 33458
rect 73166 33406 73218 33458
rect 74398 33406 74450 33458
rect 75630 33406 75682 33458
rect 3166 33294 3218 33346
rect 8206 33294 8258 33346
rect 9662 33294 9714 33346
rect 10334 33294 10386 33346
rect 12014 33294 12066 33346
rect 12686 33294 12738 33346
rect 12910 33294 12962 33346
rect 17950 33294 18002 33346
rect 18174 33294 18226 33346
rect 19742 33294 19794 33346
rect 20414 33294 20466 33346
rect 28254 33294 28306 33346
rect 28926 33294 28978 33346
rect 29822 33294 29874 33346
rect 32846 33294 32898 33346
rect 33518 33294 33570 33346
rect 34190 33294 34242 33346
rect 37998 33294 38050 33346
rect 39342 33294 39394 33346
rect 43150 33294 43202 33346
rect 44270 33294 44322 33346
rect 48190 33294 48242 33346
rect 48414 33294 48466 33346
rect 49646 33294 49698 33346
rect 49870 33294 49922 33346
rect 50430 33294 50482 33346
rect 50766 33294 50818 33346
rect 50990 33294 51042 33346
rect 54126 33294 54178 33346
rect 54574 33294 54626 33346
rect 56142 33294 56194 33346
rect 56590 33294 56642 33346
rect 57150 33294 57202 33346
rect 57710 33294 57762 33346
rect 57822 33294 57874 33346
rect 64206 33294 64258 33346
rect 65438 33294 65490 33346
rect 66558 33294 66610 33346
rect 67118 33294 67170 33346
rect 70254 33294 70306 33346
rect 70590 33294 70642 33346
rect 71934 33294 71986 33346
rect 73950 33294 74002 33346
rect 75070 33294 75122 33346
rect 76414 33294 76466 33346
rect 77534 33294 77586 33346
rect 7198 33182 7250 33234
rect 13694 33182 13746 33234
rect 13806 33182 13858 33234
rect 18846 33182 18898 33234
rect 44718 33182 44770 33234
rect 45502 33182 45554 33234
rect 45614 33182 45666 33234
rect 45838 33182 45890 33234
rect 51774 33182 51826 33234
rect 60510 33182 60562 33234
rect 61630 33182 61682 33234
rect 62526 33182 62578 33234
rect 63086 33182 63138 33234
rect 63870 33182 63922 33234
rect 63982 33182 64034 33234
rect 65662 33182 65714 33234
rect 67230 33182 67282 33234
rect 71710 33182 71762 33234
rect 2830 33070 2882 33122
rect 9438 33070 9490 33122
rect 9886 33070 9938 33122
rect 19966 33070 20018 33122
rect 28478 33070 28530 33122
rect 36878 33070 36930 33122
rect 51438 33070 51490 33122
rect 51662 33070 51714 33122
rect 52334 33070 52386 33122
rect 52782 33070 52834 33122
rect 57598 33070 57650 33122
rect 59166 33070 59218 33122
rect 60622 33070 60674 33122
rect 61518 33070 61570 33122
rect 74846 33070 74898 33122
rect 76190 33070 76242 33122
rect 77310 33070 77362 33122
rect 78094 33070 78146 33122
rect 20534 32902 20586 32954
rect 20638 32902 20690 32954
rect 20742 32902 20794 32954
rect 39854 32902 39906 32954
rect 39958 32902 40010 32954
rect 40062 32902 40114 32954
rect 59174 32902 59226 32954
rect 59278 32902 59330 32954
rect 59382 32902 59434 32954
rect 78494 32902 78546 32954
rect 78598 32902 78650 32954
rect 78702 32902 78754 32954
rect 3614 32734 3666 32786
rect 7422 32734 7474 32786
rect 7646 32734 7698 32786
rect 8206 32734 8258 32786
rect 8318 32734 8370 32786
rect 8990 32734 9042 32786
rect 13134 32734 13186 32786
rect 17614 32734 17666 32786
rect 17838 32734 17890 32786
rect 29486 32734 29538 32786
rect 34190 32734 34242 32786
rect 38558 32734 38610 32786
rect 38670 32734 38722 32786
rect 39230 32734 39282 32786
rect 42366 32734 42418 32786
rect 48078 32734 48130 32786
rect 49870 32734 49922 32786
rect 50654 32734 50706 32786
rect 56030 32734 56082 32786
rect 57934 32734 57986 32786
rect 58494 32734 58546 32786
rect 63534 32734 63586 32786
rect 67230 32734 67282 32786
rect 69582 32734 69634 32786
rect 74286 32734 74338 32786
rect 2830 32622 2882 32674
rect 3166 32622 3218 32674
rect 7310 32622 7362 32674
rect 8094 32622 8146 32674
rect 12798 32622 12850 32674
rect 14926 32622 14978 32674
rect 17950 32622 18002 32674
rect 19742 32622 19794 32674
rect 22654 32622 22706 32674
rect 24894 32622 24946 32674
rect 33630 32622 33682 32674
rect 46622 32622 46674 32674
rect 49758 32622 49810 32674
rect 50094 32622 50146 32674
rect 52222 32622 52274 32674
rect 55918 32622 55970 32674
rect 57486 32622 57538 32674
rect 58718 32622 58770 32674
rect 58830 32622 58882 32674
rect 59278 32622 59330 32674
rect 60286 32622 60338 32674
rect 66446 32622 66498 32674
rect 67454 32622 67506 32674
rect 70478 32622 70530 32674
rect 74734 32622 74786 32674
rect 76526 32622 76578 32674
rect 77198 32622 77250 32674
rect 77534 32622 77586 32674
rect 77982 32622 78034 32674
rect 13022 32510 13074 32562
rect 13246 32510 13298 32562
rect 14030 32510 14082 32562
rect 18846 32510 18898 32562
rect 19070 32510 19122 32562
rect 22430 32510 22482 32562
rect 24446 32510 24498 32562
rect 27470 32510 27522 32562
rect 28926 32510 28978 32562
rect 31166 32510 31218 32562
rect 31502 32510 31554 32562
rect 31726 32510 31778 32562
rect 33854 32510 33906 32562
rect 37326 32510 37378 32562
rect 38110 32510 38162 32562
rect 38782 32510 38834 32562
rect 47630 32510 47682 32562
rect 49534 32510 49586 32562
rect 51550 32510 51602 32562
rect 55358 32510 55410 32562
rect 55694 32510 55746 32562
rect 56366 32510 56418 32562
rect 57710 32510 57762 32562
rect 58158 32510 58210 32562
rect 60062 32510 60114 32562
rect 60398 32510 60450 32562
rect 61518 32510 61570 32562
rect 62190 32510 62242 32562
rect 63198 32510 63250 32562
rect 63534 32510 63586 32562
rect 63758 32510 63810 32562
rect 66782 32510 66834 32562
rect 67566 32510 67618 32562
rect 69918 32510 69970 32562
rect 70590 32510 70642 32562
rect 71150 32510 71202 32562
rect 74846 32510 74898 32562
rect 75182 32510 75234 32562
rect 4174 32398 4226 32450
rect 14142 32398 14194 32450
rect 16046 32398 16098 32450
rect 23438 32398 23490 32450
rect 23998 32398 24050 32450
rect 27582 32398 27634 32450
rect 28254 32398 28306 32450
rect 31390 32398 31442 32450
rect 37102 32398 37154 32450
rect 37662 32398 37714 32450
rect 42254 32398 42306 32450
rect 45390 32398 45442 32450
rect 46174 32398 46226 32450
rect 51438 32398 51490 32450
rect 53790 32398 53842 32450
rect 54350 32398 54402 32450
rect 61742 32398 61794 32450
rect 62638 32398 62690 32450
rect 66670 32398 66722 32450
rect 4398 32286 4450 32338
rect 4734 32286 4786 32338
rect 29150 32286 29202 32338
rect 54574 32286 54626 32338
rect 54910 32286 54962 32338
rect 76302 32286 76354 32338
rect 76638 32286 76690 32338
rect 10874 32118 10926 32170
rect 10978 32118 11030 32170
rect 11082 32118 11134 32170
rect 30194 32118 30246 32170
rect 30298 32118 30350 32170
rect 30402 32118 30454 32170
rect 49514 32118 49566 32170
rect 49618 32118 49670 32170
rect 49722 32118 49774 32170
rect 68834 32118 68886 32170
rect 68938 32118 68990 32170
rect 69042 32118 69094 32170
rect 14142 31950 14194 32002
rect 27582 31950 27634 32002
rect 37774 31950 37826 32002
rect 59166 31950 59218 32002
rect 60398 31950 60450 32002
rect 70254 31950 70306 32002
rect 73390 31950 73442 32002
rect 4958 31838 5010 31890
rect 9214 31838 9266 31890
rect 11454 31838 11506 31890
rect 16942 31838 16994 31890
rect 17726 31838 17778 31890
rect 20302 31838 20354 31890
rect 22654 31838 22706 31890
rect 23998 31838 24050 31890
rect 26910 31838 26962 31890
rect 31614 31838 31666 31890
rect 33406 31838 33458 31890
rect 33742 31838 33794 31890
rect 37550 31838 37602 31890
rect 38110 31838 38162 31890
rect 40126 31838 40178 31890
rect 41806 31838 41858 31890
rect 44046 31838 44098 31890
rect 46510 31838 46562 31890
rect 61742 31838 61794 31890
rect 63870 31838 63922 31890
rect 65886 31838 65938 31890
rect 74286 31838 74338 31890
rect 75518 31838 75570 31890
rect 77310 31838 77362 31890
rect 78094 31838 78146 31890
rect 2942 31726 2994 31778
rect 4622 31726 4674 31778
rect 5630 31726 5682 31778
rect 9326 31726 9378 31778
rect 10670 31726 10722 31778
rect 13918 31726 13970 31778
rect 14142 31726 14194 31778
rect 17054 31726 17106 31778
rect 20638 31726 20690 31778
rect 20862 31726 20914 31778
rect 21758 31726 21810 31778
rect 21982 31726 22034 31778
rect 24894 31726 24946 31778
rect 27246 31726 27298 31778
rect 31278 31726 31330 31778
rect 32174 31726 32226 31778
rect 33182 31726 33234 31778
rect 39678 31726 39730 31778
rect 41022 31726 41074 31778
rect 43598 31726 43650 31778
rect 43822 31726 43874 31778
rect 46174 31726 46226 31778
rect 46398 31726 46450 31778
rect 47630 31726 47682 31778
rect 49758 31726 49810 31778
rect 49982 31726 50034 31778
rect 54126 31726 54178 31778
rect 55358 31726 55410 31778
rect 56142 31726 56194 31778
rect 59502 31726 59554 31778
rect 60286 31726 60338 31778
rect 61518 31726 61570 31778
rect 61854 31726 61906 31778
rect 63310 31726 63362 31778
rect 69806 31726 69858 31778
rect 70814 31726 70866 31778
rect 76190 31726 76242 31778
rect 1934 31614 1986 31666
rect 3502 31614 3554 31666
rect 4398 31614 4450 31666
rect 6190 31614 6242 31666
rect 15486 31614 15538 31666
rect 15710 31614 15762 31666
rect 24558 31614 24610 31666
rect 46846 31614 46898 31666
rect 47294 31614 47346 31666
rect 51102 31614 51154 31666
rect 52222 31614 52274 31666
rect 53790 31614 53842 31666
rect 54910 31614 54962 31666
rect 56814 31614 56866 31666
rect 59726 31614 59778 31666
rect 60398 31614 60450 31666
rect 62526 31614 62578 31666
rect 65998 31614 66050 31666
rect 66782 31614 66834 31666
rect 69582 31614 69634 31666
rect 71262 31614 71314 31666
rect 72046 31614 72098 31666
rect 73502 31614 73554 31666
rect 74398 31614 74450 31666
rect 77422 31614 77474 31666
rect 6078 31502 6130 31554
rect 6302 31502 6354 31554
rect 11902 31502 11954 31554
rect 15598 31502 15650 31554
rect 16158 31502 16210 31554
rect 24670 31502 24722 31554
rect 25342 31502 25394 31554
rect 30606 31502 30658 31554
rect 39006 31502 39058 31554
rect 46622 31502 46674 31554
rect 47518 31502 47570 31554
rect 48078 31502 48130 31554
rect 50318 31502 50370 31554
rect 51214 31502 51266 31554
rect 51438 31502 51490 31554
rect 51774 31502 51826 31554
rect 53902 31502 53954 31554
rect 57262 31502 57314 31554
rect 57710 31502 57762 31554
rect 58270 31502 58322 31554
rect 61854 31502 61906 31554
rect 62638 31502 62690 31554
rect 63646 31502 63698 31554
rect 63870 31502 63922 31554
rect 64318 31502 64370 31554
rect 65774 31502 65826 31554
rect 66670 31502 66722 31554
rect 67230 31502 67282 31554
rect 68574 31502 68626 31554
rect 71934 31502 71986 31554
rect 73390 31502 73442 31554
rect 74174 31502 74226 31554
rect 77534 31502 77586 31554
rect 20534 31334 20586 31386
rect 20638 31334 20690 31386
rect 20742 31334 20794 31386
rect 39854 31334 39906 31386
rect 39958 31334 40010 31386
rect 40062 31334 40114 31386
rect 59174 31334 59226 31386
rect 59278 31334 59330 31386
rect 59382 31334 59434 31386
rect 78494 31334 78546 31386
rect 78598 31334 78650 31386
rect 78702 31334 78754 31386
rect 8878 31166 8930 31218
rect 13470 31166 13522 31218
rect 13694 31166 13746 31218
rect 14702 31166 14754 31218
rect 14814 31166 14866 31218
rect 14926 31166 14978 31218
rect 18622 31166 18674 31218
rect 27694 31166 27746 31218
rect 31726 31166 31778 31218
rect 44158 31166 44210 31218
rect 46510 31166 46562 31218
rect 48414 31166 48466 31218
rect 54350 31166 54402 31218
rect 58494 31166 58546 31218
rect 65550 31166 65602 31218
rect 67342 31166 67394 31218
rect 68238 31166 68290 31218
rect 69582 31166 69634 31218
rect 71822 31166 71874 31218
rect 71934 31166 71986 31218
rect 72270 31166 72322 31218
rect 74622 31166 74674 31218
rect 2718 31054 2770 31106
rect 3054 31054 3106 31106
rect 5966 31054 6018 31106
rect 7086 31054 7138 31106
rect 8206 31054 8258 31106
rect 16942 31054 16994 31106
rect 20638 31054 20690 31106
rect 24334 31054 24386 31106
rect 26686 31054 26738 31106
rect 27806 31054 27858 31106
rect 31166 31054 31218 31106
rect 35534 31054 35586 31106
rect 37102 31054 37154 31106
rect 42030 31054 42082 31106
rect 43598 31054 43650 31106
rect 50430 31054 50482 31106
rect 55358 31054 55410 31106
rect 58606 31054 58658 31106
rect 60734 31054 60786 31106
rect 65998 31054 66050 31106
rect 66894 31054 66946 31106
rect 68462 31054 68514 31106
rect 70254 31054 70306 31106
rect 74846 31054 74898 31106
rect 76862 31054 76914 31106
rect 4174 30942 4226 30994
rect 4510 30942 4562 30994
rect 5182 30942 5234 30994
rect 6638 30942 6690 30994
rect 6862 30942 6914 30994
rect 6974 30942 7026 30994
rect 9774 30942 9826 30994
rect 10446 30942 10498 30994
rect 13806 30942 13858 30994
rect 15374 30942 15426 30994
rect 16046 30942 16098 30994
rect 18510 30942 18562 30994
rect 18734 30942 18786 30994
rect 19182 30942 19234 30994
rect 19966 30942 20018 30994
rect 23886 30942 23938 30994
rect 26014 30942 26066 30994
rect 27246 30942 27298 30994
rect 27470 30942 27522 30994
rect 30494 30942 30546 30994
rect 31054 30942 31106 30994
rect 36430 30942 36482 30994
rect 39342 30942 39394 30994
rect 40462 30942 40514 30994
rect 40798 30942 40850 30994
rect 41582 30942 41634 30994
rect 41806 30942 41858 30994
rect 42142 30942 42194 30994
rect 43822 30942 43874 30994
rect 48750 30942 48802 30994
rect 50318 30942 50370 30994
rect 51550 30942 51602 30994
rect 51886 30942 51938 30994
rect 54238 30942 54290 30994
rect 54462 30942 54514 30994
rect 54910 30942 54962 30994
rect 61070 30942 61122 30994
rect 61630 30942 61682 30994
rect 63198 30942 63250 30994
rect 66110 30942 66162 30994
rect 66334 30942 66386 30994
rect 67118 30942 67170 30994
rect 67566 30942 67618 30994
rect 68574 30942 68626 30994
rect 69134 30942 69186 30994
rect 69470 30942 69522 30994
rect 69694 30942 69746 30994
rect 70702 30942 70754 30994
rect 72046 30942 72098 30994
rect 74958 30942 75010 30994
rect 75966 30942 76018 30994
rect 76078 30942 76130 30994
rect 76190 30942 76242 30994
rect 77086 30942 77138 30994
rect 77646 30942 77698 30994
rect 8990 30830 9042 30882
rect 10110 30830 10162 30882
rect 10334 30830 10386 30882
rect 16718 30830 16770 30882
rect 17614 30830 17666 30882
rect 19742 30830 19794 30882
rect 22878 30830 22930 30882
rect 23438 30830 23490 30882
rect 24894 30830 24946 30882
rect 25902 30830 25954 30882
rect 29598 30830 29650 30882
rect 32286 30830 32338 30882
rect 32734 30830 32786 30882
rect 33854 30830 33906 30882
rect 34414 30830 34466 30882
rect 34974 30830 35026 30882
rect 39118 30830 39170 30882
rect 39678 30830 39730 30882
rect 40238 30830 40290 30882
rect 45390 30830 45442 30882
rect 45950 30830 46002 30882
rect 46174 30830 46226 30882
rect 50990 30830 51042 30882
rect 52446 30830 52498 30882
rect 53566 30830 53618 30882
rect 54686 30830 54738 30882
rect 55806 30830 55858 30882
rect 56254 30830 56306 30882
rect 59726 30830 59778 30882
rect 60174 30830 60226 30882
rect 61966 30830 62018 30882
rect 63870 30830 63922 30882
rect 71150 30830 71202 30882
rect 75518 30830 75570 30882
rect 8654 30718 8706 30770
rect 32062 30718 32114 30770
rect 58382 30718 58434 30770
rect 62190 30718 62242 30770
rect 63310 30718 63362 30770
rect 10874 30550 10926 30602
rect 10978 30550 11030 30602
rect 11082 30550 11134 30602
rect 30194 30550 30246 30602
rect 30298 30550 30350 30602
rect 30402 30550 30454 30602
rect 49514 30550 49566 30602
rect 49618 30550 49670 30602
rect 49722 30550 49774 30602
rect 68834 30550 68886 30602
rect 68938 30550 68990 30602
rect 69042 30550 69094 30602
rect 4174 30382 4226 30434
rect 19182 30382 19234 30434
rect 54798 30382 54850 30434
rect 55582 30382 55634 30434
rect 57486 30382 57538 30434
rect 70142 30382 70194 30434
rect 70702 30382 70754 30434
rect 71038 30382 71090 30434
rect 71710 30382 71762 30434
rect 76414 30382 76466 30434
rect 76750 30382 76802 30434
rect 11566 30270 11618 30322
rect 16606 30270 16658 30322
rect 19294 30270 19346 30322
rect 23998 30270 24050 30322
rect 26014 30270 26066 30322
rect 30942 30270 30994 30322
rect 33854 30270 33906 30322
rect 34750 30270 34802 30322
rect 35422 30270 35474 30322
rect 44718 30270 44770 30322
rect 47854 30270 47906 30322
rect 48302 30270 48354 30322
rect 49758 30270 49810 30322
rect 50542 30270 50594 30322
rect 57150 30270 57202 30322
rect 58382 30270 58434 30322
rect 61406 30270 61458 30322
rect 61742 30270 61794 30322
rect 67006 30270 67058 30322
rect 72270 30270 72322 30322
rect 74398 30270 74450 30322
rect 74510 30270 74562 30322
rect 75406 30270 75458 30322
rect 4062 30158 4114 30210
rect 6750 30158 6802 30210
rect 6974 30158 7026 30210
rect 7646 30158 7698 30210
rect 9438 30158 9490 30210
rect 9774 30158 9826 30210
rect 10334 30158 10386 30210
rect 10558 30158 10610 30210
rect 11006 30158 11058 30210
rect 11790 30158 11842 30210
rect 12462 30158 12514 30210
rect 14030 30158 14082 30210
rect 14366 30158 14418 30210
rect 14814 30158 14866 30210
rect 15038 30158 15090 30210
rect 15822 30158 15874 30210
rect 16158 30158 16210 30210
rect 18958 30158 19010 30210
rect 23886 30158 23938 30210
rect 25790 30158 25842 30210
rect 26350 30158 26402 30210
rect 30046 30158 30098 30210
rect 30270 30158 30322 30210
rect 31502 30158 31554 30210
rect 31838 30158 31890 30210
rect 35310 30158 35362 30210
rect 35982 30158 36034 30210
rect 36318 30158 36370 30210
rect 36654 30158 36706 30210
rect 37438 30158 37490 30210
rect 46062 30158 46114 30210
rect 46958 30158 47010 30210
rect 50430 30158 50482 30210
rect 53902 30158 53954 30210
rect 54238 30158 54290 30210
rect 58494 30158 58546 30210
rect 62078 30158 62130 30210
rect 66110 30158 66162 30210
rect 66782 30158 66834 30210
rect 67566 30158 67618 30210
rect 72046 30158 72098 30210
rect 75070 30158 75122 30210
rect 75518 30158 75570 30210
rect 77310 30158 77362 30210
rect 3166 30046 3218 30098
rect 9550 30046 9602 30098
rect 10446 30046 10498 30098
rect 23550 30046 23602 30098
rect 24110 30046 24162 30098
rect 31614 30046 31666 30098
rect 32174 30046 32226 30098
rect 32734 30046 32786 30098
rect 34414 30046 34466 30098
rect 41694 30046 41746 30098
rect 44382 30046 44434 30098
rect 47182 30046 47234 30098
rect 47742 30046 47794 30098
rect 54686 30046 54738 30098
rect 55694 30046 55746 30098
rect 58158 30046 58210 30098
rect 67790 30046 67842 30098
rect 67902 30046 67954 30098
rect 68462 30046 68514 30098
rect 68574 30046 68626 30098
rect 69470 30046 69522 30098
rect 69582 30046 69634 30098
rect 69694 30046 69746 30098
rect 77534 30046 77586 30098
rect 77758 30046 77810 30098
rect 77870 30046 77922 30098
rect 2382 29934 2434 29986
rect 2830 29934 2882 29986
rect 4174 29934 4226 29986
rect 4846 29934 4898 29986
rect 12910 29934 12962 29986
rect 14142 29934 14194 29986
rect 15374 29934 15426 29986
rect 16046 29934 16098 29986
rect 17166 29934 17218 29986
rect 22990 29934 23042 29986
rect 24894 29934 24946 29986
rect 25230 29934 25282 29986
rect 26910 29934 26962 29986
rect 27358 29934 27410 29986
rect 28142 29934 28194 29986
rect 28814 29934 28866 29986
rect 32846 29934 32898 29986
rect 33070 29934 33122 29986
rect 33406 29934 33458 29986
rect 34638 29934 34690 29986
rect 35534 29934 35586 29986
rect 36542 29934 36594 29986
rect 41358 29934 41410 29986
rect 43822 29934 43874 29986
rect 44606 29934 44658 29986
rect 46286 29934 46338 29986
rect 53454 29934 53506 29986
rect 54014 29934 54066 29986
rect 54798 29934 54850 29986
rect 55582 29934 55634 29986
rect 56254 29934 56306 29986
rect 56702 29934 56754 29986
rect 57374 29934 57426 29986
rect 60622 29934 60674 29986
rect 70814 29934 70866 29986
rect 72718 29934 72770 29986
rect 74286 29934 74338 29986
rect 76638 29934 76690 29986
rect 20534 29766 20586 29818
rect 20638 29766 20690 29818
rect 20742 29766 20794 29818
rect 39854 29766 39906 29818
rect 39958 29766 40010 29818
rect 40062 29766 40114 29818
rect 59174 29766 59226 29818
rect 59278 29766 59330 29818
rect 59382 29766 59434 29818
rect 78494 29766 78546 29818
rect 78598 29766 78650 29818
rect 78702 29766 78754 29818
rect 9886 29598 9938 29650
rect 12126 29598 12178 29650
rect 13918 29598 13970 29650
rect 16382 29598 16434 29650
rect 19518 29598 19570 29650
rect 28590 29598 28642 29650
rect 28814 29598 28866 29650
rect 29822 29598 29874 29650
rect 33966 29598 34018 29650
rect 36094 29598 36146 29650
rect 40462 29598 40514 29650
rect 51102 29598 51154 29650
rect 60734 29598 60786 29650
rect 63646 29598 63698 29650
rect 70702 29598 70754 29650
rect 71710 29598 71762 29650
rect 4622 29486 4674 29538
rect 6526 29486 6578 29538
rect 12350 29486 12402 29538
rect 15486 29486 15538 29538
rect 18286 29486 18338 29538
rect 21310 29486 21362 29538
rect 23998 29486 24050 29538
rect 26910 29486 26962 29538
rect 33630 29486 33682 29538
rect 33742 29486 33794 29538
rect 37886 29486 37938 29538
rect 43710 29486 43762 29538
rect 45950 29486 46002 29538
rect 46510 29486 46562 29538
rect 51326 29486 51378 29538
rect 53006 29486 53058 29538
rect 54910 29486 54962 29538
rect 59726 29486 59778 29538
rect 59838 29486 59890 29538
rect 63870 29486 63922 29538
rect 67790 29486 67842 29538
rect 68238 29486 68290 29538
rect 71486 29486 71538 29538
rect 2830 29374 2882 29426
rect 4174 29374 4226 29426
rect 4510 29374 4562 29426
rect 7198 29374 7250 29426
rect 11454 29374 11506 29426
rect 12462 29374 12514 29426
rect 14814 29374 14866 29426
rect 18062 29374 18114 29426
rect 18398 29374 18450 29426
rect 22430 29374 22482 29426
rect 23102 29374 23154 29426
rect 23662 29374 23714 29426
rect 27358 29374 27410 29426
rect 27806 29374 27858 29426
rect 28478 29374 28530 29426
rect 32398 29374 32450 29426
rect 37326 29374 37378 29426
rect 40126 29374 40178 29426
rect 40574 29374 40626 29426
rect 40686 29374 40738 29426
rect 41806 29374 41858 29426
rect 43150 29374 43202 29426
rect 45278 29374 45330 29426
rect 46846 29374 46898 29426
rect 49646 29374 49698 29426
rect 50206 29374 50258 29426
rect 51438 29374 51490 29426
rect 54574 29374 54626 29426
rect 54686 29374 54738 29426
rect 55134 29374 55186 29426
rect 56254 29374 56306 29426
rect 58606 29374 58658 29426
rect 59502 29374 59554 29426
rect 63982 29374 64034 29426
rect 64542 29374 64594 29426
rect 70814 29374 70866 29426
rect 71374 29374 71426 29426
rect 75182 29374 75234 29426
rect 1934 29262 1986 29314
rect 5070 29262 5122 29314
rect 6862 29262 6914 29314
rect 7982 29262 8034 29314
rect 10670 29262 10722 29314
rect 11342 29262 11394 29314
rect 12910 29262 12962 29314
rect 13358 29262 13410 29314
rect 15038 29262 15090 29314
rect 18958 29262 19010 29314
rect 21198 29262 21250 29314
rect 21534 29262 21586 29314
rect 22206 29262 22258 29314
rect 24558 29262 24610 29314
rect 25902 29262 25954 29314
rect 26350 29262 26402 29314
rect 29374 29262 29426 29314
rect 32062 29262 32114 29314
rect 32734 29262 32786 29314
rect 37102 29262 37154 29314
rect 38558 29262 38610 29314
rect 39118 29262 39170 29314
rect 39678 29262 39730 29314
rect 41694 29262 41746 29314
rect 44382 29262 44434 29314
rect 45054 29262 45106 29314
rect 48190 29262 48242 29314
rect 50430 29262 50482 29314
rect 55918 29262 55970 29314
rect 56590 29262 56642 29314
rect 58158 29262 58210 29314
rect 60286 29262 60338 29314
rect 64654 29262 64706 29314
rect 67342 29262 67394 29314
rect 68798 29262 68850 29314
rect 70030 29262 70082 29314
rect 72046 29262 72098 29314
rect 76078 29262 76130 29314
rect 76750 29262 76802 29314
rect 77086 29262 77138 29314
rect 77646 29262 77698 29314
rect 77982 29262 78034 29314
rect 19182 29150 19234 29202
rect 39342 29150 39394 29202
rect 48414 29150 48466 29202
rect 48750 29150 48802 29202
rect 52782 29150 52834 29202
rect 53118 29150 53170 29202
rect 58942 29150 58994 29202
rect 70702 29150 70754 29202
rect 76638 29150 76690 29202
rect 77646 29150 77698 29202
rect 10874 28982 10926 29034
rect 10978 28982 11030 29034
rect 11082 28982 11134 29034
rect 30194 28982 30246 29034
rect 30298 28982 30350 29034
rect 30402 28982 30454 29034
rect 49514 28982 49566 29034
rect 49618 28982 49670 29034
rect 49722 28982 49774 29034
rect 68834 28982 68886 29034
rect 68938 28982 68990 29034
rect 69042 28982 69094 29034
rect 6750 28814 6802 28866
rect 10670 28814 10722 28866
rect 14254 28814 14306 28866
rect 28814 28814 28866 28866
rect 33742 28814 33794 28866
rect 40574 28814 40626 28866
rect 40910 28814 40962 28866
rect 69470 28814 69522 28866
rect 77310 28814 77362 28866
rect 3614 28702 3666 28754
rect 4958 28702 5010 28754
rect 10446 28702 10498 28754
rect 14814 28702 14866 28754
rect 17838 28702 17890 28754
rect 18622 28702 18674 28754
rect 20862 28702 20914 28754
rect 22878 28702 22930 28754
rect 24782 28702 24834 28754
rect 27022 28702 27074 28754
rect 30606 28702 30658 28754
rect 32062 28702 32114 28754
rect 32398 28702 32450 28754
rect 40014 28702 40066 28754
rect 41134 28702 41186 28754
rect 46398 28702 46450 28754
rect 52334 28702 52386 28754
rect 65102 28702 65154 28754
rect 65774 28702 65826 28754
rect 71486 28702 71538 28754
rect 73838 28702 73890 28754
rect 74622 28702 74674 28754
rect 76190 28702 76242 28754
rect 77870 28702 77922 28754
rect 7086 28590 7138 28642
rect 7310 28590 7362 28642
rect 7758 28590 7810 28642
rect 10334 28590 10386 28642
rect 12126 28590 12178 28642
rect 12574 28590 12626 28642
rect 14590 28590 14642 28642
rect 15374 28590 15426 28642
rect 17726 28590 17778 28642
rect 18846 28590 18898 28642
rect 20190 28590 20242 28642
rect 23998 28590 24050 28642
rect 24446 28590 24498 28642
rect 25566 28590 25618 28642
rect 26462 28590 26514 28642
rect 28478 28590 28530 28642
rect 29710 28590 29762 28642
rect 29934 28590 29986 28642
rect 31614 28590 31666 28642
rect 32510 28590 32562 28642
rect 34302 28590 34354 28642
rect 36878 28590 36930 28642
rect 37438 28590 37490 28642
rect 46622 28590 46674 28642
rect 48302 28590 48354 28642
rect 48638 28590 48690 28642
rect 49870 28590 49922 28642
rect 50318 28590 50370 28642
rect 54014 28590 54066 28642
rect 56030 28590 56082 28642
rect 58830 28590 58882 28642
rect 59726 28590 59778 28642
rect 60174 28590 60226 28642
rect 61966 28590 62018 28642
rect 64206 28590 64258 28642
rect 64654 28590 64706 28642
rect 65998 28590 66050 28642
rect 67342 28590 67394 28642
rect 67566 28590 67618 28642
rect 71038 28590 71090 28642
rect 71934 28590 71986 28642
rect 74510 28590 74562 28642
rect 75406 28590 75458 28642
rect 76302 28590 76354 28642
rect 77646 28590 77698 28642
rect 2830 28478 2882 28530
rect 3166 28478 3218 28530
rect 4622 28478 4674 28530
rect 13806 28478 13858 28530
rect 17390 28478 17442 28530
rect 17950 28478 18002 28530
rect 25902 28478 25954 28530
rect 27582 28478 27634 28530
rect 28702 28478 28754 28530
rect 33630 28478 33682 28530
rect 33742 28478 33794 28530
rect 36542 28478 36594 28530
rect 37998 28478 38050 28530
rect 47294 28478 47346 28530
rect 48414 28478 48466 28530
rect 50430 28478 50482 28530
rect 50542 28478 50594 28530
rect 53454 28478 53506 28530
rect 54574 28478 54626 28530
rect 54798 28478 54850 28530
rect 55246 28478 55298 28530
rect 55582 28478 55634 28530
rect 58158 28478 58210 28530
rect 60622 28478 60674 28530
rect 61406 28478 61458 28530
rect 61518 28478 61570 28530
rect 66670 28478 66722 28530
rect 68238 28478 68290 28530
rect 69470 28478 69522 28530
rect 69582 28478 69634 28530
rect 4846 28366 4898 28418
rect 5630 28366 5682 28418
rect 16942 28366 16994 28418
rect 22430 28366 22482 28418
rect 22990 28366 23042 28418
rect 23438 28366 23490 28418
rect 25790 28366 25842 28418
rect 26798 28366 26850 28418
rect 27022 28366 27074 28418
rect 27694 28366 27746 28418
rect 27918 28366 27970 28418
rect 31166 28366 31218 28418
rect 35646 28366 35698 28418
rect 36094 28366 36146 28418
rect 36654 28366 36706 28418
rect 37886 28366 37938 28418
rect 38110 28366 38162 28418
rect 52446 28366 52498 28418
rect 53678 28366 53730 28418
rect 53902 28366 53954 28418
rect 54686 28366 54738 28418
rect 55470 28366 55522 28418
rect 58270 28366 58322 28418
rect 58494 28366 58546 28418
rect 61630 28366 61682 28418
rect 20534 28198 20586 28250
rect 20638 28198 20690 28250
rect 20742 28198 20794 28250
rect 39854 28198 39906 28250
rect 39958 28198 40010 28250
rect 40062 28198 40114 28250
rect 59174 28198 59226 28250
rect 59278 28198 59330 28250
rect 59382 28198 59434 28250
rect 78494 28198 78546 28250
rect 78598 28198 78650 28250
rect 78702 28198 78754 28250
rect 5294 28030 5346 28082
rect 5406 28030 5458 28082
rect 6526 28030 6578 28082
rect 13918 28030 13970 28082
rect 14702 28030 14754 28082
rect 18286 28030 18338 28082
rect 19070 28030 19122 28082
rect 23662 28030 23714 28082
rect 24894 28030 24946 28082
rect 28702 28030 28754 28082
rect 42142 28030 42194 28082
rect 56814 28030 56866 28082
rect 61966 28030 62018 28082
rect 65438 28030 65490 28082
rect 71486 28030 71538 28082
rect 75070 28030 75122 28082
rect 76526 28030 76578 28082
rect 3166 27918 3218 27970
rect 4734 27918 4786 27970
rect 8766 27918 8818 27970
rect 13358 27918 13410 27970
rect 14142 27918 14194 27970
rect 14926 27918 14978 27970
rect 19182 27918 19234 27970
rect 22430 27918 22482 27970
rect 26798 27918 26850 27970
rect 28142 27918 28194 27970
rect 28590 27918 28642 27970
rect 30718 27918 30770 27970
rect 37214 27918 37266 27970
rect 40798 27918 40850 27970
rect 46286 27918 46338 27970
rect 53790 27918 53842 27970
rect 54574 27918 54626 27970
rect 56590 27918 56642 27970
rect 59278 27918 59330 27970
rect 61406 27918 61458 27970
rect 61854 27918 61906 27970
rect 62862 27918 62914 27970
rect 65998 27918 66050 27970
rect 70030 27918 70082 27970
rect 71374 27918 71426 27970
rect 71598 27918 71650 27970
rect 75518 27918 75570 27970
rect 75742 27918 75794 27970
rect 76750 27918 76802 27970
rect 77758 27918 77810 27970
rect 3390 27806 3442 27858
rect 4286 27806 4338 27858
rect 5518 27806 5570 27858
rect 5966 27806 6018 27858
rect 6302 27806 6354 27858
rect 6638 27806 6690 27858
rect 8318 27806 8370 27858
rect 11006 27806 11058 27858
rect 13246 27806 13298 27858
rect 13582 27806 13634 27858
rect 14254 27806 14306 27858
rect 15038 27806 15090 27858
rect 18846 27806 18898 27858
rect 21870 27806 21922 27858
rect 22654 27806 22706 27858
rect 22878 27806 22930 27858
rect 26574 27806 26626 27858
rect 27358 27806 27410 27858
rect 28030 27806 28082 27858
rect 28926 27806 28978 27858
rect 29038 27806 29090 27858
rect 30046 27806 30098 27858
rect 30830 27806 30882 27858
rect 31614 27806 31666 27858
rect 36318 27806 36370 27858
rect 40126 27806 40178 27858
rect 45054 27806 45106 27858
rect 45278 27806 45330 27858
rect 46062 27806 46114 27858
rect 46622 27806 46674 27858
rect 49870 27806 49922 27858
rect 52558 27806 52610 27858
rect 52894 27806 52946 27858
rect 53566 27806 53618 27858
rect 54350 27806 54402 27858
rect 54686 27806 54738 27858
rect 56478 27806 56530 27858
rect 58494 27806 58546 27858
rect 60398 27806 60450 27858
rect 61630 27806 61682 27858
rect 62750 27806 62802 27858
rect 63086 27806 63138 27858
rect 65774 27806 65826 27858
rect 69470 27806 69522 27858
rect 75630 27806 75682 27858
rect 76414 27806 76466 27858
rect 76974 27806 77026 27858
rect 7086 27694 7138 27746
rect 7870 27694 7922 27746
rect 10446 27694 10498 27746
rect 11118 27694 11170 27746
rect 12014 27694 12066 27746
rect 12686 27694 12738 27746
rect 15598 27694 15650 27746
rect 15934 27694 15986 27746
rect 16494 27694 16546 27746
rect 17054 27694 17106 27746
rect 17726 27694 17778 27746
rect 19742 27694 19794 27746
rect 20078 27694 20130 27746
rect 20526 27694 20578 27746
rect 21086 27694 21138 27746
rect 21422 27694 21474 27746
rect 22766 27694 22818 27746
rect 24222 27694 24274 27746
rect 25566 27694 25618 27746
rect 26014 27694 26066 27746
rect 32062 27694 32114 27746
rect 32398 27694 32450 27746
rect 35086 27694 35138 27746
rect 35534 27694 35586 27746
rect 36430 27694 36482 27746
rect 39342 27694 39394 27746
rect 39902 27694 39954 27746
rect 41582 27694 41634 27746
rect 45390 27694 45442 27746
rect 46510 27694 46562 27746
rect 49758 27694 49810 27746
rect 55918 27694 55970 27746
rect 57374 27694 57426 27746
rect 59390 27694 59442 27746
rect 59838 27694 59890 27746
rect 60846 27694 60898 27746
rect 69582 27694 69634 27746
rect 72046 27694 72098 27746
rect 74174 27694 74226 27746
rect 74510 27694 74562 27746
rect 77870 27694 77922 27746
rect 17950 27582 18002 27634
rect 23438 27582 23490 27634
rect 23774 27582 23826 27634
rect 30718 27582 30770 27634
rect 41806 27582 41858 27634
rect 50206 27582 50258 27634
rect 52670 27582 52722 27634
rect 55134 27582 55186 27634
rect 58158 27582 58210 27634
rect 58494 27582 58546 27634
rect 59054 27582 59106 27634
rect 60622 27582 60674 27634
rect 60846 27582 60898 27634
rect 61182 27582 61234 27634
rect 77534 27582 77586 27634
rect 10874 27414 10926 27466
rect 10978 27414 11030 27466
rect 11082 27414 11134 27466
rect 30194 27414 30246 27466
rect 30298 27414 30350 27466
rect 30402 27414 30454 27466
rect 49514 27414 49566 27466
rect 49618 27414 49670 27466
rect 49722 27414 49774 27466
rect 68834 27414 68886 27466
rect 68938 27414 68990 27466
rect 69042 27414 69094 27466
rect 10110 27246 10162 27298
rect 16942 27246 16994 27298
rect 17390 27246 17442 27298
rect 17726 27246 17778 27298
rect 18958 27246 19010 27298
rect 28366 27246 28418 27298
rect 36318 27246 36370 27298
rect 39678 27246 39730 27298
rect 45950 27246 46002 27298
rect 48078 27246 48130 27298
rect 48302 27246 48354 27298
rect 48750 27246 48802 27298
rect 54574 27246 54626 27298
rect 54910 27246 54962 27298
rect 56142 27246 56194 27298
rect 56478 27246 56530 27298
rect 57598 27246 57650 27298
rect 62974 27246 63026 27298
rect 63982 27246 64034 27298
rect 65998 27246 66050 27298
rect 66334 27246 66386 27298
rect 73054 27246 73106 27298
rect 76414 27246 76466 27298
rect 77310 27246 77362 27298
rect 4174 27134 4226 27186
rect 4958 27134 5010 27186
rect 5854 27134 5906 27186
rect 8878 27134 8930 27186
rect 9550 27134 9602 27186
rect 23102 27134 23154 27186
rect 28254 27134 28306 27186
rect 30942 27134 30994 27186
rect 31838 27134 31890 27186
rect 34638 27134 34690 27186
rect 35646 27134 35698 27186
rect 39230 27134 39282 27186
rect 42142 27134 42194 27186
rect 44718 27134 44770 27186
rect 57038 27134 57090 27186
rect 58270 27134 58322 27186
rect 74846 27134 74898 27186
rect 78094 27134 78146 27186
rect 3726 27022 3778 27074
rect 4062 27022 4114 27074
rect 5742 27022 5794 27074
rect 6078 27022 6130 27074
rect 10446 27022 10498 27074
rect 10558 27022 10610 27074
rect 11342 27022 11394 27074
rect 14030 27022 14082 27074
rect 14814 27022 14866 27074
rect 17502 27022 17554 27074
rect 19070 27022 19122 27074
rect 19966 27022 20018 27074
rect 23214 27022 23266 27074
rect 23886 27022 23938 27074
rect 24334 27022 24386 27074
rect 25230 27022 25282 27074
rect 26574 27022 26626 27074
rect 27694 27022 27746 27074
rect 32062 27022 32114 27074
rect 34302 27022 34354 27074
rect 34862 27022 34914 27074
rect 35982 27022 36034 27074
rect 38558 27022 38610 27074
rect 39790 27022 39842 27074
rect 40574 27022 40626 27074
rect 41246 27022 41298 27074
rect 44046 27022 44098 27074
rect 44606 27022 44658 27074
rect 45502 27022 45554 27074
rect 45726 27022 45778 27074
rect 46062 27022 46114 27074
rect 48526 27022 48578 27074
rect 48974 27022 49026 27074
rect 49422 27022 49474 27074
rect 53902 27022 53954 27074
rect 57262 27022 57314 27074
rect 58606 27022 58658 27074
rect 63870 27022 63922 27074
rect 64878 27022 64930 27074
rect 68350 27022 68402 27074
rect 69470 27022 69522 27074
rect 69918 27022 69970 27074
rect 71038 27022 71090 27074
rect 71262 27022 71314 27074
rect 71934 27022 71986 27074
rect 72494 27022 72546 27074
rect 72718 27022 72770 27074
rect 75630 27022 75682 27074
rect 77310 27022 77362 27074
rect 8654 26910 8706 26962
rect 8878 26910 8930 26962
rect 9102 26910 9154 26962
rect 10670 26910 10722 26962
rect 11678 26910 11730 26962
rect 13694 26910 13746 26962
rect 14366 26910 14418 26962
rect 15150 26910 15202 26962
rect 16158 26910 16210 26962
rect 16718 26910 16770 26962
rect 17054 26910 17106 26962
rect 18062 26910 18114 26962
rect 20750 26910 20802 26962
rect 22542 26910 22594 26962
rect 22766 26910 22818 26962
rect 24782 26910 24834 26962
rect 26686 26910 26738 26962
rect 27358 26910 27410 26962
rect 28814 26910 28866 26962
rect 31502 26910 31554 26962
rect 31726 26910 31778 26962
rect 32398 26910 32450 26962
rect 34414 26910 34466 26962
rect 39902 26910 39954 26962
rect 52670 26910 52722 26962
rect 54686 26910 54738 26962
rect 56366 26910 56418 26962
rect 59166 26910 59218 26962
rect 61630 26910 61682 26962
rect 63310 26910 63362 26962
rect 65214 26910 65266 26962
rect 65774 26910 65826 26962
rect 70366 26910 70418 26962
rect 74174 26910 74226 26962
rect 74734 26910 74786 26962
rect 75854 26910 75906 26962
rect 75966 26910 76018 26962
rect 77646 26910 77698 26962
rect 7086 26798 7138 26850
rect 8206 26798 8258 26850
rect 10782 26798 10834 26850
rect 11566 26798 11618 26850
rect 12462 26798 12514 26850
rect 12910 26798 12962 26850
rect 14254 26798 14306 26850
rect 15038 26798 15090 26850
rect 15598 26798 15650 26850
rect 18174 26798 18226 26850
rect 18398 26798 18450 26850
rect 18958 26798 19010 26850
rect 19630 26798 19682 26850
rect 19854 26798 19906 26850
rect 21534 26798 21586 26850
rect 21982 26798 22034 26850
rect 22990 26798 23042 26850
rect 26014 26798 26066 26850
rect 26910 26798 26962 26850
rect 27470 26798 27522 26850
rect 33742 26798 33794 26850
rect 39118 26798 39170 26850
rect 41694 26798 41746 26850
rect 46286 26798 46338 26850
rect 49422 26798 49474 26850
rect 52334 26798 52386 26850
rect 53566 26798 53618 26850
rect 53790 26798 53842 26850
rect 54014 26798 54066 26850
rect 61742 26798 61794 26850
rect 61966 26798 62018 26850
rect 63086 26798 63138 26850
rect 63982 26798 64034 26850
rect 65102 26798 65154 26850
rect 68462 26798 68514 26850
rect 68686 26798 68738 26850
rect 74958 26798 75010 26850
rect 20534 26630 20586 26682
rect 20638 26630 20690 26682
rect 20742 26630 20794 26682
rect 39854 26630 39906 26682
rect 39958 26630 40010 26682
rect 40062 26630 40114 26682
rect 59174 26630 59226 26682
rect 59278 26630 59330 26682
rect 59382 26630 59434 26682
rect 78494 26630 78546 26682
rect 78598 26630 78650 26682
rect 78702 26630 78754 26682
rect 5406 26462 5458 26514
rect 6190 26462 6242 26514
rect 6302 26462 6354 26514
rect 7646 26462 7698 26514
rect 8654 26462 8706 26514
rect 10446 26462 10498 26514
rect 12910 26462 12962 26514
rect 13582 26462 13634 26514
rect 13806 26462 13858 26514
rect 19630 26462 19682 26514
rect 22990 26462 23042 26514
rect 24558 26462 24610 26514
rect 25566 26462 25618 26514
rect 36542 26462 36594 26514
rect 43150 26462 43202 26514
rect 45054 26462 45106 26514
rect 45502 26462 45554 26514
rect 48750 26462 48802 26514
rect 49646 26462 49698 26514
rect 57934 26462 57986 26514
rect 65438 26462 65490 26514
rect 69694 26462 69746 26514
rect 69806 26462 69858 26514
rect 70478 26462 70530 26514
rect 74286 26462 74338 26514
rect 6526 26350 6578 26402
rect 7422 26350 7474 26402
rect 7982 26350 8034 26402
rect 8878 26350 8930 26402
rect 12014 26350 12066 26402
rect 13694 26350 13746 26402
rect 16718 26350 16770 26402
rect 16830 26350 16882 26402
rect 18398 26350 18450 26402
rect 20638 26350 20690 26402
rect 28366 26350 28418 26402
rect 31390 26350 31442 26402
rect 35422 26350 35474 26402
rect 38670 26350 38722 26402
rect 41918 26350 41970 26402
rect 43822 26350 43874 26402
rect 43934 26350 43986 26402
rect 49758 26350 49810 26402
rect 50430 26350 50482 26402
rect 60062 26350 60114 26402
rect 63758 26350 63810 26402
rect 65550 26350 65602 26402
rect 67006 26350 67058 26402
rect 67902 26350 67954 26402
rect 70366 26350 70418 26402
rect 73838 26350 73890 26402
rect 2830 26238 2882 26290
rect 4062 26238 4114 26290
rect 4510 26238 4562 26290
rect 4846 26238 4898 26290
rect 5294 26238 5346 26290
rect 5518 26238 5570 26290
rect 6078 26238 6130 26290
rect 7310 26238 7362 26290
rect 8990 26238 9042 26290
rect 10334 26238 10386 26290
rect 10558 26238 10610 26290
rect 11006 26238 11058 26290
rect 11454 26238 11506 26290
rect 11790 26238 11842 26290
rect 13918 26238 13970 26290
rect 14142 26238 14194 26290
rect 14814 26238 14866 26290
rect 15262 26238 15314 26290
rect 17054 26238 17106 26290
rect 19518 26238 19570 26290
rect 20750 26238 20802 26290
rect 23550 26238 23602 26290
rect 27470 26238 27522 26290
rect 27694 26238 27746 26290
rect 29822 26238 29874 26290
rect 30942 26238 30994 26290
rect 31950 26238 32002 26290
rect 32286 26238 32338 26290
rect 32510 26238 32562 26290
rect 34750 26238 34802 26290
rect 36206 26238 36258 26290
rect 38334 26238 38386 26290
rect 39902 26238 39954 26290
rect 41470 26238 41522 26290
rect 42030 26238 42082 26290
rect 42142 26238 42194 26290
rect 44494 26238 44546 26290
rect 50766 26238 50818 26290
rect 52670 26238 52722 26290
rect 53118 26238 53170 26290
rect 53566 26238 53618 26290
rect 57486 26238 57538 26290
rect 57710 26238 57762 26290
rect 58158 26238 58210 26290
rect 61294 26238 61346 26290
rect 61518 26238 61570 26290
rect 62190 26238 62242 26290
rect 62862 26238 62914 26290
rect 63086 26238 63138 26290
rect 69134 26238 69186 26290
rect 69582 26238 69634 26290
rect 71934 26238 71986 26290
rect 72382 26238 72434 26290
rect 74174 26238 74226 26290
rect 74398 26238 74450 26290
rect 76190 26238 76242 26290
rect 77422 26238 77474 26290
rect 1934 26126 1986 26178
rect 3614 26126 3666 26178
rect 9662 26126 9714 26178
rect 11678 26126 11730 26178
rect 12462 26126 12514 26178
rect 15710 26126 15762 26178
rect 16158 26126 16210 26178
rect 17950 26126 18002 26178
rect 21534 26126 21586 26178
rect 21982 26126 22034 26178
rect 22430 26126 22482 26178
rect 24110 26126 24162 26178
rect 29710 26126 29762 26178
rect 30494 26126 30546 26178
rect 32398 26126 32450 26178
rect 33854 26126 33906 26178
rect 34974 26126 35026 26178
rect 35982 26126 36034 26178
rect 39454 26126 39506 26178
rect 40238 26126 40290 26178
rect 48190 26126 48242 26178
rect 56254 26126 56306 26178
rect 56702 26126 56754 26178
rect 57598 26126 57650 26178
rect 58606 26126 58658 26178
rect 59054 26126 59106 26178
rect 60622 26126 60674 26178
rect 64654 26126 64706 26178
rect 65998 26126 66050 26178
rect 68014 26126 68066 26178
rect 75518 26126 75570 26178
rect 77310 26126 77362 26178
rect 77758 26126 77810 26178
rect 3838 26014 3890 26066
rect 20638 26014 20690 26066
rect 21534 26014 21586 26066
rect 21982 26014 22034 26066
rect 38334 26014 38386 26066
rect 43822 26014 43874 26066
rect 44718 26014 44770 26066
rect 48414 26014 48466 26066
rect 49534 26014 49586 26066
rect 66782 26014 66834 26066
rect 67118 26014 67170 26066
rect 67678 26014 67730 26066
rect 72270 26014 72322 26066
rect 10874 25846 10926 25898
rect 10978 25846 11030 25898
rect 11082 25846 11134 25898
rect 30194 25846 30246 25898
rect 30298 25846 30350 25898
rect 30402 25846 30454 25898
rect 49514 25846 49566 25898
rect 49618 25846 49670 25898
rect 49722 25846 49774 25898
rect 68834 25846 68886 25898
rect 68938 25846 68990 25898
rect 69042 25846 69094 25898
rect 18286 25678 18338 25730
rect 23662 25678 23714 25730
rect 27470 25678 27522 25730
rect 57150 25678 57202 25730
rect 66782 25678 66834 25730
rect 72382 25678 72434 25730
rect 77310 25678 77362 25730
rect 3278 25566 3330 25618
rect 4398 25566 4450 25618
rect 6190 25566 6242 25618
rect 7086 25566 7138 25618
rect 7758 25566 7810 25618
rect 10334 25566 10386 25618
rect 14702 25566 14754 25618
rect 15150 25566 15202 25618
rect 19294 25566 19346 25618
rect 25678 25566 25730 25618
rect 27694 25566 27746 25618
rect 28030 25566 28082 25618
rect 34750 25566 34802 25618
rect 38670 25566 38722 25618
rect 39118 25566 39170 25618
rect 39790 25566 39842 25618
rect 40798 25566 40850 25618
rect 43374 25566 43426 25618
rect 53454 25566 53506 25618
rect 54238 25566 54290 25618
rect 58382 25566 58434 25618
rect 61294 25566 61346 25618
rect 62750 25566 62802 25618
rect 64206 25566 64258 25618
rect 64654 25566 64706 25618
rect 66110 25566 66162 25618
rect 67790 25566 67842 25618
rect 69806 25566 69858 25618
rect 76526 25566 76578 25618
rect 77422 25566 77474 25618
rect 77870 25566 77922 25618
rect 3166 25454 3218 25506
rect 3726 25454 3778 25506
rect 4622 25454 4674 25506
rect 6638 25454 6690 25506
rect 7982 25454 8034 25506
rect 10782 25454 10834 25506
rect 17950 25454 18002 25506
rect 18398 25454 18450 25506
rect 19406 25454 19458 25506
rect 20190 25454 20242 25506
rect 21982 25454 22034 25506
rect 23438 25454 23490 25506
rect 27022 25454 27074 25506
rect 27918 25454 27970 25506
rect 33854 25454 33906 25506
rect 34302 25454 34354 25506
rect 39678 25454 39730 25506
rect 39902 25454 39954 25506
rect 40126 25454 40178 25506
rect 43486 25454 43538 25506
rect 43822 25454 43874 25506
rect 45838 25454 45890 25506
rect 53902 25454 53954 25506
rect 57822 25454 57874 25506
rect 58046 25454 58098 25506
rect 59054 25454 59106 25506
rect 62414 25454 62466 25506
rect 62638 25454 62690 25506
rect 62862 25454 62914 25506
rect 63310 25454 63362 25506
rect 65998 25454 66050 25506
rect 67678 25454 67730 25506
rect 69246 25454 69298 25506
rect 75854 25454 75906 25506
rect 76414 25454 76466 25506
rect 4286 25342 4338 25394
rect 7646 25342 7698 25394
rect 11230 25342 11282 25394
rect 20414 25342 20466 25394
rect 20526 25342 20578 25394
rect 21870 25342 21922 25394
rect 22318 25342 22370 25394
rect 23998 25342 24050 25394
rect 24558 25342 24610 25394
rect 24894 25342 24946 25394
rect 26238 25342 26290 25394
rect 26686 25342 26738 25394
rect 26798 25342 26850 25394
rect 33070 25342 33122 25394
rect 33182 25342 33234 25394
rect 40350 25342 40402 25394
rect 41246 25342 41298 25394
rect 45502 25342 45554 25394
rect 57038 25342 57090 25394
rect 57150 25342 57202 25394
rect 62190 25342 62242 25394
rect 63870 25342 63922 25394
rect 68574 25342 68626 25394
rect 69918 25342 69970 25394
rect 72494 25342 72546 25394
rect 8654 25230 8706 25282
rect 9214 25230 9266 25282
rect 9774 25230 9826 25282
rect 11790 25230 11842 25282
rect 12126 25230 12178 25282
rect 12574 25230 12626 25282
rect 17390 25230 17442 25282
rect 21758 25230 21810 25282
rect 22094 25230 22146 25282
rect 22878 25230 22930 25282
rect 28142 25230 28194 25282
rect 32846 25230 32898 25282
rect 38110 25230 38162 25282
rect 45614 25230 45666 25282
rect 56478 25230 56530 25282
rect 58270 25230 58322 25282
rect 58494 25230 58546 25282
rect 59502 25230 59554 25282
rect 59950 25230 60002 25282
rect 69694 25230 69746 25282
rect 72382 25230 72434 25282
rect 20534 25062 20586 25114
rect 20638 25062 20690 25114
rect 20742 25062 20794 25114
rect 39854 25062 39906 25114
rect 39958 25062 40010 25114
rect 40062 25062 40114 25114
rect 59174 25062 59226 25114
rect 59278 25062 59330 25114
rect 59382 25062 59434 25114
rect 78494 25062 78546 25114
rect 78598 25062 78650 25114
rect 78702 25062 78754 25114
rect 4286 24894 4338 24946
rect 10446 24894 10498 24946
rect 11454 24894 11506 24946
rect 15934 24894 15986 24946
rect 22654 24894 22706 24946
rect 27582 24894 27634 24946
rect 27694 24894 27746 24946
rect 44494 24894 44546 24946
rect 44606 24894 44658 24946
rect 44942 24894 44994 24946
rect 46846 24894 46898 24946
rect 59054 24894 59106 24946
rect 63422 24894 63474 24946
rect 64542 24894 64594 24946
rect 64766 24894 64818 24946
rect 65550 24894 65602 24946
rect 65774 24894 65826 24946
rect 66670 24894 66722 24946
rect 66782 24894 66834 24946
rect 72270 24894 72322 24946
rect 73278 24894 73330 24946
rect 74958 24894 75010 24946
rect 3614 24782 3666 24834
rect 4398 24782 4450 24834
rect 6414 24782 6466 24834
rect 8094 24782 8146 24834
rect 9886 24782 9938 24834
rect 10670 24782 10722 24834
rect 10782 24782 10834 24834
rect 12014 24782 12066 24834
rect 14254 24782 14306 24834
rect 18622 24782 18674 24834
rect 24446 24782 24498 24834
rect 26126 24782 26178 24834
rect 26686 24782 26738 24834
rect 30942 24782 30994 24834
rect 32734 24782 32786 24834
rect 32846 24782 32898 24834
rect 35422 24782 35474 24834
rect 37774 24782 37826 24834
rect 39454 24782 39506 24834
rect 43486 24782 43538 24834
rect 44046 24782 44098 24834
rect 48078 24782 48130 24834
rect 53342 24782 53394 24834
rect 53902 24782 53954 24834
rect 59278 24782 59330 24834
rect 59390 24782 59442 24834
rect 62414 24782 62466 24834
rect 64430 24782 64482 24834
rect 66558 24782 66610 24834
rect 69022 24782 69074 24834
rect 69806 24782 69858 24834
rect 72046 24782 72098 24834
rect 73502 24782 73554 24834
rect 75182 24782 75234 24834
rect 76862 24782 76914 24834
rect 77534 24782 77586 24834
rect 77646 24782 77698 24834
rect 2942 24670 2994 24722
rect 4062 24670 4114 24722
rect 7086 24670 7138 24722
rect 9662 24670 9714 24722
rect 9998 24670 10050 24722
rect 11566 24670 11618 24722
rect 13022 24670 13074 24722
rect 13582 24670 13634 24722
rect 13694 24670 13746 24722
rect 14366 24670 14418 24722
rect 14926 24670 14978 24722
rect 15822 24670 15874 24722
rect 16046 24670 16098 24722
rect 16494 24670 16546 24722
rect 19182 24670 19234 24722
rect 19854 24670 19906 24722
rect 20302 24670 20354 24722
rect 22766 24670 22818 24722
rect 22990 24670 23042 24722
rect 23102 24670 23154 24722
rect 26350 24670 26402 24722
rect 26574 24670 26626 24722
rect 30494 24670 30546 24722
rect 32510 24670 32562 24722
rect 33854 24670 33906 24722
rect 34526 24670 34578 24722
rect 35310 24670 35362 24722
rect 37102 24670 37154 24722
rect 37662 24670 37714 24722
rect 38894 24670 38946 24722
rect 42590 24670 42642 24722
rect 44270 24670 44322 24722
rect 46958 24670 47010 24722
rect 47854 24670 47906 24722
rect 52558 24670 52610 24722
rect 54014 24670 54066 24722
rect 54350 24670 54402 24722
rect 57710 24670 57762 24722
rect 58046 24670 58098 24722
rect 61854 24670 61906 24722
rect 65438 24670 65490 24722
rect 67790 24670 67842 24722
rect 70702 24670 70754 24722
rect 71374 24670 71426 24722
rect 71934 24670 71986 24722
rect 73614 24670 73666 24722
rect 75294 24670 75346 24722
rect 76302 24670 76354 24722
rect 3166 24558 3218 24610
rect 4846 24558 4898 24610
rect 7310 24558 7362 24610
rect 7982 24558 8034 24610
rect 9102 24558 9154 24610
rect 21534 24558 21586 24610
rect 21982 24558 22034 24610
rect 22878 24558 22930 24610
rect 23998 24558 24050 24610
rect 24894 24558 24946 24610
rect 25566 24558 25618 24610
rect 26686 24558 26738 24610
rect 28254 24558 28306 24610
rect 30046 24558 30098 24610
rect 34638 24558 34690 24610
rect 38782 24558 38834 24610
rect 42702 24558 42754 24610
rect 45390 24558 45442 24610
rect 52446 24558 52498 24610
rect 59950 24558 60002 24610
rect 60286 24558 60338 24610
rect 60734 24558 60786 24610
rect 61742 24558 61794 24610
rect 63870 24558 63922 24610
rect 67342 24558 67394 24610
rect 70590 24558 70642 24610
rect 74062 24558 74114 24610
rect 76414 24558 76466 24610
rect 8318 24446 8370 24498
rect 11454 24446 11506 24498
rect 21534 24446 21586 24498
rect 21758 24446 21810 24498
rect 22318 24446 22370 24498
rect 27806 24446 27858 24498
rect 35422 24446 35474 24498
rect 57934 24446 57986 24498
rect 63870 24446 63922 24498
rect 64206 24446 64258 24498
rect 77534 24446 77586 24498
rect 10874 24278 10926 24330
rect 10978 24278 11030 24330
rect 11082 24278 11134 24330
rect 30194 24278 30246 24330
rect 30298 24278 30350 24330
rect 30402 24278 30454 24330
rect 49514 24278 49566 24330
rect 49618 24278 49670 24330
rect 49722 24278 49774 24330
rect 68834 24278 68886 24330
rect 68938 24278 68990 24330
rect 69042 24278 69094 24330
rect 7310 24110 7362 24162
rect 7422 24110 7474 24162
rect 7646 24110 7698 24162
rect 9102 24110 9154 24162
rect 9550 24110 9602 24162
rect 9886 24110 9938 24162
rect 10110 24110 10162 24162
rect 19294 24110 19346 24162
rect 40462 24110 40514 24162
rect 41022 24110 41074 24162
rect 54014 24110 54066 24162
rect 64430 24110 64482 24162
rect 64766 24110 64818 24162
rect 65102 24110 65154 24162
rect 3950 23998 4002 24050
rect 4398 23998 4450 24050
rect 8430 23998 8482 24050
rect 11790 23998 11842 24050
rect 12238 23998 12290 24050
rect 12910 23998 12962 24050
rect 14478 23998 14530 24050
rect 17726 23998 17778 24050
rect 19518 23998 19570 24050
rect 19854 23998 19906 24050
rect 20862 23998 20914 24050
rect 21870 23998 21922 24050
rect 22990 23998 23042 24050
rect 26014 23998 26066 24050
rect 27246 23998 27298 24050
rect 34078 23998 34130 24050
rect 38110 23998 38162 24050
rect 39566 23998 39618 24050
rect 42030 23998 42082 24050
rect 44718 23998 44770 24050
rect 48414 23998 48466 24050
rect 49310 23998 49362 24050
rect 49758 23998 49810 24050
rect 57934 23998 57986 24050
rect 60398 23998 60450 24050
rect 64766 23998 64818 24050
rect 71822 23998 71874 24050
rect 75518 23998 75570 24050
rect 77310 23998 77362 24050
rect 2830 23886 2882 23938
rect 7870 23886 7922 23938
rect 10558 23886 10610 23938
rect 11118 23886 11170 23938
rect 13694 23886 13746 23938
rect 14030 23886 14082 23938
rect 18622 23886 18674 23938
rect 19742 23886 19794 23938
rect 23102 23886 23154 23938
rect 23326 23886 23378 23938
rect 26126 23886 26178 23938
rect 27470 23886 27522 23938
rect 30606 23886 30658 23938
rect 33630 23886 33682 23938
rect 33966 23886 34018 23938
rect 34638 23886 34690 23938
rect 35422 23886 35474 23938
rect 35758 23886 35810 23938
rect 37998 23886 38050 23938
rect 38782 23886 38834 23938
rect 39118 23886 39170 23938
rect 41918 23886 41970 23938
rect 44270 23886 44322 23938
rect 44494 23886 44546 23938
rect 47518 23886 47570 23938
rect 47742 23886 47794 23938
rect 52782 23886 52834 23938
rect 53454 23886 53506 23938
rect 53678 23886 53730 23938
rect 56814 23886 56866 23938
rect 57822 23886 57874 23938
rect 58382 23886 58434 23938
rect 58942 23886 58994 23938
rect 61742 23886 61794 23938
rect 62078 23886 62130 23938
rect 65326 23886 65378 23938
rect 66334 23886 66386 23938
rect 66670 23886 66722 23938
rect 72158 23886 72210 23938
rect 76190 23886 76242 23938
rect 1934 23774 1986 23826
rect 3614 23774 3666 23826
rect 10670 23774 10722 23826
rect 11006 23774 11058 23826
rect 13918 23774 13970 23826
rect 18286 23774 18338 23826
rect 18398 23774 18450 23826
rect 23550 23774 23602 23826
rect 23998 23774 24050 23826
rect 24894 23774 24946 23826
rect 25454 23774 25506 23826
rect 27918 23774 27970 23826
rect 30270 23774 30322 23826
rect 38894 23774 38946 23826
rect 40126 23774 40178 23826
rect 41134 23774 41186 23826
rect 42366 23774 42418 23826
rect 52446 23774 52498 23826
rect 59054 23774 59106 23826
rect 59726 23774 59778 23826
rect 65438 23774 65490 23826
rect 72606 23774 72658 23826
rect 3838 23662 3890 23714
rect 9214 23662 9266 23714
rect 9662 23662 9714 23714
rect 17278 23662 17330 23714
rect 19966 23662 20018 23714
rect 22318 23662 22370 23714
rect 22990 23662 23042 23714
rect 24446 23662 24498 23714
rect 25678 23662 25730 23714
rect 25902 23662 25954 23714
rect 26798 23662 26850 23714
rect 26910 23662 26962 23714
rect 27022 23662 27074 23714
rect 30382 23662 30434 23714
rect 32622 23662 32674 23714
rect 34750 23662 34802 23714
rect 34974 23662 35026 23714
rect 35534 23662 35586 23714
rect 36878 23662 36930 23714
rect 37774 23662 37826 23714
rect 38222 23662 38274 23714
rect 40350 23662 40402 23714
rect 41246 23662 41298 23714
rect 42142 23662 42194 23714
rect 50990 23662 51042 23714
rect 52558 23662 52610 23714
rect 59278 23662 59330 23714
rect 59838 23662 59890 23714
rect 60062 23662 60114 23714
rect 61854 23662 61906 23714
rect 65662 23662 65714 23714
rect 66446 23662 66498 23714
rect 67006 23662 67058 23714
rect 67454 23662 67506 23714
rect 67902 23662 67954 23714
rect 20534 23494 20586 23546
rect 20638 23494 20690 23546
rect 20742 23494 20794 23546
rect 39854 23494 39906 23546
rect 39958 23494 40010 23546
rect 40062 23494 40114 23546
rect 59174 23494 59226 23546
rect 59278 23494 59330 23546
rect 59382 23494 59434 23546
rect 78494 23494 78546 23546
rect 78598 23494 78650 23546
rect 78702 23494 78754 23546
rect 11342 23326 11394 23378
rect 18062 23326 18114 23378
rect 18510 23326 18562 23378
rect 26798 23326 26850 23378
rect 35086 23326 35138 23378
rect 40462 23326 40514 23378
rect 41694 23326 41746 23378
rect 48078 23326 48130 23378
rect 50094 23326 50146 23378
rect 50318 23326 50370 23378
rect 53454 23326 53506 23378
rect 53566 23326 53618 23378
rect 57598 23326 57650 23378
rect 65326 23326 65378 23378
rect 73502 23326 73554 23378
rect 74846 23326 74898 23378
rect 4286 23214 4338 23266
rect 4510 23214 4562 23266
rect 9886 23214 9938 23266
rect 15038 23214 15090 23266
rect 19070 23214 19122 23266
rect 19182 23214 19234 23266
rect 20078 23214 20130 23266
rect 25902 23214 25954 23266
rect 26462 23214 26514 23266
rect 26574 23214 26626 23266
rect 28254 23214 28306 23266
rect 29822 23214 29874 23266
rect 34638 23214 34690 23266
rect 46174 23214 46226 23266
rect 47182 23214 47234 23266
rect 49870 23214 49922 23266
rect 52894 23214 52946 23266
rect 53678 23214 53730 23266
rect 53790 23214 53842 23266
rect 53902 23214 53954 23266
rect 67454 23214 67506 23266
rect 76414 23214 76466 23266
rect 3502 23102 3554 23154
rect 6974 23102 7026 23154
rect 8206 23102 8258 23154
rect 9774 23102 9826 23154
rect 13470 23102 13522 23154
rect 14814 23102 14866 23154
rect 16606 23102 16658 23154
rect 19406 23102 19458 23154
rect 20302 23102 20354 23154
rect 21310 23102 21362 23154
rect 21646 23102 21698 23154
rect 24110 23102 24162 23154
rect 24670 23102 24722 23154
rect 29150 23102 29202 23154
rect 34078 23102 34130 23154
rect 36766 23102 36818 23154
rect 38670 23102 38722 23154
rect 39566 23102 39618 23154
rect 40238 23102 40290 23154
rect 40574 23102 40626 23154
rect 41918 23102 41970 23154
rect 44718 23102 44770 23154
rect 45502 23102 45554 23154
rect 47854 23102 47906 23154
rect 50542 23102 50594 23154
rect 50990 23102 51042 23154
rect 52446 23102 52498 23154
rect 55582 23102 55634 23154
rect 56142 23102 56194 23154
rect 56702 23102 56754 23154
rect 57486 23102 57538 23154
rect 59950 23102 60002 23154
rect 60062 23102 60114 23154
rect 60174 23102 60226 23154
rect 60286 23102 60338 23154
rect 60622 23102 60674 23154
rect 61406 23102 61458 23154
rect 62750 23102 62802 23154
rect 64094 23102 64146 23154
rect 64654 23102 64706 23154
rect 66110 23102 66162 23154
rect 68574 23102 68626 23154
rect 71262 23102 71314 23154
rect 72158 23102 72210 23154
rect 73390 23102 73442 23154
rect 73614 23102 73666 23154
rect 73950 23102 74002 23154
rect 75742 23102 75794 23154
rect 3390 22990 3442 23042
rect 5070 22990 5122 23042
rect 6414 22990 6466 23042
rect 7758 22990 7810 23042
rect 13022 22990 13074 23042
rect 16382 22990 16434 23042
rect 23550 22990 23602 23042
rect 27806 22990 27858 23042
rect 34190 22990 34242 23042
rect 36206 22990 36258 23042
rect 37214 22990 37266 23042
rect 38110 22990 38162 23042
rect 39454 22990 39506 23042
rect 45614 22990 45666 23042
rect 48638 22990 48690 23042
rect 50206 22990 50258 23042
rect 52558 22990 52610 23042
rect 58158 22990 58210 23042
rect 58718 22990 58770 23042
rect 58942 22990 58994 23042
rect 61294 22990 61346 23042
rect 63534 22990 63586 23042
rect 65886 22990 65938 23042
rect 67118 22990 67170 23042
rect 69246 22990 69298 23042
rect 70590 22990 70642 23042
rect 71374 22990 71426 23042
rect 74734 22990 74786 23042
rect 75630 22990 75682 23042
rect 76862 22990 76914 23042
rect 3166 22878 3218 22930
rect 4622 22878 4674 22930
rect 6638 22878 6690 22930
rect 9886 22878 9938 22930
rect 16046 22878 16098 22930
rect 40798 22878 40850 22930
rect 41022 22878 41074 22930
rect 41582 22878 41634 22930
rect 46958 22878 47010 22930
rect 47294 22878 47346 22930
rect 48190 22878 48242 22930
rect 57598 22878 57650 22930
rect 59278 22878 59330 22930
rect 66446 22878 66498 22930
rect 10874 22710 10926 22762
rect 10978 22710 11030 22762
rect 11082 22710 11134 22762
rect 30194 22710 30246 22762
rect 30298 22710 30350 22762
rect 30402 22710 30454 22762
rect 49514 22710 49566 22762
rect 49618 22710 49670 22762
rect 49722 22710 49774 22762
rect 68834 22710 68886 22762
rect 68938 22710 68990 22762
rect 69042 22710 69094 22762
rect 3502 22542 3554 22594
rect 3838 22542 3890 22594
rect 10110 22542 10162 22594
rect 12574 22542 12626 22594
rect 16494 22542 16546 22594
rect 20638 22542 20690 22594
rect 40126 22542 40178 22594
rect 44494 22542 44546 22594
rect 48078 22542 48130 22594
rect 49534 22542 49586 22594
rect 59502 22542 59554 22594
rect 60286 22542 60338 22594
rect 2494 22430 2546 22482
rect 3054 22430 3106 22482
rect 5630 22430 5682 22482
rect 6190 22430 6242 22482
rect 8542 22430 8594 22482
rect 9438 22430 9490 22482
rect 12126 22430 12178 22482
rect 12910 22430 12962 22482
rect 13806 22430 13858 22482
rect 24222 22430 24274 22482
rect 25790 22430 25842 22482
rect 38558 22430 38610 22482
rect 40798 22430 40850 22482
rect 43822 22430 43874 22482
rect 48190 22430 48242 22482
rect 54350 22430 54402 22482
rect 54910 22430 54962 22482
rect 55918 22430 55970 22482
rect 56926 22430 56978 22482
rect 59838 22430 59890 22482
rect 60622 22430 60674 22482
rect 64206 22430 64258 22482
rect 66894 22430 66946 22482
rect 70590 22430 70642 22482
rect 72494 22430 72546 22482
rect 77422 22430 77474 22482
rect 4622 22318 4674 22370
rect 6526 22318 6578 22370
rect 6862 22318 6914 22370
rect 7646 22318 7698 22370
rect 8094 22318 8146 22370
rect 9326 22318 9378 22370
rect 13694 22318 13746 22370
rect 13918 22318 13970 22370
rect 14366 22318 14418 22370
rect 14702 22318 14754 22370
rect 16382 22318 16434 22370
rect 20190 22318 20242 22370
rect 20414 22318 20466 22370
rect 26686 22318 26738 22370
rect 32062 22318 32114 22370
rect 32510 22318 32562 22370
rect 32958 22318 33010 22370
rect 33406 22318 33458 22370
rect 33854 22318 33906 22370
rect 34078 22318 34130 22370
rect 37662 22318 37714 22370
rect 37886 22318 37938 22370
rect 40910 22318 40962 22370
rect 44270 22318 44322 22370
rect 45502 22318 45554 22370
rect 45726 22318 45778 22370
rect 45950 22318 46002 22370
rect 49422 22318 49474 22370
rect 52670 22318 52722 22370
rect 53902 22318 53954 22370
rect 57822 22318 57874 22370
rect 64766 22318 64818 22370
rect 65102 22318 65154 22370
rect 66670 22318 66722 22370
rect 67342 22318 67394 22370
rect 71150 22318 71202 22370
rect 71486 22318 71538 22370
rect 72270 22318 72322 22370
rect 72942 22318 72994 22370
rect 74398 22318 74450 22370
rect 74622 22318 74674 22370
rect 75630 22318 75682 22370
rect 75854 22318 75906 22370
rect 3726 22206 3778 22258
rect 4510 22206 4562 22258
rect 6750 22206 6802 22258
rect 12798 22206 12850 22258
rect 14926 22206 14978 22258
rect 15038 22206 15090 22258
rect 16494 22206 16546 22258
rect 20078 22206 20130 22258
rect 24782 22206 24834 22258
rect 25230 22206 25282 22258
rect 26350 22206 26402 22258
rect 27694 22206 27746 22258
rect 43038 22206 43090 22258
rect 47854 22206 47906 22258
rect 51438 22206 51490 22258
rect 51774 22206 51826 22258
rect 52334 22206 52386 22258
rect 53454 22206 53506 22258
rect 57486 22206 57538 22258
rect 58270 22206 58322 22258
rect 58606 22206 58658 22258
rect 59054 22206 59106 22258
rect 59166 22206 59218 22258
rect 63758 22206 63810 22258
rect 64878 22206 64930 22258
rect 65550 22206 65602 22258
rect 65662 22206 65714 22258
rect 68350 22206 68402 22258
rect 71262 22206 71314 22258
rect 74846 22206 74898 22258
rect 75406 22206 75458 22258
rect 77534 22206 77586 22258
rect 2158 22094 2210 22146
rect 4286 22094 4338 22146
rect 15486 22094 15538 22146
rect 17166 22094 17218 22146
rect 19966 22094 20018 22146
rect 21870 22094 21922 22146
rect 22318 22094 22370 22146
rect 26462 22094 26514 22146
rect 27358 22094 27410 22146
rect 27582 22094 27634 22146
rect 28142 22094 28194 22146
rect 28590 22094 28642 22146
rect 33966 22094 34018 22146
rect 36430 22094 36482 22146
rect 36766 22094 36818 22146
rect 41582 22094 41634 22146
rect 47294 22094 47346 22146
rect 52446 22094 52498 22146
rect 55470 22094 55522 22146
rect 56478 22094 56530 22146
rect 57598 22094 57650 22146
rect 58382 22094 58434 22146
rect 59390 22094 59442 22146
rect 60174 22094 60226 22146
rect 61294 22094 61346 22146
rect 65886 22094 65938 22146
rect 67118 22094 67170 22146
rect 67230 22094 67282 22146
rect 67902 22094 67954 22146
rect 77310 22094 77362 22146
rect 77758 22094 77810 22146
rect 20534 21926 20586 21978
rect 20638 21926 20690 21978
rect 20742 21926 20794 21978
rect 39854 21926 39906 21978
rect 39958 21926 40010 21978
rect 40062 21926 40114 21978
rect 59174 21926 59226 21978
rect 59278 21926 59330 21978
rect 59382 21926 59434 21978
rect 78494 21926 78546 21978
rect 78598 21926 78650 21978
rect 78702 21926 78754 21978
rect 2718 21758 2770 21810
rect 2942 21758 2994 21810
rect 5518 21758 5570 21810
rect 7758 21758 7810 21810
rect 8990 21758 9042 21810
rect 9774 21758 9826 21810
rect 10222 21758 10274 21810
rect 18286 21758 18338 21810
rect 20638 21758 20690 21810
rect 21198 21758 21250 21810
rect 24446 21758 24498 21810
rect 26238 21758 26290 21810
rect 32958 21758 33010 21810
rect 36654 21758 36706 21810
rect 37998 21758 38050 21810
rect 38446 21758 38498 21810
rect 40350 21758 40402 21810
rect 44494 21758 44546 21810
rect 44830 21758 44882 21810
rect 45390 21758 45442 21810
rect 47854 21758 47906 21810
rect 48078 21758 48130 21810
rect 49982 21758 50034 21810
rect 54238 21758 54290 21810
rect 56366 21758 56418 21810
rect 57822 21758 57874 21810
rect 59502 21758 59554 21810
rect 63198 21758 63250 21810
rect 63758 21758 63810 21810
rect 65774 21758 65826 21810
rect 76862 21758 76914 21810
rect 77086 21758 77138 21810
rect 2606 21646 2658 21698
rect 4062 21646 4114 21698
rect 5406 21646 5458 21698
rect 6974 21646 7026 21698
rect 7198 21646 7250 21698
rect 8206 21646 8258 21698
rect 8878 21646 8930 21698
rect 12574 21646 12626 21698
rect 16830 21646 16882 21698
rect 18174 21646 18226 21698
rect 21422 21646 21474 21698
rect 22094 21646 22146 21698
rect 23662 21646 23714 21698
rect 25678 21646 25730 21698
rect 29710 21646 29762 21698
rect 31950 21646 32002 21698
rect 32734 21646 32786 21698
rect 35758 21646 35810 21698
rect 37886 21646 37938 21698
rect 40126 21646 40178 21698
rect 42478 21646 42530 21698
rect 44270 21646 44322 21698
rect 48638 21646 48690 21698
rect 53566 21646 53618 21698
rect 60510 21646 60562 21698
rect 61518 21646 61570 21698
rect 65550 21646 65602 21698
rect 71710 21646 71762 21698
rect 76750 21646 76802 21698
rect 4286 21534 4338 21586
rect 6638 21534 6690 21586
rect 7310 21534 7362 21586
rect 9998 21534 10050 21586
rect 13022 21534 13074 21586
rect 16718 21534 16770 21586
rect 17054 21534 17106 21586
rect 18062 21534 18114 21586
rect 18398 21534 18450 21586
rect 19518 21534 19570 21586
rect 20750 21534 20802 21586
rect 21534 21534 21586 21586
rect 24894 21534 24946 21586
rect 25902 21534 25954 21586
rect 26126 21534 26178 21586
rect 27582 21534 27634 21586
rect 29150 21534 29202 21586
rect 32062 21534 32114 21586
rect 32622 21534 32674 21586
rect 36094 21534 36146 21586
rect 36654 21534 36706 21586
rect 37326 21534 37378 21586
rect 37774 21534 37826 21586
rect 40014 21534 40066 21586
rect 42142 21534 42194 21586
rect 44158 21534 44210 21586
rect 47742 21534 47794 21586
rect 48526 21534 48578 21586
rect 48862 21534 48914 21586
rect 49422 21534 49474 21586
rect 49870 21534 49922 21586
rect 50094 21534 50146 21586
rect 55918 21534 55970 21586
rect 58046 21534 58098 21586
rect 59054 21534 59106 21586
rect 60734 21534 60786 21586
rect 61294 21534 61346 21586
rect 61630 21534 61682 21586
rect 64318 21534 64370 21586
rect 65438 21534 65490 21586
rect 66558 21534 66610 21586
rect 71150 21534 71202 21586
rect 74398 21534 74450 21586
rect 74958 21534 75010 21586
rect 2158 21422 2210 21474
rect 9886 21422 9938 21474
rect 13470 21422 13522 21474
rect 15262 21422 15314 21474
rect 16158 21422 16210 21474
rect 19966 21422 20018 21474
rect 22542 21422 22594 21474
rect 23102 21422 23154 21474
rect 26014 21422 26066 21474
rect 26798 21422 26850 21474
rect 27470 21422 27522 21474
rect 39006 21422 39058 21474
rect 39454 21422 39506 21474
rect 40686 21422 40738 21474
rect 42030 21422 42082 21474
rect 45838 21422 45890 21474
rect 53678 21422 53730 21474
rect 53790 21422 53842 21474
rect 55470 21422 55522 21474
rect 58606 21422 58658 21474
rect 59950 21422 60002 21474
rect 66334 21422 66386 21474
rect 67454 21422 67506 21474
rect 67790 21422 67842 21474
rect 69470 21422 69522 21474
rect 69806 21422 69858 21474
rect 70814 21422 70866 21474
rect 76078 21422 76130 21474
rect 17726 21310 17778 21362
rect 20638 21310 20690 21362
rect 40462 21310 40514 21362
rect 40686 21310 40738 21362
rect 55694 21310 55746 21362
rect 66894 21310 66946 21362
rect 10874 21142 10926 21194
rect 10978 21142 11030 21194
rect 11082 21142 11134 21194
rect 30194 21142 30246 21194
rect 30298 21142 30350 21194
rect 30402 21142 30454 21194
rect 49514 21142 49566 21194
rect 49618 21142 49670 21194
rect 49722 21142 49774 21194
rect 68834 21142 68886 21194
rect 68938 21142 68990 21194
rect 69042 21142 69094 21194
rect 3950 20974 4002 21026
rect 16382 20974 16434 21026
rect 26574 20974 26626 21026
rect 27246 20974 27298 21026
rect 34974 20974 35026 21026
rect 36542 20974 36594 21026
rect 41582 20974 41634 21026
rect 49870 20974 49922 21026
rect 55806 20974 55858 21026
rect 62302 20974 62354 21026
rect 69918 20974 69970 21026
rect 1934 20862 1986 20914
rect 4174 20862 4226 20914
rect 6526 20862 6578 20914
rect 7646 20862 7698 20914
rect 8654 20862 8706 20914
rect 11118 20862 11170 20914
rect 13806 20862 13858 20914
rect 17726 20862 17778 20914
rect 21870 20862 21922 20914
rect 22990 20862 23042 20914
rect 23998 20862 24050 20914
rect 25902 20862 25954 20914
rect 27470 20862 27522 20914
rect 30270 20862 30322 20914
rect 36094 20862 36146 20914
rect 38110 20862 38162 20914
rect 39230 20862 39282 20914
rect 40686 20862 40738 20914
rect 41918 20862 41970 20914
rect 46062 20862 46114 20914
rect 46510 20862 46562 20914
rect 48638 20862 48690 20914
rect 55022 20862 55074 20914
rect 56142 20862 56194 20914
rect 57934 20862 57986 20914
rect 58718 20862 58770 20914
rect 64542 20862 64594 20914
rect 66110 20862 66162 20914
rect 71038 20862 71090 20914
rect 72158 20862 72210 20914
rect 72718 20862 72770 20914
rect 74062 20862 74114 20914
rect 75518 20862 75570 20914
rect 77534 20862 77586 20914
rect 3054 20750 3106 20802
rect 4622 20750 4674 20802
rect 7198 20750 7250 20802
rect 8206 20750 8258 20802
rect 10670 20750 10722 20802
rect 11566 20750 11618 20802
rect 13694 20750 13746 20802
rect 14366 20750 14418 20802
rect 16606 20750 16658 20802
rect 17950 20750 18002 20802
rect 21646 20750 21698 20802
rect 22094 20750 22146 20802
rect 23550 20750 23602 20802
rect 27694 20750 27746 20802
rect 28478 20750 28530 20802
rect 33854 20750 33906 20802
rect 34414 20750 34466 20802
rect 34638 20750 34690 20802
rect 35758 20750 35810 20802
rect 38670 20750 38722 20802
rect 39342 20750 39394 20802
rect 40350 20750 40402 20802
rect 45838 20750 45890 20802
rect 48302 20750 48354 20802
rect 49646 20750 49698 20802
rect 54126 20750 54178 20802
rect 54350 20750 54402 20802
rect 55582 20750 55634 20802
rect 58606 20750 58658 20802
rect 59838 20750 59890 20802
rect 60398 20750 60450 20802
rect 60622 20750 60674 20802
rect 61742 20750 61794 20802
rect 61966 20750 62018 20802
rect 62974 20750 63026 20802
rect 63422 20750 63474 20802
rect 63870 20750 63922 20802
rect 65214 20750 65266 20802
rect 65550 20750 65602 20802
rect 67566 20750 67618 20802
rect 69582 20750 69634 20802
rect 70366 20750 70418 20802
rect 71598 20750 71650 20802
rect 73726 20750 73778 20802
rect 74286 20750 74338 20802
rect 75182 20750 75234 20802
rect 77310 20750 77362 20802
rect 77870 20750 77922 20802
rect 4958 20638 5010 20690
rect 6078 20638 6130 20690
rect 9214 20638 9266 20690
rect 9326 20638 9378 20690
rect 9886 20638 9938 20690
rect 10558 20638 10610 20690
rect 19630 20638 19682 20690
rect 20526 20638 20578 20690
rect 20750 20638 20802 20690
rect 20862 20638 20914 20690
rect 21870 20638 21922 20690
rect 22318 20638 22370 20690
rect 25566 20638 25618 20690
rect 26462 20638 26514 20690
rect 28814 20638 28866 20690
rect 30606 20638 30658 20690
rect 32062 20638 32114 20690
rect 39902 20638 39954 20690
rect 42142 20638 42194 20690
rect 44606 20638 44658 20690
rect 44718 20638 44770 20690
rect 52334 20638 52386 20690
rect 52670 20638 52722 20690
rect 53454 20638 53506 20690
rect 56142 20638 56194 20690
rect 56366 20638 56418 20690
rect 65326 20638 65378 20690
rect 66334 20638 66386 20690
rect 68238 20638 68290 20690
rect 69358 20638 69410 20690
rect 70814 20638 70866 20690
rect 72270 20638 72322 20690
rect 73838 20638 73890 20690
rect 74734 20638 74786 20690
rect 3614 20526 3666 20578
rect 4846 20526 4898 20578
rect 5630 20526 5682 20578
rect 9550 20526 9602 20578
rect 10334 20526 10386 20578
rect 13918 20526 13970 20578
rect 18734 20526 18786 20578
rect 19182 20526 19234 20578
rect 20078 20526 20130 20578
rect 24558 20526 24610 20578
rect 25118 20526 25170 20578
rect 26574 20526 26626 20578
rect 27806 20526 27858 20578
rect 27918 20526 27970 20578
rect 28702 20526 28754 20578
rect 29598 20526 29650 20578
rect 31950 20526 32002 20578
rect 37774 20526 37826 20578
rect 38894 20526 38946 20578
rect 39118 20526 39170 20578
rect 44382 20526 44434 20578
rect 69806 20526 69858 20578
rect 70926 20526 70978 20578
rect 71150 20526 71202 20578
rect 72046 20526 72098 20578
rect 20534 20358 20586 20410
rect 20638 20358 20690 20410
rect 20742 20358 20794 20410
rect 39854 20358 39906 20410
rect 39958 20358 40010 20410
rect 40062 20358 40114 20410
rect 59174 20358 59226 20410
rect 59278 20358 59330 20410
rect 59382 20358 59434 20410
rect 78494 20358 78546 20410
rect 78598 20358 78650 20410
rect 78702 20358 78754 20410
rect 14814 20190 14866 20242
rect 20862 20190 20914 20242
rect 27246 20190 27298 20242
rect 27470 20190 27522 20242
rect 29710 20190 29762 20242
rect 39790 20190 39842 20242
rect 44494 20190 44546 20242
rect 45390 20190 45442 20242
rect 54238 20190 54290 20242
rect 55918 20190 55970 20242
rect 59838 20190 59890 20242
rect 65326 20190 65378 20242
rect 67342 20190 67394 20242
rect 74398 20190 74450 20242
rect 4622 20078 4674 20130
rect 5854 20078 5906 20130
rect 10110 20078 10162 20130
rect 11678 20078 11730 20130
rect 12014 20078 12066 20130
rect 15038 20078 15090 20130
rect 17838 20078 17890 20130
rect 24222 20078 24274 20130
rect 25902 20078 25954 20130
rect 28254 20078 28306 20130
rect 35982 20078 36034 20130
rect 39566 20078 39618 20130
rect 40574 20078 40626 20130
rect 41582 20078 41634 20130
rect 41806 20078 41858 20130
rect 46286 20078 46338 20130
rect 46510 20078 46562 20130
rect 48414 20078 48466 20130
rect 48526 20078 48578 20130
rect 48638 20078 48690 20130
rect 60062 20078 60114 20130
rect 63086 20078 63138 20130
rect 67230 20078 67282 20130
rect 70366 20078 70418 20130
rect 76974 20078 77026 20130
rect 77534 20078 77586 20130
rect 1822 19966 1874 20018
rect 2382 19966 2434 20018
rect 3502 19966 3554 20018
rect 3726 19966 3778 20018
rect 3838 19966 3890 20018
rect 4174 19966 4226 20018
rect 5070 19966 5122 20018
rect 5742 19966 5794 20018
rect 5966 19966 6018 20018
rect 6414 19966 6466 20018
rect 14142 19966 14194 20018
rect 15150 19966 15202 20018
rect 18398 19966 18450 20018
rect 19182 19966 19234 20018
rect 19518 19966 19570 20018
rect 22318 19966 22370 20018
rect 24110 19966 24162 20018
rect 24334 19966 24386 20018
rect 24782 19966 24834 20018
rect 27582 19966 27634 20018
rect 28366 19966 28418 20018
rect 29598 19966 29650 20018
rect 29934 19966 29986 20018
rect 30382 19966 30434 20018
rect 30718 19966 30770 20018
rect 30830 19966 30882 20018
rect 31054 19966 31106 20018
rect 33742 19966 33794 20018
rect 35310 19966 35362 20018
rect 38670 19966 38722 20018
rect 39902 19966 39954 20018
rect 40686 19966 40738 20018
rect 44158 19966 44210 20018
rect 44942 19966 44994 20018
rect 45614 19966 45666 20018
rect 46174 19966 46226 20018
rect 49534 19966 49586 20018
rect 53566 19966 53618 20018
rect 54126 19966 54178 20018
rect 54462 19966 54514 20018
rect 55806 19966 55858 20018
rect 56030 19966 56082 20018
rect 56478 19966 56530 20018
rect 59614 19966 59666 20018
rect 60174 19966 60226 20018
rect 61966 19966 62018 20018
rect 64206 19966 64258 20018
rect 66670 19966 66722 20018
rect 66894 19966 66946 20018
rect 67118 19966 67170 20018
rect 69022 19966 69074 20018
rect 71262 19966 71314 20018
rect 71710 19966 71762 20018
rect 74062 19966 74114 20018
rect 74174 19966 74226 20018
rect 74622 19966 74674 20018
rect 75294 19966 75346 20018
rect 76750 19966 76802 20018
rect 77086 19966 77138 20018
rect 2718 19854 2770 19906
rect 3614 19854 3666 19906
rect 9886 19854 9938 19906
rect 13918 19854 13970 19906
rect 17054 19854 17106 19906
rect 21310 19854 21362 19906
rect 22766 19854 22818 19906
rect 23550 19854 23602 19906
rect 26350 19854 26402 19906
rect 26910 19854 26962 19906
rect 29038 19854 29090 19906
rect 30942 19854 30994 19906
rect 34302 19854 34354 19906
rect 35198 19854 35250 19906
rect 37102 19854 37154 19906
rect 39118 19854 39170 19906
rect 41918 19854 41970 19906
rect 43374 19854 43426 19906
rect 43934 19854 43986 19906
rect 45502 19854 45554 19906
rect 46846 19854 46898 19906
rect 53006 19854 53058 19906
rect 61630 19854 61682 19906
rect 62414 19854 62466 19906
rect 64766 19854 64818 19906
rect 65774 19854 65826 19906
rect 67902 19854 67954 19906
rect 68686 19854 68738 19906
rect 69694 19854 69746 19906
rect 70254 19854 70306 19906
rect 71934 19854 71986 19906
rect 73278 19854 73330 19906
rect 75406 19854 75458 19906
rect 4398 19742 4450 19794
rect 4958 19742 5010 19794
rect 13694 19742 13746 19794
rect 28254 19742 28306 19794
rect 34414 19742 34466 19794
rect 40798 19742 40850 19794
rect 49534 19742 49586 19794
rect 49870 19742 49922 19794
rect 53230 19742 53282 19794
rect 65662 19742 65714 19794
rect 65886 19742 65938 19794
rect 75630 19742 75682 19794
rect 10874 19574 10926 19626
rect 10978 19574 11030 19626
rect 11082 19574 11134 19626
rect 30194 19574 30246 19626
rect 30298 19574 30350 19626
rect 30402 19574 30454 19626
rect 49514 19574 49566 19626
rect 49618 19574 49670 19626
rect 49722 19574 49774 19626
rect 68834 19574 68886 19626
rect 68938 19574 68990 19626
rect 69042 19574 69094 19626
rect 4958 19406 5010 19458
rect 9438 19406 9490 19458
rect 25006 19406 25058 19458
rect 26238 19406 26290 19458
rect 30830 19406 30882 19458
rect 37550 19406 37602 19458
rect 38446 19406 38498 19458
rect 40462 19406 40514 19458
rect 43934 19406 43986 19458
rect 54350 19406 54402 19458
rect 60062 19406 60114 19458
rect 61854 19406 61906 19458
rect 64318 19406 64370 19458
rect 69470 19406 69522 19458
rect 4846 19294 4898 19346
rect 5854 19294 5906 19346
rect 6750 19294 6802 19346
rect 8318 19294 8370 19346
rect 14254 19294 14306 19346
rect 14702 19294 14754 19346
rect 16942 19294 16994 19346
rect 17278 19294 17330 19346
rect 18174 19294 18226 19346
rect 19630 19294 19682 19346
rect 22206 19294 22258 19346
rect 22654 19294 22706 19346
rect 28814 19294 28866 19346
rect 30270 19294 30322 19346
rect 35310 19294 35362 19346
rect 36094 19294 36146 19346
rect 36766 19294 36818 19346
rect 37662 19294 37714 19346
rect 38110 19294 38162 19346
rect 42702 19294 42754 19346
rect 43598 19294 43650 19346
rect 48078 19294 48130 19346
rect 50318 19294 50370 19346
rect 52334 19294 52386 19346
rect 53790 19294 53842 19346
rect 56590 19294 56642 19346
rect 57822 19294 57874 19346
rect 59726 19294 59778 19346
rect 63646 19294 63698 19346
rect 70478 19294 70530 19346
rect 74398 19294 74450 19346
rect 75518 19294 75570 19346
rect 77310 19294 77362 19346
rect 3054 19182 3106 19234
rect 3950 19182 4002 19234
rect 6078 19182 6130 19234
rect 8542 19182 8594 19234
rect 8878 19182 8930 19234
rect 9662 19182 9714 19234
rect 9886 19182 9938 19234
rect 13806 19182 13858 19234
rect 17054 19182 17106 19234
rect 17502 19182 17554 19234
rect 18286 19182 18338 19234
rect 19742 19182 19794 19234
rect 21534 19182 21586 19234
rect 23438 19182 23490 19234
rect 24110 19182 24162 19234
rect 25006 19182 25058 19234
rect 26350 19182 26402 19234
rect 27806 19182 27858 19234
rect 30494 19182 30546 19234
rect 31726 19182 31778 19234
rect 33854 19182 33906 19234
rect 34078 19182 34130 19234
rect 35870 19182 35922 19234
rect 39006 19182 39058 19234
rect 48190 19182 48242 19234
rect 49870 19182 49922 19234
rect 51102 19182 51154 19234
rect 53678 19182 53730 19234
rect 55806 19182 55858 19234
rect 56254 19182 56306 19234
rect 58046 19182 58098 19234
rect 59390 19182 59442 19234
rect 61518 19182 61570 19234
rect 61854 19182 61906 19234
rect 63198 19182 63250 19234
rect 64094 19182 64146 19234
rect 65438 19182 65490 19234
rect 66110 19182 66162 19234
rect 66782 19182 66834 19234
rect 70366 19182 70418 19234
rect 71262 19182 71314 19234
rect 76190 19182 76242 19234
rect 1934 19070 1986 19122
rect 3614 19070 3666 19122
rect 18174 19070 18226 19122
rect 18734 19070 18786 19122
rect 20190 19070 20242 19122
rect 26238 19070 26290 19122
rect 26910 19070 26962 19122
rect 27470 19070 27522 19122
rect 31390 19070 31442 19122
rect 34750 19070 34802 19122
rect 39566 19070 39618 19122
rect 39678 19070 39730 19122
rect 40350 19070 40402 19122
rect 40462 19070 40514 19122
rect 41582 19070 41634 19122
rect 42366 19070 42418 19122
rect 50990 19070 51042 19122
rect 57710 19070 57762 19122
rect 67566 19070 67618 19122
rect 69358 19070 69410 19122
rect 9998 18958 10050 19010
rect 10110 18958 10162 19010
rect 16270 18958 16322 19010
rect 16830 18958 16882 19010
rect 18510 18958 18562 19010
rect 19630 18958 19682 19010
rect 19966 18958 20018 19010
rect 20862 18958 20914 19010
rect 27582 18958 27634 19010
rect 28254 18958 28306 19010
rect 29710 18958 29762 19010
rect 31502 18958 31554 19010
rect 32174 18958 32226 19010
rect 38670 18958 38722 19010
rect 39902 18958 39954 19010
rect 41022 18958 41074 19010
rect 42590 18958 42642 19010
rect 43822 18958 43874 19010
rect 44494 18958 44546 19010
rect 45390 18958 45442 19010
rect 50766 18958 50818 19010
rect 51550 18958 51602 19010
rect 64654 18958 64706 19010
rect 68014 18958 68066 19010
rect 68574 18958 68626 19010
rect 69470 18958 69522 19010
rect 71710 18958 71762 19010
rect 20534 18790 20586 18842
rect 20638 18790 20690 18842
rect 20742 18790 20794 18842
rect 39854 18790 39906 18842
rect 39958 18790 40010 18842
rect 40062 18790 40114 18842
rect 59174 18790 59226 18842
rect 59278 18790 59330 18842
rect 59382 18790 59434 18842
rect 78494 18790 78546 18842
rect 78598 18790 78650 18842
rect 78702 18790 78754 18842
rect 2382 18622 2434 18674
rect 3838 18622 3890 18674
rect 8878 18622 8930 18674
rect 9886 18622 9938 18674
rect 16606 18622 16658 18674
rect 16830 18622 16882 18674
rect 18062 18622 18114 18674
rect 19854 18622 19906 18674
rect 23438 18622 23490 18674
rect 24222 18622 24274 18674
rect 24334 18622 24386 18674
rect 31390 18622 31442 18674
rect 34638 18622 34690 18674
rect 35646 18622 35698 18674
rect 35870 18622 35922 18674
rect 36654 18622 36706 18674
rect 37550 18622 37602 18674
rect 38894 18622 38946 18674
rect 45838 18622 45890 18674
rect 49534 18622 49586 18674
rect 49646 18622 49698 18674
rect 49758 18622 49810 18674
rect 51326 18622 51378 18674
rect 51662 18622 51714 18674
rect 55358 18622 55410 18674
rect 57598 18622 57650 18674
rect 59390 18622 59442 18674
rect 65550 18622 65602 18674
rect 71710 18622 71762 18674
rect 77646 18622 77698 18674
rect 1934 18510 1986 18562
rect 2830 18510 2882 18562
rect 3166 18510 3218 18562
rect 5854 18510 5906 18562
rect 6526 18510 6578 18562
rect 9774 18510 9826 18562
rect 11566 18510 11618 18562
rect 13246 18510 13298 18562
rect 15822 18510 15874 18562
rect 16942 18510 16994 18562
rect 17726 18510 17778 18562
rect 17838 18510 17890 18562
rect 18622 18510 18674 18562
rect 20078 18510 20130 18562
rect 20190 18510 20242 18562
rect 23550 18510 23602 18562
rect 25678 18510 25730 18562
rect 27806 18510 27858 18562
rect 29934 18510 29986 18562
rect 31278 18510 31330 18562
rect 34526 18510 34578 18562
rect 36542 18510 36594 18562
rect 38446 18510 38498 18562
rect 39006 18510 39058 18562
rect 43710 18510 43762 18562
rect 45614 18510 45666 18562
rect 47630 18510 47682 18562
rect 51886 18510 51938 18562
rect 53230 18510 53282 18562
rect 58942 18510 58994 18562
rect 59166 18510 59218 18562
rect 65662 18510 65714 18562
rect 68910 18510 68962 18562
rect 70030 18510 70082 18562
rect 73838 18510 73890 18562
rect 77534 18510 77586 18562
rect 77758 18510 77810 18562
rect 3950 18398 4002 18450
rect 5406 18398 5458 18450
rect 6414 18398 6466 18450
rect 8318 18398 8370 18450
rect 8654 18398 8706 18450
rect 8990 18398 9042 18450
rect 10110 18398 10162 18450
rect 14030 18398 14082 18450
rect 14478 18398 14530 18450
rect 18398 18398 18450 18450
rect 18734 18398 18786 18450
rect 19406 18398 19458 18450
rect 20638 18398 20690 18450
rect 21870 18398 21922 18450
rect 22878 18398 22930 18450
rect 23326 18398 23378 18450
rect 24894 18398 24946 18450
rect 26686 18398 26738 18450
rect 27134 18398 27186 18450
rect 27694 18398 27746 18450
rect 28030 18398 28082 18450
rect 30158 18398 30210 18450
rect 34862 18398 34914 18450
rect 35198 18398 35250 18450
rect 38670 18398 38722 18450
rect 40574 18398 40626 18450
rect 42254 18398 42306 18450
rect 45502 18398 45554 18450
rect 46958 18398 47010 18450
rect 50206 18398 50258 18450
rect 50654 18398 50706 18450
rect 51438 18398 51490 18450
rect 52334 18398 52386 18450
rect 53790 18398 53842 18450
rect 54798 18398 54850 18450
rect 58046 18398 58098 18450
rect 58158 18398 58210 18450
rect 58270 18398 58322 18450
rect 59726 18398 59778 18450
rect 61294 18398 61346 18450
rect 62078 18398 62130 18450
rect 64094 18398 64146 18450
rect 64654 18398 64706 18450
rect 65774 18398 65826 18450
rect 65886 18398 65938 18450
rect 67118 18398 67170 18450
rect 70702 18398 70754 18450
rect 71598 18398 71650 18450
rect 71822 18398 71874 18450
rect 72158 18398 72210 18450
rect 74622 18398 74674 18450
rect 75182 18398 75234 18450
rect 76078 18398 76130 18450
rect 76750 18398 76802 18450
rect 78094 18398 78146 18450
rect 4958 18286 5010 18338
rect 7870 18286 7922 18338
rect 10446 18286 10498 18338
rect 11342 18286 11394 18338
rect 13470 18286 13522 18338
rect 15262 18286 15314 18338
rect 16158 18286 16210 18338
rect 21422 18286 21474 18338
rect 22206 18286 22258 18338
rect 26238 18286 26290 18338
rect 28590 18286 28642 18338
rect 32062 18286 32114 18338
rect 32286 18286 32338 18338
rect 35758 18286 35810 18338
rect 37998 18286 38050 18338
rect 38894 18286 38946 18338
rect 40462 18286 40514 18338
rect 42590 18286 42642 18338
rect 43486 18286 43538 18338
rect 43822 18286 43874 18338
rect 44942 18286 44994 18338
rect 47182 18286 47234 18338
rect 51550 18286 51602 18338
rect 54126 18286 54178 18338
rect 55022 18286 55074 18338
rect 61742 18286 61794 18338
rect 66670 18286 66722 18338
rect 68350 18286 68402 18338
rect 69358 18286 69410 18338
rect 70926 18286 70978 18338
rect 73726 18286 73778 18338
rect 3838 18174 3890 18226
rect 6526 18174 6578 18226
rect 24446 18174 24498 18226
rect 32622 18174 32674 18226
rect 36654 18174 36706 18226
rect 39790 18174 39842 18226
rect 42366 18174 42418 18226
rect 59502 18174 59554 18226
rect 66222 18174 66274 18226
rect 74062 18174 74114 18226
rect 10874 18006 10926 18058
rect 10978 18006 11030 18058
rect 11082 18006 11134 18058
rect 30194 18006 30246 18058
rect 30298 18006 30350 18058
rect 30402 18006 30454 18058
rect 49514 18006 49566 18058
rect 49618 18006 49670 18058
rect 49722 18006 49774 18058
rect 68834 18006 68886 18058
rect 68938 18006 68990 18058
rect 69042 18006 69094 18058
rect 3950 17838 4002 17890
rect 5854 17838 5906 17890
rect 10110 17838 10162 17890
rect 12462 17838 12514 17890
rect 16270 17838 16322 17890
rect 19182 17838 19234 17890
rect 63870 17838 63922 17890
rect 64206 17838 64258 17890
rect 64878 17838 64930 17890
rect 65550 17838 65602 17890
rect 65774 17838 65826 17890
rect 74510 17838 74562 17890
rect 3838 17726 3890 17778
rect 4622 17726 4674 17778
rect 5742 17726 5794 17778
rect 7982 17726 8034 17778
rect 9550 17726 9602 17778
rect 10558 17726 10610 17778
rect 19742 17726 19794 17778
rect 20414 17726 20466 17778
rect 20974 17726 21026 17778
rect 22766 17726 22818 17778
rect 31166 17726 31218 17778
rect 32174 17726 32226 17778
rect 33630 17726 33682 17778
rect 34190 17726 34242 17778
rect 34526 17726 34578 17778
rect 37774 17726 37826 17778
rect 39678 17726 39730 17778
rect 41694 17726 41746 17778
rect 45838 17726 45890 17778
rect 47630 17726 47682 17778
rect 53342 17726 53394 17778
rect 58494 17726 58546 17778
rect 61854 17726 61906 17778
rect 63422 17726 63474 17778
rect 64878 17726 64930 17778
rect 65774 17726 65826 17778
rect 70142 17726 70194 17778
rect 71150 17726 71202 17778
rect 75182 17726 75234 17778
rect 2270 17614 2322 17666
rect 3614 17614 3666 17666
rect 6974 17614 7026 17666
rect 7534 17614 7586 17666
rect 8878 17614 8930 17666
rect 9662 17614 9714 17666
rect 9774 17614 9826 17666
rect 13582 17614 13634 17666
rect 16942 17614 16994 17666
rect 17614 17614 17666 17666
rect 18286 17614 18338 17666
rect 19070 17614 19122 17666
rect 22206 17614 22258 17666
rect 26798 17614 26850 17666
rect 28814 17614 28866 17666
rect 30494 17614 30546 17666
rect 31614 17614 31666 17666
rect 32510 17614 32562 17666
rect 35310 17614 35362 17666
rect 36430 17614 36482 17666
rect 36766 17614 36818 17666
rect 37886 17614 37938 17666
rect 39342 17614 39394 17666
rect 45726 17614 45778 17666
rect 46622 17614 46674 17666
rect 47518 17614 47570 17666
rect 51326 17614 51378 17666
rect 62078 17614 62130 17666
rect 69358 17614 69410 17666
rect 69806 17614 69858 17666
rect 71262 17614 71314 17666
rect 71486 17614 71538 17666
rect 74622 17614 74674 17666
rect 75630 17614 75682 17666
rect 76078 17614 76130 17666
rect 77310 17614 77362 17666
rect 77646 17614 77698 17666
rect 8542 17502 8594 17554
rect 11790 17502 11842 17554
rect 12574 17502 12626 17554
rect 13918 17502 13970 17554
rect 21870 17502 21922 17554
rect 26350 17502 26402 17554
rect 30158 17502 30210 17554
rect 31726 17502 31778 17554
rect 35198 17502 35250 17554
rect 35982 17502 36034 17554
rect 36542 17502 36594 17554
rect 38558 17502 38610 17554
rect 40238 17502 40290 17554
rect 41806 17502 41858 17554
rect 42030 17502 42082 17554
rect 50766 17502 50818 17554
rect 51438 17502 51490 17554
rect 52446 17502 52498 17554
rect 58046 17502 58098 17554
rect 58270 17502 58322 17554
rect 58606 17502 58658 17554
rect 61742 17502 61794 17554
rect 71038 17502 71090 17554
rect 73950 17502 74002 17554
rect 74510 17502 74562 17554
rect 77422 17502 77474 17554
rect 2046 17390 2098 17442
rect 4958 17390 5010 17442
rect 6862 17390 6914 17442
rect 7086 17390 7138 17442
rect 8654 17390 8706 17442
rect 9438 17390 9490 17442
rect 12462 17390 12514 17442
rect 13806 17390 13858 17442
rect 14366 17390 14418 17442
rect 14814 17390 14866 17442
rect 19182 17390 19234 17442
rect 21982 17390 22034 17442
rect 25790 17390 25842 17442
rect 26238 17390 26290 17442
rect 26462 17390 26514 17442
rect 28142 17390 28194 17442
rect 29598 17390 29650 17442
rect 30270 17390 30322 17442
rect 33294 17390 33346 17442
rect 34974 17390 35026 17442
rect 39566 17390 39618 17442
rect 40350 17390 40402 17442
rect 40574 17390 40626 17442
rect 40910 17390 40962 17442
rect 44718 17390 44770 17442
rect 47294 17390 47346 17442
rect 47742 17390 47794 17442
rect 48974 17390 49026 17442
rect 49422 17390 49474 17442
rect 50318 17390 50370 17442
rect 51662 17390 51714 17442
rect 52222 17390 52274 17442
rect 52334 17390 52386 17442
rect 63086 17390 63138 17442
rect 63870 17390 63922 17442
rect 64430 17390 64482 17442
rect 65326 17390 65378 17442
rect 73502 17390 73554 17442
rect 77982 17390 78034 17442
rect 20534 17222 20586 17274
rect 20638 17222 20690 17274
rect 20742 17222 20794 17274
rect 39854 17222 39906 17274
rect 39958 17222 40010 17274
rect 40062 17222 40114 17274
rect 59174 17222 59226 17274
rect 59278 17222 59330 17274
rect 59382 17222 59434 17274
rect 78494 17222 78546 17274
rect 78598 17222 78650 17274
rect 78702 17222 78754 17274
rect 9774 17054 9826 17106
rect 11902 17054 11954 17106
rect 12350 17054 12402 17106
rect 12798 17054 12850 17106
rect 13470 17054 13522 17106
rect 14590 17054 14642 17106
rect 17054 17054 17106 17106
rect 18174 17054 18226 17106
rect 19182 17054 19234 17106
rect 19630 17054 19682 17106
rect 20190 17054 20242 17106
rect 29150 17054 29202 17106
rect 30270 17054 30322 17106
rect 30494 17054 30546 17106
rect 32734 17054 32786 17106
rect 33518 17054 33570 17106
rect 38670 17054 38722 17106
rect 39230 17054 39282 17106
rect 40686 17054 40738 17106
rect 40910 17054 40962 17106
rect 47630 17054 47682 17106
rect 48638 17054 48690 17106
rect 50542 17054 50594 17106
rect 52782 17054 52834 17106
rect 52894 17054 52946 17106
rect 53678 17054 53730 17106
rect 58046 17054 58098 17106
rect 60286 17054 60338 17106
rect 60734 17054 60786 17106
rect 63086 17054 63138 17106
rect 70030 17054 70082 17106
rect 74062 17054 74114 17106
rect 3950 16942 4002 16994
rect 4734 16942 4786 16994
rect 13582 16942 13634 16994
rect 16830 16942 16882 16994
rect 32510 16942 32562 16994
rect 32846 16942 32898 16994
rect 42478 16942 42530 16994
rect 43822 16942 43874 16994
rect 46174 16942 46226 16994
rect 46286 16942 46338 16994
rect 49982 16942 50034 16994
rect 55470 16942 55522 16994
rect 61406 16942 61458 16994
rect 64654 16942 64706 16994
rect 67566 16942 67618 16994
rect 73726 16942 73778 16994
rect 76750 16942 76802 16994
rect 2046 16830 2098 16882
rect 3614 16830 3666 16882
rect 5294 16830 5346 16882
rect 6974 16830 7026 16882
rect 7870 16830 7922 16882
rect 10334 16830 10386 16882
rect 13246 16830 13298 16882
rect 14142 16830 14194 16882
rect 15710 16830 15762 16882
rect 16158 16830 16210 16882
rect 16718 16830 16770 16882
rect 17726 16830 17778 16882
rect 18286 16830 18338 16882
rect 18398 16830 18450 16882
rect 21534 16830 21586 16882
rect 22206 16830 22258 16882
rect 24334 16830 24386 16882
rect 24670 16830 24722 16882
rect 24782 16830 24834 16882
rect 24894 16830 24946 16882
rect 25902 16830 25954 16882
rect 27246 16830 27298 16882
rect 30158 16830 30210 16882
rect 31166 16830 31218 16882
rect 31838 16830 31890 16882
rect 32062 16830 32114 16882
rect 34974 16830 35026 16882
rect 35870 16830 35922 16882
rect 36542 16830 36594 16882
rect 36878 16830 36930 16882
rect 37550 16830 37602 16882
rect 37774 16830 37826 16882
rect 40126 16830 40178 16882
rect 40574 16830 40626 16882
rect 46510 16830 46562 16882
rect 46958 16830 47010 16882
rect 48190 16830 48242 16882
rect 49534 16830 49586 16882
rect 49758 16830 49810 16882
rect 50318 16830 50370 16882
rect 50990 16830 51042 16882
rect 51662 16830 51714 16882
rect 54238 16830 54290 16882
rect 55918 16830 55970 16882
rect 57486 16830 57538 16882
rect 61294 16830 61346 16882
rect 61630 16830 61682 16882
rect 61854 16830 61906 16882
rect 64094 16830 64146 16882
rect 64206 16830 64258 16882
rect 64430 16830 64482 16882
rect 65774 16830 65826 16882
rect 66894 16830 66946 16882
rect 67342 16830 67394 16882
rect 67454 16830 67506 16882
rect 69470 16830 69522 16882
rect 69694 16830 69746 16882
rect 73950 16830 74002 16882
rect 74174 16830 74226 16882
rect 75182 16830 75234 16882
rect 76078 16830 76130 16882
rect 77422 16830 77474 16882
rect 2494 16718 2546 16770
rect 3838 16718 3890 16770
rect 4510 16718 4562 16770
rect 4846 16718 4898 16770
rect 7086 16718 7138 16770
rect 8990 16718 9042 16770
rect 17950 16718 18002 16770
rect 20638 16718 20690 16770
rect 22878 16718 22930 16770
rect 23774 16718 23826 16770
rect 25790 16718 25842 16770
rect 28030 16718 28082 16770
rect 29598 16718 29650 16770
rect 35086 16718 35138 16770
rect 39566 16718 39618 16770
rect 42030 16718 42082 16770
rect 44046 16718 44098 16770
rect 45614 16718 45666 16770
rect 47070 16718 47122 16770
rect 51886 16718 51938 16770
rect 52670 16718 52722 16770
rect 54462 16718 54514 16770
rect 56366 16718 56418 16770
rect 57710 16718 57762 16770
rect 62638 16718 62690 16770
rect 64766 16718 64818 16770
rect 65550 16718 65602 16770
rect 66446 16718 66498 16770
rect 77086 16718 77138 16770
rect 10110 16606 10162 16658
rect 12014 16606 12066 16658
rect 13134 16606 13186 16658
rect 22094 16606 22146 16658
rect 37886 16606 37938 16658
rect 38782 16606 38834 16658
rect 39678 16606 39730 16658
rect 54798 16606 54850 16658
rect 62302 16606 62354 16658
rect 10874 16438 10926 16490
rect 10978 16438 11030 16490
rect 11082 16438 11134 16490
rect 30194 16438 30246 16490
rect 30298 16438 30350 16490
rect 30402 16438 30454 16490
rect 49514 16438 49566 16490
rect 49618 16438 49670 16490
rect 49722 16438 49774 16490
rect 68834 16438 68886 16490
rect 68938 16438 68990 16490
rect 69042 16438 69094 16490
rect 3054 16270 3106 16322
rect 4734 16270 4786 16322
rect 6862 16270 6914 16322
rect 7758 16270 7810 16322
rect 10222 16270 10274 16322
rect 11006 16270 11058 16322
rect 11902 16270 11954 16322
rect 41582 16270 41634 16322
rect 51550 16270 51602 16322
rect 51886 16270 51938 16322
rect 59502 16270 59554 16322
rect 64990 16270 65042 16322
rect 77422 16270 77474 16322
rect 2270 16158 2322 16210
rect 3166 16158 3218 16210
rect 4398 16158 4450 16210
rect 6190 16158 6242 16210
rect 14366 16158 14418 16210
rect 14814 16158 14866 16210
rect 16270 16158 16322 16210
rect 16718 16158 16770 16210
rect 17166 16158 17218 16210
rect 17950 16158 18002 16210
rect 19182 16158 19234 16210
rect 20302 16158 20354 16210
rect 26238 16158 26290 16210
rect 30270 16158 30322 16210
rect 32174 16158 32226 16210
rect 33854 16158 33906 16210
rect 35870 16158 35922 16210
rect 40238 16158 40290 16210
rect 40910 16158 40962 16210
rect 42142 16158 42194 16210
rect 48862 16158 48914 16210
rect 49870 16158 49922 16210
rect 50654 16158 50706 16210
rect 51326 16158 51378 16210
rect 55022 16158 55074 16210
rect 57486 16158 57538 16210
rect 59838 16158 59890 16210
rect 60622 16158 60674 16210
rect 61966 16158 62018 16210
rect 62638 16158 62690 16210
rect 62862 16158 62914 16210
rect 63646 16158 63698 16210
rect 66446 16158 66498 16210
rect 70366 16158 70418 16210
rect 72494 16158 72546 16210
rect 74398 16158 74450 16210
rect 75518 16158 75570 16210
rect 77982 16158 78034 16210
rect 3614 16046 3666 16098
rect 6638 16046 6690 16098
rect 7646 16046 7698 16098
rect 9662 16046 9714 16098
rect 11342 16046 11394 16098
rect 11454 16046 11506 16098
rect 11566 16046 11618 16098
rect 13918 16046 13970 16098
rect 18174 16046 18226 16098
rect 20414 16046 20466 16098
rect 21646 16046 21698 16098
rect 22206 16046 22258 16098
rect 22654 16046 22706 16098
rect 24222 16046 24274 16098
rect 24782 16046 24834 16098
rect 24894 16046 24946 16098
rect 26126 16046 26178 16098
rect 26910 16046 26962 16098
rect 27246 16046 27298 16098
rect 30830 16046 30882 16098
rect 31950 16046 32002 16098
rect 35086 16046 35138 16098
rect 35422 16046 35474 16098
rect 38446 16046 38498 16098
rect 39006 16046 39058 16098
rect 39902 16046 39954 16098
rect 40126 16046 40178 16098
rect 46286 16046 46338 16098
rect 46398 16046 46450 16098
rect 47630 16046 47682 16098
rect 48526 16046 48578 16098
rect 49422 16046 49474 16098
rect 54574 16046 54626 16098
rect 55582 16046 55634 16098
rect 55918 16046 55970 16098
rect 56590 16046 56642 16098
rect 56926 16046 56978 16098
rect 59950 16046 60002 16098
rect 61406 16046 61458 16098
rect 61854 16046 61906 16098
rect 62078 16046 62130 16098
rect 64318 16046 64370 16098
rect 65326 16046 65378 16098
rect 66222 16046 66274 16098
rect 69918 16046 69970 16098
rect 70142 16046 70194 16098
rect 72382 16046 72434 16098
rect 73278 16046 73330 16098
rect 74174 16046 74226 16098
rect 74846 16046 74898 16098
rect 75966 16046 76018 16098
rect 76302 16046 76354 16098
rect 4622 15934 4674 15986
rect 7758 15934 7810 15986
rect 9998 15934 10050 15986
rect 12574 15934 12626 15986
rect 12686 15934 12738 15986
rect 13806 15934 13858 15986
rect 17950 15934 18002 15986
rect 18398 15934 18450 15986
rect 19630 15934 19682 15986
rect 20302 15934 20354 15986
rect 20862 15934 20914 15986
rect 26462 15934 26514 15986
rect 27134 15934 27186 15986
rect 29598 15934 29650 15986
rect 32622 15934 32674 15986
rect 33518 15934 33570 15986
rect 34414 15934 34466 15986
rect 39118 15934 39170 15986
rect 39678 15934 39730 15986
rect 41582 15934 41634 15986
rect 41694 15934 41746 15986
rect 46622 15934 46674 15986
rect 47742 15934 47794 15986
rect 56366 15934 56418 15986
rect 57822 15934 57874 15986
rect 64878 15934 64930 15986
rect 66894 15934 66946 15986
rect 76078 15934 76130 15986
rect 77310 15934 77362 15986
rect 9214 15822 9266 15874
rect 9886 15822 9938 15874
rect 10446 15822 10498 15874
rect 11230 15822 11282 15874
rect 12350 15822 12402 15874
rect 13582 15822 13634 15874
rect 15262 15822 15314 15874
rect 15934 15822 15986 15874
rect 17838 15822 17890 15874
rect 20638 15822 20690 15874
rect 23326 15822 23378 15874
rect 25454 15822 25506 15874
rect 28814 15822 28866 15874
rect 29710 15822 29762 15874
rect 29934 15822 29986 15874
rect 30942 15822 30994 15874
rect 31166 15822 31218 15874
rect 33742 15822 33794 15874
rect 34526 15822 34578 15874
rect 34750 15822 34802 15874
rect 35310 15822 35362 15874
rect 37662 15822 37714 15874
rect 40238 15822 40290 15874
rect 42702 15822 42754 15874
rect 46174 15822 46226 15874
rect 47966 15822 48018 15874
rect 55694 15822 55746 15874
rect 56590 15822 56642 15874
rect 57598 15822 57650 15874
rect 61630 15822 61682 15874
rect 63198 15822 63250 15874
rect 64654 15822 64706 15874
rect 70814 15822 70866 15874
rect 71262 15822 71314 15874
rect 77422 15822 77474 15874
rect 20534 15654 20586 15706
rect 20638 15654 20690 15706
rect 20742 15654 20794 15706
rect 39854 15654 39906 15706
rect 39958 15654 40010 15706
rect 40062 15654 40114 15706
rect 59174 15654 59226 15706
rect 59278 15654 59330 15706
rect 59382 15654 59434 15706
rect 78494 15654 78546 15706
rect 78598 15654 78650 15706
rect 78702 15654 78754 15706
rect 2382 15486 2434 15538
rect 5854 15486 5906 15538
rect 11566 15486 11618 15538
rect 14478 15486 14530 15538
rect 15262 15486 15314 15538
rect 15710 15486 15762 15538
rect 17054 15486 17106 15538
rect 18510 15486 18562 15538
rect 19182 15486 19234 15538
rect 19406 15486 19458 15538
rect 19966 15486 20018 15538
rect 20638 15486 20690 15538
rect 21534 15486 21586 15538
rect 21646 15486 21698 15538
rect 28142 15486 28194 15538
rect 30494 15486 30546 15538
rect 31726 15486 31778 15538
rect 31950 15486 32002 15538
rect 34190 15486 34242 15538
rect 34302 15486 34354 15538
rect 35198 15486 35250 15538
rect 35646 15486 35698 15538
rect 39678 15486 39730 15538
rect 45502 15486 45554 15538
rect 46174 15486 46226 15538
rect 47294 15486 47346 15538
rect 50878 15486 50930 15538
rect 57374 15486 57426 15538
rect 60286 15486 60338 15538
rect 61294 15486 61346 15538
rect 61966 15486 62018 15538
rect 62302 15486 62354 15538
rect 64318 15486 64370 15538
rect 65886 15486 65938 15538
rect 69470 15486 69522 15538
rect 70254 15486 70306 15538
rect 71038 15486 71090 15538
rect 73726 15486 73778 15538
rect 75406 15486 75458 15538
rect 78094 15486 78146 15538
rect 2830 15374 2882 15426
rect 12686 15374 12738 15426
rect 16718 15374 16770 15426
rect 16830 15374 16882 15426
rect 21086 15374 21138 15426
rect 24558 15374 24610 15426
rect 43374 15374 43426 15426
rect 44046 15374 44098 15426
rect 44158 15374 44210 15426
rect 46398 15374 46450 15426
rect 46734 15374 46786 15426
rect 50542 15374 50594 15426
rect 50654 15374 50706 15426
rect 51214 15374 51266 15426
rect 70926 15374 70978 15426
rect 71598 15374 71650 15426
rect 73390 15374 73442 15426
rect 73502 15374 73554 15426
rect 74062 15374 74114 15426
rect 74510 15374 74562 15426
rect 76862 15374 76914 15426
rect 77534 15374 77586 15426
rect 3054 15262 3106 15314
rect 3950 15262 4002 15314
rect 5406 15262 5458 15314
rect 8542 15262 8594 15314
rect 11006 15262 11058 15314
rect 13246 15262 13298 15314
rect 13918 15262 13970 15314
rect 18062 15262 18114 15314
rect 18286 15262 18338 15314
rect 18734 15262 18786 15314
rect 19518 15262 19570 15314
rect 21310 15262 21362 15314
rect 22878 15262 22930 15314
rect 23998 15262 24050 15314
rect 28030 15262 28082 15314
rect 28254 15262 28306 15314
rect 28702 15262 28754 15314
rect 31838 15262 31890 15314
rect 32398 15262 32450 15314
rect 34414 15262 34466 15314
rect 34750 15262 34802 15314
rect 38782 15262 38834 15314
rect 39118 15262 39170 15314
rect 42478 15262 42530 15314
rect 43038 15262 43090 15314
rect 43822 15262 43874 15314
rect 44606 15262 44658 15314
rect 45950 15262 46002 15314
rect 46286 15262 46338 15314
rect 46846 15262 46898 15314
rect 47966 15262 48018 15314
rect 48414 15262 48466 15314
rect 51662 15262 51714 15314
rect 52782 15262 52834 15314
rect 53118 15262 53170 15314
rect 54126 15262 54178 15314
rect 60062 15262 60114 15314
rect 60398 15262 60450 15314
rect 60734 15262 60786 15314
rect 62974 15262 63026 15314
rect 63310 15262 63362 15314
rect 68910 15262 68962 15314
rect 70030 15262 70082 15314
rect 71262 15262 71314 15314
rect 76190 15262 76242 15314
rect 76750 15262 76802 15314
rect 77422 15262 77474 15314
rect 4510 15150 4562 15202
rect 4958 15150 5010 15202
rect 8990 15150 9042 15202
rect 9662 15150 9714 15202
rect 11230 15150 11282 15202
rect 16270 15150 16322 15202
rect 18398 15150 18450 15202
rect 21422 15150 21474 15202
rect 22430 15150 22482 15202
rect 23886 15150 23938 15202
rect 27470 15150 27522 15202
rect 30046 15150 30098 15202
rect 32174 15150 32226 15202
rect 38222 15150 38274 15202
rect 43150 15150 43202 15202
rect 62862 15150 62914 15202
rect 65326 15150 65378 15202
rect 70366 15150 70418 15202
rect 72494 15150 72546 15202
rect 54014 15038 54066 15090
rect 72606 15038 72658 15090
rect 77534 15038 77586 15090
rect 10874 14870 10926 14922
rect 10978 14870 11030 14922
rect 11082 14870 11134 14922
rect 30194 14870 30246 14922
rect 30298 14870 30350 14922
rect 30402 14870 30454 14922
rect 49514 14870 49566 14922
rect 49618 14870 49670 14922
rect 49722 14870 49774 14922
rect 68834 14870 68886 14922
rect 68938 14870 68990 14922
rect 69042 14870 69094 14922
rect 3726 14702 3778 14754
rect 13806 14702 13858 14754
rect 28030 14702 28082 14754
rect 28702 14702 28754 14754
rect 39790 14702 39842 14754
rect 46734 14702 46786 14754
rect 56702 14702 56754 14754
rect 58046 14702 58098 14754
rect 63870 14702 63922 14754
rect 64206 14702 64258 14754
rect 77422 14702 77474 14754
rect 5630 14590 5682 14642
rect 9438 14590 9490 14642
rect 17054 14590 17106 14642
rect 17614 14590 17666 14642
rect 19854 14590 19906 14642
rect 20302 14590 20354 14642
rect 20862 14590 20914 14642
rect 21646 14590 21698 14642
rect 22542 14590 22594 14642
rect 24670 14590 24722 14642
rect 26126 14590 26178 14642
rect 32510 14590 32562 14642
rect 36206 14590 36258 14642
rect 38222 14590 38274 14642
rect 42254 14590 42306 14642
rect 46174 14590 46226 14642
rect 49422 14590 49474 14642
rect 51998 14590 52050 14642
rect 57038 14590 57090 14642
rect 59614 14590 59666 14642
rect 61518 14590 61570 14642
rect 63646 14590 63698 14642
rect 67006 14590 67058 14642
rect 67902 14590 67954 14642
rect 69694 14590 69746 14642
rect 72382 14590 72434 14642
rect 73054 14590 73106 14642
rect 73950 14590 74002 14642
rect 74510 14590 74562 14642
rect 2830 14478 2882 14530
rect 4622 14478 4674 14530
rect 8094 14478 8146 14530
rect 8654 14478 8706 14530
rect 8766 14478 8818 14530
rect 9998 14478 10050 14530
rect 12462 14478 12514 14530
rect 12574 14478 12626 14530
rect 12910 14478 12962 14530
rect 13694 14478 13746 14530
rect 18062 14478 18114 14530
rect 19182 14478 19234 14530
rect 24222 14478 24274 14530
rect 25454 14478 25506 14530
rect 26014 14478 26066 14530
rect 28030 14478 28082 14530
rect 32398 14478 32450 14530
rect 33518 14478 33570 14530
rect 34750 14478 34802 14530
rect 34974 14478 35026 14530
rect 38446 14478 38498 14530
rect 40686 14478 40738 14530
rect 45950 14478 46002 14530
rect 48750 14478 48802 14530
rect 49310 14478 49362 14530
rect 51102 14478 51154 14530
rect 54014 14478 54066 14530
rect 54238 14478 54290 14530
rect 54910 14478 54962 14530
rect 57150 14478 57202 14530
rect 60062 14478 60114 14530
rect 60510 14478 60562 14530
rect 62078 14478 62130 14530
rect 62414 14478 62466 14530
rect 66894 14478 66946 14530
rect 67678 14478 67730 14530
rect 68014 14478 68066 14530
rect 70030 14478 70082 14530
rect 70478 14478 70530 14530
rect 71486 14478 71538 14530
rect 71710 14478 71762 14530
rect 73502 14478 73554 14530
rect 75070 14478 75122 14530
rect 77534 14478 77586 14530
rect 1934 14366 1986 14418
rect 3838 14366 3890 14418
rect 4510 14366 4562 14418
rect 7086 14366 7138 14418
rect 9326 14366 9378 14418
rect 12238 14366 12290 14418
rect 13806 14366 13858 14418
rect 14366 14366 14418 14418
rect 14590 14366 14642 14418
rect 14702 14366 14754 14418
rect 15598 14366 15650 14418
rect 23886 14366 23938 14418
rect 27694 14366 27746 14418
rect 28814 14366 28866 14418
rect 33966 14366 34018 14418
rect 39118 14366 39170 14418
rect 39902 14366 39954 14418
rect 40350 14366 40402 14418
rect 40574 14366 40626 14418
rect 42478 14366 42530 14418
rect 44158 14366 44210 14418
rect 44382 14366 44434 14418
rect 49982 14366 50034 14418
rect 50318 14366 50370 14418
rect 50766 14366 50818 14418
rect 54462 14366 54514 14418
rect 58158 14366 58210 14418
rect 62750 14366 62802 14418
rect 66110 14366 66162 14418
rect 68350 14366 68402 14418
rect 76078 14366 76130 14418
rect 3726 14254 3778 14306
rect 4286 14254 4338 14306
rect 6078 14254 6130 14306
rect 6638 14254 6690 14306
rect 7198 14254 7250 14306
rect 9550 14254 9602 14306
rect 12350 14254 12402 14306
rect 15150 14254 15202 14306
rect 16158 14254 16210 14306
rect 16494 14254 16546 14306
rect 21982 14254 22034 14306
rect 23998 14254 24050 14306
rect 28702 14254 28754 14306
rect 35310 14254 35362 14306
rect 35758 14254 35810 14306
rect 37662 14254 37714 14306
rect 39790 14254 39842 14306
rect 41582 14254 41634 14306
rect 50094 14254 50146 14306
rect 50878 14254 50930 14306
rect 58046 14254 58098 14306
rect 61406 14254 61458 14306
rect 61630 14254 61682 14306
rect 62638 14254 62690 14306
rect 77422 14254 77474 14306
rect 20534 14086 20586 14138
rect 20638 14086 20690 14138
rect 20742 14086 20794 14138
rect 39854 14086 39906 14138
rect 39958 14086 40010 14138
rect 40062 14086 40114 14138
rect 59174 14086 59226 14138
rect 59278 14086 59330 14138
rect 59382 14086 59434 14138
rect 78494 14086 78546 14138
rect 78598 14086 78650 14138
rect 78702 14086 78754 14138
rect 4510 13918 4562 13970
rect 9886 13918 9938 13970
rect 12014 13918 12066 13970
rect 16830 13918 16882 13970
rect 17054 13918 17106 13970
rect 18846 13918 18898 13970
rect 18958 13918 19010 13970
rect 19854 13918 19906 13970
rect 26238 13918 26290 13970
rect 35086 13918 35138 13970
rect 37662 13918 37714 13970
rect 40686 13918 40738 13970
rect 43150 13918 43202 13970
rect 43262 13918 43314 13970
rect 43374 13918 43426 13970
rect 46286 13918 46338 13970
rect 46510 13918 46562 13970
rect 48414 13918 48466 13970
rect 55134 13918 55186 13970
rect 64654 13918 64706 13970
rect 67230 13918 67282 13970
rect 67454 13918 67506 13970
rect 67790 13918 67842 13970
rect 72046 13918 72098 13970
rect 72158 13918 72210 13970
rect 2382 13806 2434 13858
rect 4062 13806 4114 13858
rect 4734 13806 4786 13858
rect 8654 13806 8706 13858
rect 12910 13806 12962 13858
rect 14814 13806 14866 13858
rect 23102 13806 23154 13858
rect 24782 13806 24834 13858
rect 26014 13806 26066 13858
rect 26686 13806 26738 13858
rect 30158 13806 30210 13858
rect 37886 13806 37938 13858
rect 37998 13806 38050 13858
rect 45390 13806 45442 13858
rect 46174 13806 46226 13858
rect 48638 13806 48690 13858
rect 49534 13806 49586 13858
rect 53790 13806 53842 13858
rect 61070 13806 61122 13858
rect 62526 13806 62578 13858
rect 65438 13806 65490 13858
rect 65550 13806 65602 13858
rect 67118 13806 67170 13858
rect 68238 13806 68290 13858
rect 73502 13806 73554 13858
rect 73614 13806 73666 13858
rect 75406 13806 75458 13858
rect 2270 13694 2322 13746
rect 2606 13694 2658 13746
rect 3390 13694 3442 13746
rect 4846 13694 4898 13746
rect 5742 13694 5794 13746
rect 8206 13694 8258 13746
rect 9774 13694 9826 13746
rect 11454 13694 11506 13746
rect 14142 13694 14194 13746
rect 16718 13694 16770 13746
rect 17838 13694 17890 13746
rect 18398 13694 18450 13746
rect 18622 13694 18674 13746
rect 19070 13694 19122 13746
rect 20974 13694 21026 13746
rect 22542 13694 22594 13746
rect 24670 13694 24722 13746
rect 25006 13694 25058 13746
rect 25566 13694 25618 13746
rect 27470 13694 27522 13746
rect 28142 13694 28194 13746
rect 29486 13694 29538 13746
rect 34750 13694 34802 13746
rect 34862 13694 34914 13746
rect 35310 13694 35362 13746
rect 35982 13694 36034 13746
rect 38894 13694 38946 13746
rect 39678 13694 39730 13746
rect 40238 13694 40290 13746
rect 40574 13694 40626 13746
rect 40798 13694 40850 13746
rect 43822 13694 43874 13746
rect 44942 13694 44994 13746
rect 48750 13694 48802 13746
rect 49982 13694 50034 13746
rect 54014 13694 54066 13746
rect 54910 13694 54962 13746
rect 55134 13694 55186 13746
rect 55470 13694 55522 13746
rect 59838 13694 59890 13746
rect 60286 13694 60338 13746
rect 62750 13694 62802 13746
rect 62974 13694 63026 13746
rect 65774 13694 65826 13746
rect 66558 13694 66610 13746
rect 71486 13694 71538 13746
rect 72270 13694 72322 13746
rect 72718 13694 72770 13746
rect 73278 13694 73330 13746
rect 75294 13694 75346 13746
rect 76862 13694 76914 13746
rect 1822 13582 1874 13634
rect 3614 13582 3666 13634
rect 5294 13582 5346 13634
rect 7758 13582 7810 13634
rect 12798 13582 12850 13634
rect 15262 13582 15314 13634
rect 15710 13582 15762 13634
rect 16158 13582 16210 13634
rect 20862 13582 20914 13634
rect 26126 13582 26178 13634
rect 28030 13582 28082 13634
rect 34078 13582 34130 13634
rect 35758 13582 35810 13634
rect 36318 13582 36370 13634
rect 37214 13582 37266 13634
rect 39118 13582 39170 13634
rect 44494 13582 44546 13634
rect 49870 13582 49922 13634
rect 59390 13582 59442 13634
rect 60958 13582 61010 13634
rect 61966 13582 62018 13634
rect 66110 13582 66162 13634
rect 69806 13582 69858 13634
rect 70366 13582 70418 13634
rect 70814 13582 70866 13634
rect 71374 13582 71426 13634
rect 76190 13582 76242 13634
rect 76974 13582 77026 13634
rect 9886 13470 9938 13522
rect 11678 13470 11730 13522
rect 17614 13470 17666 13522
rect 18174 13470 18226 13522
rect 54350 13470 54402 13522
rect 61294 13470 61346 13522
rect 75406 13470 75458 13522
rect 10874 13302 10926 13354
rect 10978 13302 11030 13354
rect 11082 13302 11134 13354
rect 30194 13302 30246 13354
rect 30298 13302 30350 13354
rect 30402 13302 30454 13354
rect 49514 13302 49566 13354
rect 49618 13302 49670 13354
rect 49722 13302 49774 13354
rect 68834 13302 68886 13354
rect 68938 13302 68990 13354
rect 69042 13302 69094 13354
rect 3390 13134 3442 13186
rect 13806 13134 13858 13186
rect 36654 13134 36706 13186
rect 38334 13134 38386 13186
rect 42590 13134 42642 13186
rect 44270 13134 44322 13186
rect 55358 13134 55410 13186
rect 55694 13134 55746 13186
rect 68462 13134 68514 13186
rect 76414 13134 76466 13186
rect 77310 13134 77362 13186
rect 2830 13022 2882 13074
rect 3614 13022 3666 13074
rect 3950 13022 4002 13074
rect 8990 13022 9042 13074
rect 12350 13022 12402 13074
rect 14366 13022 14418 13074
rect 15262 13022 15314 13074
rect 17166 13022 17218 13074
rect 17838 13022 17890 13074
rect 25230 13022 25282 13074
rect 32174 13022 32226 13074
rect 37886 13022 37938 13074
rect 43598 13022 43650 13074
rect 45950 13022 46002 13074
rect 48974 13022 49026 13074
rect 50990 13022 51042 13074
rect 54350 13022 54402 13074
rect 54462 13022 54514 13074
rect 59278 13022 59330 13074
rect 61518 13022 61570 13074
rect 64430 13022 64482 13074
rect 65438 13022 65490 13074
rect 66334 13022 66386 13074
rect 67230 13022 67282 13074
rect 71710 13022 71762 13074
rect 77870 13022 77922 13074
rect 3838 12910 3890 12962
rect 4062 12910 4114 12962
rect 18398 12910 18450 12962
rect 19070 12910 19122 12962
rect 19406 12910 19458 12962
rect 20414 12910 20466 12962
rect 20750 12910 20802 12962
rect 25006 12910 25058 12962
rect 25902 12910 25954 12962
rect 32622 12910 32674 12962
rect 33966 12910 34018 12962
rect 37774 12910 37826 12962
rect 39902 12910 39954 12962
rect 40350 12910 40402 12962
rect 40798 12910 40850 12962
rect 42478 12910 42530 12962
rect 43486 12910 43538 12962
rect 45838 12910 45890 12962
rect 49646 12910 49698 12962
rect 49870 12910 49922 12962
rect 53790 12910 53842 12962
rect 55134 12910 55186 12962
rect 56142 12910 56194 12962
rect 59950 12910 60002 12962
rect 60174 12910 60226 12962
rect 61294 12910 61346 12962
rect 61854 12910 61906 12962
rect 63982 12910 64034 12962
rect 64990 12910 65042 12962
rect 66782 12910 66834 12962
rect 67902 12910 67954 12962
rect 68126 12910 68178 12962
rect 71150 12910 71202 12962
rect 71374 12910 71426 12962
rect 71822 12910 71874 12962
rect 76078 12910 76130 12962
rect 76302 12910 76354 12962
rect 4846 12798 4898 12850
rect 4958 12798 5010 12850
rect 8430 12798 8482 12850
rect 8542 12798 8594 12850
rect 13694 12798 13746 12850
rect 13806 12798 13858 12850
rect 18510 12798 18562 12850
rect 18734 12798 18786 12850
rect 20302 12798 20354 12850
rect 21646 12798 21698 12850
rect 22094 12798 22146 12850
rect 29598 12798 29650 12850
rect 34190 12798 34242 12850
rect 36542 12798 36594 12850
rect 46062 12798 46114 12850
rect 51102 12798 51154 12850
rect 61742 12798 61794 12850
rect 70142 12798 70194 12850
rect 70254 12798 70306 12850
rect 77422 12798 77474 12850
rect 2046 12686 2098 12738
rect 2494 12686 2546 12738
rect 4622 12686 4674 12738
rect 7758 12686 7810 12738
rect 8206 12686 8258 12738
rect 11790 12686 11842 12738
rect 12798 12686 12850 12738
rect 14814 12686 14866 12738
rect 16158 12686 16210 12738
rect 16718 12686 16770 12738
rect 19294 12686 19346 12738
rect 20078 12686 20130 12738
rect 20190 12686 20242 12738
rect 27358 12686 27410 12738
rect 28030 12686 28082 12738
rect 29710 12686 29762 12738
rect 29934 12686 29986 12738
rect 30270 12686 30322 12738
rect 31502 12686 31554 12738
rect 35534 12686 35586 12738
rect 35982 12686 36034 12738
rect 36654 12686 36706 12738
rect 41918 12686 41970 12738
rect 42590 12686 42642 12738
rect 45614 12686 45666 12738
rect 50654 12686 50706 12738
rect 50878 12686 50930 12738
rect 52670 12686 52722 12738
rect 56926 12686 56978 12738
rect 62414 12686 62466 12738
rect 62862 12686 62914 12738
rect 69246 12686 69298 12738
rect 70478 12686 70530 12738
rect 71598 12686 71650 12738
rect 72382 12686 72434 12738
rect 20534 12518 20586 12570
rect 20638 12518 20690 12570
rect 20742 12518 20794 12570
rect 39854 12518 39906 12570
rect 39958 12518 40010 12570
rect 40062 12518 40114 12570
rect 59174 12518 59226 12570
rect 59278 12518 59330 12570
rect 59382 12518 59434 12570
rect 78494 12518 78546 12570
rect 78598 12518 78650 12570
rect 78702 12518 78754 12570
rect 8878 12350 8930 12402
rect 16158 12350 16210 12402
rect 17054 12350 17106 12402
rect 18286 12350 18338 12402
rect 19070 12350 19122 12402
rect 19294 12350 19346 12402
rect 19854 12350 19906 12402
rect 21086 12350 21138 12402
rect 22542 12350 22594 12402
rect 23326 12350 23378 12402
rect 37214 12350 37266 12402
rect 42926 12350 42978 12402
rect 48862 12350 48914 12402
rect 53118 12350 53170 12402
rect 55918 12350 55970 12402
rect 56590 12350 56642 12402
rect 58046 12350 58098 12402
rect 58494 12350 58546 12402
rect 61294 12350 61346 12402
rect 64654 12350 64706 12402
rect 65998 12350 66050 12402
rect 73502 12350 73554 12402
rect 74062 12350 74114 12402
rect 4174 12238 4226 12290
rect 5854 12238 5906 12290
rect 6078 12238 6130 12290
rect 8542 12238 8594 12290
rect 11790 12238 11842 12290
rect 12350 12238 12402 12290
rect 12462 12238 12514 12290
rect 13470 12238 13522 12290
rect 18174 12238 18226 12290
rect 20526 12238 20578 12290
rect 22206 12238 22258 12290
rect 22318 12238 22370 12290
rect 26686 12238 26738 12290
rect 30830 12238 30882 12290
rect 34750 12238 34802 12290
rect 48638 12238 48690 12290
rect 53566 12238 53618 12290
rect 55246 12238 55298 12290
rect 57486 12238 57538 12290
rect 60174 12238 60226 12290
rect 61966 12238 62018 12290
rect 62078 12238 62130 12290
rect 62526 12238 62578 12290
rect 63422 12238 63474 12290
rect 66670 12238 66722 12290
rect 66782 12238 66834 12290
rect 68798 12238 68850 12290
rect 71262 12238 71314 12290
rect 76750 12238 76802 12290
rect 2942 12126 2994 12178
rect 4510 12126 4562 12178
rect 8766 12126 8818 12178
rect 8990 12126 9042 12178
rect 9998 12126 10050 12178
rect 12686 12126 12738 12178
rect 13806 12126 13858 12178
rect 14814 12126 14866 12178
rect 16494 12126 16546 12178
rect 18958 12126 19010 12178
rect 20638 12126 20690 12178
rect 26014 12126 26066 12178
rect 27918 12126 27970 12178
rect 28814 12126 28866 12178
rect 30046 12126 30098 12178
rect 34190 12126 34242 12178
rect 39230 12126 39282 12178
rect 43822 12126 43874 12178
rect 48526 12126 48578 12178
rect 49758 12126 49810 12178
rect 54014 12126 54066 12178
rect 54462 12126 54514 12178
rect 56478 12126 56530 12178
rect 56814 12126 56866 12178
rect 59502 12126 59554 12178
rect 63198 12126 63250 12178
rect 63534 12126 63586 12178
rect 67006 12126 67058 12178
rect 67678 12126 67730 12178
rect 68238 12126 68290 12178
rect 70478 12126 70530 12178
rect 73390 12126 73442 12178
rect 73726 12126 73778 12178
rect 76190 12126 76242 12178
rect 77198 12126 77250 12178
rect 1934 12014 1986 12066
rect 10110 12014 10162 12066
rect 15374 12014 15426 12066
rect 17614 12014 17666 12066
rect 21534 12014 21586 12066
rect 22878 12014 22930 12066
rect 24894 12014 24946 12066
rect 25790 12014 25842 12066
rect 28590 12014 28642 12066
rect 34414 12014 34466 12066
rect 35982 12014 36034 12066
rect 38558 12014 38610 12066
rect 39566 12014 39618 12066
rect 42590 12014 42642 12066
rect 44158 12014 44210 12066
rect 49870 12014 49922 12066
rect 55134 12014 55186 12066
rect 59726 12014 59778 12066
rect 60734 12014 60786 12066
rect 63982 12014 64034 12066
rect 65550 12014 65602 12066
rect 69582 12014 69634 12066
rect 70366 12014 70418 12066
rect 75518 12014 75570 12066
rect 77534 12014 77586 12066
rect 10782 11902 10834 11954
rect 18286 11902 18338 11954
rect 20526 11902 20578 11954
rect 27582 11902 27634 11954
rect 27918 11902 27970 11954
rect 39678 11902 39730 11954
rect 44494 11902 44546 11954
rect 50094 11902 50146 11954
rect 60958 11902 61010 11954
rect 61966 11902 62018 11954
rect 10874 11734 10926 11786
rect 10978 11734 11030 11786
rect 11082 11734 11134 11786
rect 30194 11734 30246 11786
rect 30298 11734 30350 11786
rect 30402 11734 30454 11786
rect 49514 11734 49566 11786
rect 49618 11734 49670 11786
rect 49722 11734 49774 11786
rect 68834 11734 68886 11786
rect 68938 11734 68990 11786
rect 69042 11734 69094 11786
rect 8990 11566 9042 11618
rect 13694 11566 13746 11618
rect 44270 11566 44322 11618
rect 70030 11566 70082 11618
rect 71262 11566 71314 11618
rect 2046 11454 2098 11506
rect 3278 11454 3330 11506
rect 5742 11454 5794 11506
rect 8654 11454 8706 11506
rect 13022 11454 13074 11506
rect 16158 11454 16210 11506
rect 18622 11454 18674 11506
rect 20862 11454 20914 11506
rect 21646 11454 21698 11506
rect 21870 11454 21922 11506
rect 25006 11454 25058 11506
rect 26798 11454 26850 11506
rect 29710 11454 29762 11506
rect 34302 11454 34354 11506
rect 36206 11454 36258 11506
rect 43598 11454 43650 11506
rect 52334 11454 52386 11506
rect 54238 11454 54290 11506
rect 56366 11454 56418 11506
rect 57262 11454 57314 11506
rect 57934 11454 57986 11506
rect 62302 11454 62354 11506
rect 63310 11454 63362 11506
rect 63758 11454 63810 11506
rect 66222 11454 66274 11506
rect 66558 11454 66610 11506
rect 67006 11454 67058 11506
rect 67454 11454 67506 11506
rect 71150 11454 71202 11506
rect 74846 11454 74898 11506
rect 76526 11454 76578 11506
rect 77422 11454 77474 11506
rect 3166 11342 3218 11394
rect 3614 11342 3666 11394
rect 4174 11342 4226 11394
rect 4510 11342 4562 11394
rect 4734 11342 4786 11394
rect 8766 11342 8818 11394
rect 13918 11342 13970 11394
rect 14142 11342 14194 11394
rect 14254 11342 14306 11394
rect 15262 11342 15314 11394
rect 18062 11342 18114 11394
rect 18958 11342 19010 11394
rect 20190 11342 20242 11394
rect 22094 11342 22146 11394
rect 22206 11342 22258 11394
rect 24894 11342 24946 11394
rect 25790 11342 25842 11394
rect 26238 11342 26290 11394
rect 26686 11342 26738 11394
rect 26910 11342 26962 11394
rect 29598 11342 29650 11394
rect 33742 11342 33794 11394
rect 34190 11342 34242 11394
rect 34414 11342 34466 11394
rect 35534 11342 35586 11394
rect 40014 11342 40066 11394
rect 44158 11342 44210 11394
rect 48862 11342 48914 11394
rect 49310 11342 49362 11394
rect 51550 11342 51602 11394
rect 51998 11342 52050 11394
rect 54126 11342 54178 11394
rect 57038 11342 57090 11394
rect 58270 11342 58322 11394
rect 62190 11342 62242 11394
rect 63870 11342 63922 11394
rect 70142 11342 70194 11394
rect 71374 11342 71426 11394
rect 73838 11342 73890 11394
rect 74958 11342 75010 11394
rect 75630 11342 75682 11394
rect 75854 11342 75906 11394
rect 77758 11342 77810 11394
rect 5854 11230 5906 11282
rect 6078 11230 6130 11282
rect 16718 11230 16770 11282
rect 17726 11230 17778 11282
rect 30046 11230 30098 11282
rect 39678 11230 39730 11282
rect 40574 11230 40626 11282
rect 48750 11230 48802 11282
rect 53454 11230 53506 11282
rect 58942 11230 58994 11282
rect 60510 11230 60562 11282
rect 61518 11230 61570 11282
rect 77310 11230 77362 11282
rect 77646 11230 77698 11282
rect 4622 11118 4674 11170
rect 12014 11118 12066 11170
rect 12462 11118 12514 11170
rect 14366 11118 14418 11170
rect 14926 11118 14978 11170
rect 15150 11118 15202 11170
rect 15710 11118 15762 11170
rect 17278 11118 17330 11170
rect 17838 11118 17890 11170
rect 22318 11118 22370 11170
rect 28142 11118 28194 11170
rect 28814 11118 28866 11170
rect 29822 11118 29874 11170
rect 31054 11118 31106 11170
rect 34974 11118 35026 11170
rect 35646 11118 35698 11170
rect 35870 11118 35922 11170
rect 39118 11118 39170 11170
rect 39790 11118 39842 11170
rect 40462 11118 40514 11170
rect 41022 11118 41074 11170
rect 44270 11118 44322 11170
rect 48638 11118 48690 11170
rect 50990 11118 51042 11170
rect 55022 11118 55074 11170
rect 58046 11118 58098 11170
rect 64766 11118 64818 11170
rect 69470 11118 69522 11170
rect 70030 11118 70082 11170
rect 72270 11118 72322 11170
rect 74510 11118 74562 11170
rect 74734 11118 74786 11170
rect 20534 10950 20586 11002
rect 20638 10950 20690 11002
rect 20742 10950 20794 11002
rect 39854 10950 39906 11002
rect 39958 10950 40010 11002
rect 40062 10950 40114 11002
rect 59174 10950 59226 11002
rect 59278 10950 59330 11002
rect 59382 10950 59434 11002
rect 78494 10950 78546 11002
rect 78598 10950 78650 11002
rect 78702 10950 78754 11002
rect 2830 10782 2882 10834
rect 3838 10782 3890 10834
rect 8766 10782 8818 10834
rect 10558 10782 10610 10834
rect 11342 10782 11394 10834
rect 12798 10782 12850 10834
rect 13358 10782 13410 10834
rect 13582 10782 13634 10834
rect 14926 10782 14978 10834
rect 15934 10782 15986 10834
rect 17614 10782 17666 10834
rect 18622 10782 18674 10834
rect 20638 10782 20690 10834
rect 21310 10782 21362 10834
rect 25790 10782 25842 10834
rect 26014 10782 26066 10834
rect 26462 10782 26514 10834
rect 30830 10782 30882 10834
rect 45390 10782 45442 10834
rect 49422 10782 49474 10834
rect 52446 10782 52498 10834
rect 53006 10782 53058 10834
rect 53118 10782 53170 10834
rect 55806 10782 55858 10834
rect 56478 10782 56530 10834
rect 57710 10782 57762 10834
rect 62302 10782 62354 10834
rect 63086 10782 63138 10834
rect 63534 10782 63586 10834
rect 69358 10782 69410 10834
rect 70478 10782 70530 10834
rect 70814 10782 70866 10834
rect 2606 10670 2658 10722
rect 7870 10670 7922 10722
rect 8654 10670 8706 10722
rect 12462 10670 12514 10722
rect 12574 10670 12626 10722
rect 18174 10670 18226 10722
rect 21534 10670 21586 10722
rect 24334 10670 24386 10722
rect 25678 10670 25730 10722
rect 30494 10670 30546 10722
rect 30606 10670 30658 10722
rect 32958 10670 33010 10722
rect 44382 10670 44434 10722
rect 49646 10670 49698 10722
rect 53230 10670 53282 10722
rect 54238 10670 54290 10722
rect 54350 10670 54402 10722
rect 57822 10670 57874 10722
rect 61966 10670 62018 10722
rect 66670 10670 66722 10722
rect 69470 10670 69522 10722
rect 70142 10670 70194 10722
rect 70254 10670 70306 10722
rect 75742 10670 75794 10722
rect 77982 10670 78034 10722
rect 2494 10558 2546 10610
rect 3278 10558 3330 10610
rect 4398 10558 4450 10610
rect 6078 10558 6130 10610
rect 6414 10558 6466 10610
rect 7422 10558 7474 10610
rect 11118 10558 11170 10610
rect 11230 10558 11282 10610
rect 11678 10558 11730 10610
rect 13470 10558 13522 10610
rect 13694 10558 13746 10610
rect 13918 10558 13970 10610
rect 14366 10558 14418 10610
rect 15486 10558 15538 10610
rect 17054 10558 17106 10610
rect 18398 10558 18450 10610
rect 18734 10558 18786 10610
rect 19518 10558 19570 10610
rect 19966 10558 20018 10610
rect 21198 10558 21250 10610
rect 22318 10558 22370 10610
rect 23550 10558 23602 10610
rect 28254 10558 28306 10610
rect 29486 10558 29538 10610
rect 31502 10558 31554 10610
rect 32398 10558 32450 10610
rect 33854 10558 33906 10610
rect 35422 10558 35474 10610
rect 35870 10558 35922 10610
rect 38334 10558 38386 10610
rect 39230 10558 39282 10610
rect 40126 10558 40178 10610
rect 40798 10558 40850 10610
rect 42814 10558 42866 10610
rect 43822 10558 43874 10610
rect 44830 10558 44882 10610
rect 45278 10558 45330 10610
rect 45502 10558 45554 10610
rect 46958 10558 47010 10610
rect 47294 10558 47346 10610
rect 48302 10558 48354 10610
rect 49758 10558 49810 10610
rect 53678 10558 53730 10610
rect 54014 10558 54066 10610
rect 54798 10558 54850 10610
rect 56590 10558 56642 10610
rect 57486 10558 57538 10610
rect 62190 10558 62242 10610
rect 62414 10558 62466 10610
rect 63310 10558 63362 10610
rect 63422 10558 63474 10610
rect 65550 10558 65602 10610
rect 65998 10558 66050 10610
rect 67342 10558 67394 10610
rect 68574 10558 68626 10610
rect 72158 10558 72210 10610
rect 73726 10558 73778 10610
rect 74846 10558 74898 10610
rect 76414 10558 76466 10610
rect 76750 10558 76802 10610
rect 78094 10558 78146 10610
rect 1934 10446 1986 10498
rect 10446 10446 10498 10498
rect 16606 10446 16658 10498
rect 18510 10446 18562 10498
rect 22094 10446 22146 10498
rect 27806 10446 27858 10498
rect 29374 10446 29426 10498
rect 29822 10446 29874 10498
rect 31838 10446 31890 10498
rect 33966 10446 34018 10498
rect 36318 10446 36370 10498
rect 36878 10446 36930 10498
rect 38670 10446 38722 10498
rect 40014 10446 40066 10498
rect 41470 10446 41522 10498
rect 44046 10446 44098 10498
rect 50318 10446 50370 10498
rect 56702 10446 56754 10498
rect 58382 10446 58434 10498
rect 64654 10446 64706 10498
rect 67566 10446 67618 10498
rect 71822 10446 71874 10498
rect 72494 10446 72546 10498
rect 73390 10446 73442 10498
rect 73502 10446 73554 10498
rect 74958 10446 75010 10498
rect 76302 10446 76354 10498
rect 3502 10334 3554 10386
rect 4622 10334 4674 10386
rect 4958 10334 5010 10386
rect 8766 10334 8818 10386
rect 14142 10334 14194 10386
rect 14702 10334 14754 10386
rect 34414 10334 34466 10386
rect 42478 10334 42530 10386
rect 42814 10334 42866 10386
rect 48414 10334 48466 10386
rect 68238 10334 68290 10386
rect 68574 10334 68626 10386
rect 69246 10334 69298 10386
rect 77982 10334 78034 10386
rect 10874 10166 10926 10218
rect 10978 10166 11030 10218
rect 11082 10166 11134 10218
rect 30194 10166 30246 10218
rect 30298 10166 30350 10218
rect 30402 10166 30454 10218
rect 49514 10166 49566 10218
rect 49618 10166 49670 10218
rect 49722 10166 49774 10218
rect 68834 10166 68886 10218
rect 68938 10166 68990 10218
rect 69042 10166 69094 10218
rect 4510 9998 4562 10050
rect 7646 9998 7698 10050
rect 17390 9998 17442 10050
rect 19518 9998 19570 10050
rect 35534 9998 35586 10050
rect 43150 9998 43202 10050
rect 44606 9998 44658 10050
rect 57262 9998 57314 10050
rect 62414 9998 62466 10050
rect 63422 9998 63474 10050
rect 67566 9998 67618 10050
rect 72046 9998 72098 10050
rect 73278 9998 73330 10050
rect 76526 9998 76578 10050
rect 77646 9998 77698 10050
rect 77870 9998 77922 10050
rect 3726 9886 3778 9938
rect 7870 9886 7922 9938
rect 8206 9886 8258 9938
rect 11342 9886 11394 9938
rect 12574 9886 12626 9938
rect 15038 9886 15090 9938
rect 15598 9886 15650 9938
rect 18846 9886 18898 9938
rect 20750 9886 20802 9938
rect 21646 9886 21698 9938
rect 22318 9886 22370 9938
rect 26910 9886 26962 9938
rect 30270 9886 30322 9938
rect 30942 9886 30994 9938
rect 32286 9886 32338 9938
rect 35758 9886 35810 9938
rect 48526 9886 48578 9938
rect 65550 9886 65602 9938
rect 67230 9886 67282 9938
rect 68350 9886 68402 9938
rect 69470 9886 69522 9938
rect 72382 9886 72434 9938
rect 74958 9886 75010 9938
rect 76414 9886 76466 9938
rect 77982 9886 78034 9938
rect 4622 9774 4674 9826
rect 5630 9774 5682 9826
rect 8094 9774 8146 9826
rect 8878 9774 8930 9826
rect 11006 9774 11058 9826
rect 11678 9774 11730 9826
rect 13694 9774 13746 9826
rect 18398 9774 18450 9826
rect 18510 9774 18562 9826
rect 22878 9774 22930 9826
rect 25454 9774 25506 9826
rect 26014 9774 26066 9826
rect 26238 9774 26290 9826
rect 28478 9774 28530 9826
rect 29934 9774 29986 9826
rect 33518 9774 33570 9826
rect 35870 9774 35922 9826
rect 36430 9774 36482 9826
rect 38558 9774 38610 9826
rect 38894 9774 38946 9826
rect 39454 9774 39506 9826
rect 39902 9774 39954 9826
rect 40126 9774 40178 9826
rect 41134 9774 41186 9826
rect 41358 9774 41410 9826
rect 44718 9774 44770 9826
rect 45502 9774 45554 9826
rect 45726 9774 45778 9826
rect 45950 9774 46002 9826
rect 48638 9774 48690 9826
rect 49758 9774 49810 9826
rect 49982 9774 50034 9826
rect 51550 9774 51602 9826
rect 56702 9774 56754 9826
rect 57374 9774 57426 9826
rect 62414 9774 62466 9826
rect 67006 9774 67058 9826
rect 69694 9774 69746 9826
rect 70590 9774 70642 9826
rect 71038 9774 71090 9826
rect 71374 9774 71426 9826
rect 72942 9774 72994 9826
rect 2382 9662 2434 9714
rect 5966 9662 6018 9714
rect 17278 9662 17330 9714
rect 18174 9662 18226 9714
rect 19406 9662 19458 9714
rect 19518 9662 19570 9714
rect 23662 9662 23714 9714
rect 29598 9662 29650 9714
rect 33182 9662 33234 9714
rect 34974 9662 35026 9714
rect 36542 9662 36594 9714
rect 43486 9662 43538 9714
rect 44606 9662 44658 9714
rect 48302 9662 48354 9714
rect 50878 9662 50930 9714
rect 50990 9662 51042 9714
rect 59950 9662 60002 9714
rect 62750 9662 62802 9714
rect 63422 9662 63474 9714
rect 63534 9662 63586 9714
rect 70254 9662 70306 9714
rect 71150 9662 71202 9714
rect 72270 9662 72322 9714
rect 72494 9662 72546 9714
rect 72830 9662 72882 9714
rect 73166 9662 73218 9714
rect 73390 9662 73442 9714
rect 73614 9662 73666 9714
rect 73726 9662 73778 9714
rect 1934 9550 1986 9602
rect 2718 9550 2770 9602
rect 3278 9550 3330 9602
rect 4510 9550 4562 9602
rect 5854 9550 5906 9602
rect 6414 9550 6466 9602
rect 7086 9550 7138 9602
rect 8318 9550 8370 9602
rect 9438 9550 9490 9602
rect 9774 9550 9826 9602
rect 12910 9550 12962 9602
rect 13806 9550 13858 9602
rect 14030 9550 14082 9602
rect 14590 9550 14642 9602
rect 16270 9550 16322 9602
rect 16718 9550 16770 9602
rect 17390 9550 17442 9602
rect 18286 9550 18338 9602
rect 20190 9550 20242 9602
rect 22990 9550 23042 9602
rect 23214 9550 23266 9602
rect 23774 9550 23826 9602
rect 23998 9550 24050 9602
rect 24446 9550 24498 9602
rect 28142 9550 28194 9602
rect 29710 9550 29762 9602
rect 33294 9550 33346 9602
rect 33854 9550 33906 9602
rect 36766 9550 36818 9602
rect 37438 9550 37490 9602
rect 38670 9550 38722 9602
rect 40014 9550 40066 9602
rect 40574 9550 40626 9602
rect 41694 9550 41746 9602
rect 42142 9550 42194 9602
rect 42702 9550 42754 9602
rect 43262 9550 43314 9602
rect 43934 9550 43986 9602
rect 49198 9550 49250 9602
rect 50318 9550 50370 9602
rect 51214 9550 51266 9602
rect 52110 9550 52162 9602
rect 52558 9550 52610 9602
rect 53790 9550 53842 9602
rect 54350 9550 54402 9602
rect 54798 9550 54850 9602
rect 55246 9550 55298 9602
rect 55918 9550 55970 9602
rect 58046 9550 58098 9602
rect 58494 9550 58546 9602
rect 59054 9550 59106 9602
rect 59502 9550 59554 9602
rect 65102 9550 65154 9602
rect 66110 9550 66162 9602
rect 69470 9550 69522 9602
rect 70366 9550 70418 9602
rect 74622 9550 74674 9602
rect 75518 9550 75570 9602
rect 75854 9550 75906 9602
rect 77534 9550 77586 9602
rect 20534 9382 20586 9434
rect 20638 9382 20690 9434
rect 20742 9382 20794 9434
rect 39854 9382 39906 9434
rect 39958 9382 40010 9434
rect 40062 9382 40114 9434
rect 59174 9382 59226 9434
rect 59278 9382 59330 9434
rect 59382 9382 59434 9434
rect 78494 9382 78546 9434
rect 78598 9382 78650 9434
rect 78702 9382 78754 9434
rect 4734 9214 4786 9266
rect 7870 9214 7922 9266
rect 8094 9214 8146 9266
rect 8654 9214 8706 9266
rect 8878 9214 8930 9266
rect 14702 9214 14754 9266
rect 15150 9214 15202 9266
rect 20078 9214 20130 9266
rect 21646 9214 21698 9266
rect 22654 9214 22706 9266
rect 25006 9214 25058 9266
rect 25902 9214 25954 9266
rect 26126 9214 26178 9266
rect 26238 9214 26290 9266
rect 27022 9214 27074 9266
rect 28814 9214 28866 9266
rect 29486 9214 29538 9266
rect 30830 9214 30882 9266
rect 31390 9214 31442 9266
rect 32734 9214 32786 9266
rect 33854 9214 33906 9266
rect 34302 9214 34354 9266
rect 34974 9214 35026 9266
rect 35758 9214 35810 9266
rect 36542 9214 36594 9266
rect 37886 9214 37938 9266
rect 39566 9214 39618 9266
rect 40686 9214 40738 9266
rect 42142 9214 42194 9266
rect 43038 9214 43090 9266
rect 43598 9214 43650 9266
rect 44046 9214 44098 9266
rect 49982 9214 50034 9266
rect 62750 9214 62802 9266
rect 62862 9214 62914 9266
rect 63534 9214 63586 9266
rect 67230 9214 67282 9266
rect 69022 9214 69074 9266
rect 69582 9214 69634 9266
rect 70030 9214 70082 9266
rect 70926 9214 70978 9266
rect 71710 9214 71762 9266
rect 72270 9214 72322 9266
rect 73502 9214 73554 9266
rect 73614 9214 73666 9266
rect 77086 9214 77138 9266
rect 77422 9214 77474 9266
rect 5742 9102 5794 9154
rect 8990 9102 9042 9154
rect 11342 9102 11394 9154
rect 12014 9102 12066 9154
rect 19294 9102 19346 9154
rect 24334 9102 24386 9154
rect 26350 9102 26402 9154
rect 30606 9102 30658 9154
rect 32846 9102 32898 9154
rect 34862 9102 34914 9154
rect 36430 9102 36482 9154
rect 37326 9102 37378 9154
rect 40014 9102 40066 9154
rect 40574 9102 40626 9154
rect 48750 9102 48802 9154
rect 49422 9102 49474 9154
rect 50878 9102 50930 9154
rect 54350 9102 54402 9154
rect 56142 9102 56194 9154
rect 66782 9102 66834 9154
rect 67454 9102 67506 9154
rect 67566 9102 67618 9154
rect 68238 9102 68290 9154
rect 73390 9102 73442 9154
rect 76862 9102 76914 9154
rect 2830 8990 2882 9042
rect 4286 8990 4338 9042
rect 4622 8990 4674 9042
rect 4958 8990 5010 9042
rect 5518 8990 5570 9042
rect 5854 8990 5906 9042
rect 6750 8990 6802 9042
rect 7198 8990 7250 9042
rect 8206 8990 8258 9042
rect 10894 8990 10946 9042
rect 11902 8990 11954 9042
rect 13246 8990 13298 9042
rect 18062 8990 18114 9042
rect 18622 8990 18674 9042
rect 19182 8990 19234 9042
rect 19518 8990 19570 9042
rect 22094 8990 22146 9042
rect 23550 8990 23602 9042
rect 28142 8990 28194 9042
rect 28702 8990 28754 9042
rect 30494 8990 30546 9042
rect 31502 8990 31554 9042
rect 31614 8990 31666 9042
rect 31726 8990 31778 9042
rect 32062 8990 32114 9042
rect 32510 8990 32562 9042
rect 35198 8990 35250 9042
rect 35646 8990 35698 9042
rect 35982 8990 36034 9042
rect 37214 8990 37266 9042
rect 37550 8990 37602 9042
rect 40910 8990 40962 9042
rect 41582 8990 41634 9042
rect 41806 8990 41858 9042
rect 42030 8990 42082 9042
rect 42254 8990 42306 9042
rect 42926 8990 42978 9042
rect 43262 8990 43314 9042
rect 51214 8990 51266 9042
rect 52110 8990 52162 9042
rect 54798 8990 54850 9042
rect 55918 8990 55970 9042
rect 56590 8990 56642 9042
rect 57486 8990 57538 9042
rect 58046 8990 58098 9042
rect 58494 8990 58546 9042
rect 60174 8990 60226 9042
rect 60846 8990 60898 9042
rect 61518 8990 61570 9042
rect 62302 8990 62354 9042
rect 62974 8990 63026 9042
rect 64094 8990 64146 9042
rect 65438 8990 65490 9042
rect 68350 8990 68402 9042
rect 69134 8990 69186 9042
rect 71598 8990 71650 9042
rect 71934 8990 71986 9042
rect 73950 8990 74002 9042
rect 75966 8990 76018 9042
rect 76750 8990 76802 9042
rect 1934 8878 1986 8930
rect 3726 8878 3778 8930
rect 4846 8878 4898 8930
rect 9662 8878 9714 8930
rect 10446 8878 10498 8930
rect 15486 8878 15538 8930
rect 20526 8878 20578 8930
rect 20974 8878 21026 8930
rect 23774 8878 23826 8930
rect 27694 8878 27746 8930
rect 29934 8878 29986 8930
rect 38334 8878 38386 8930
rect 52782 8878 52834 8930
rect 53566 8878 53618 8930
rect 54686 8878 54738 8930
rect 56030 8878 56082 8930
rect 62526 8878 62578 8930
rect 64542 8878 64594 8930
rect 65774 8878 65826 8930
rect 66334 8878 66386 8930
rect 70478 8878 70530 8930
rect 74510 8878 74562 8930
rect 75518 8878 75570 8930
rect 77870 8878 77922 8930
rect 12014 8766 12066 8818
rect 13470 8766 13522 8818
rect 13806 8766 13858 8818
rect 28814 8766 28866 8818
rect 36542 8766 36594 8818
rect 59726 8766 59778 8818
rect 68238 8766 68290 8818
rect 69022 8766 69074 8818
rect 10874 8598 10926 8650
rect 10978 8598 11030 8650
rect 11082 8598 11134 8650
rect 30194 8598 30246 8650
rect 30298 8598 30350 8650
rect 30402 8598 30454 8650
rect 49514 8598 49566 8650
rect 49618 8598 49670 8650
rect 49722 8598 49774 8650
rect 68834 8598 68886 8650
rect 68938 8598 68990 8650
rect 69042 8598 69094 8650
rect 36430 8430 36482 8482
rect 51102 8430 51154 8482
rect 54910 8430 54962 8482
rect 56590 8430 56642 8482
rect 57374 8430 57426 8482
rect 2158 8318 2210 8370
rect 7198 8318 7250 8370
rect 7758 8318 7810 8370
rect 13918 8318 13970 8370
rect 20078 8318 20130 8370
rect 23438 8318 23490 8370
rect 24222 8318 24274 8370
rect 28590 8318 28642 8370
rect 30158 8318 30210 8370
rect 34862 8318 34914 8370
rect 35310 8318 35362 8370
rect 35758 8318 35810 8370
rect 38110 8318 38162 8370
rect 41470 8318 41522 8370
rect 45838 8318 45890 8370
rect 47518 8318 47570 8370
rect 50542 8318 50594 8370
rect 55582 8318 55634 8370
rect 60398 8318 60450 8370
rect 61630 8318 61682 8370
rect 63086 8318 63138 8370
rect 65774 8318 65826 8370
rect 67566 8318 67618 8370
rect 69246 8318 69298 8370
rect 70478 8318 70530 8370
rect 75406 8318 75458 8370
rect 77870 8318 77922 8370
rect 3054 8206 3106 8258
rect 3390 8206 3442 8258
rect 4286 8206 4338 8258
rect 4622 8206 4674 8258
rect 4846 8206 4898 8258
rect 8878 8206 8930 8258
rect 9326 8206 9378 8258
rect 9774 8206 9826 8258
rect 15262 8206 15314 8258
rect 16606 8206 16658 8258
rect 17166 8206 17218 8258
rect 17502 8206 17554 8258
rect 18286 8206 18338 8258
rect 18846 8206 18898 8258
rect 19518 8206 19570 8258
rect 22654 8206 22706 8258
rect 23550 8206 23602 8258
rect 26910 8206 26962 8258
rect 28366 8206 28418 8258
rect 28814 8206 28866 8258
rect 31390 8206 31442 8258
rect 31838 8206 31890 8258
rect 33182 8206 33234 8258
rect 36206 8206 36258 8258
rect 36766 8206 36818 8258
rect 37550 8206 37602 8258
rect 37774 8206 37826 8258
rect 43486 8206 43538 8258
rect 46286 8206 46338 8258
rect 46734 8206 46786 8258
rect 47406 8206 47458 8258
rect 48078 8206 48130 8258
rect 50766 8206 50818 8258
rect 55470 8206 55522 8258
rect 56702 8206 56754 8258
rect 57486 8206 57538 8258
rect 58382 8206 58434 8258
rect 59614 8206 59666 8258
rect 60286 8206 60338 8258
rect 62078 8206 62130 8258
rect 63310 8206 63362 8258
rect 63534 8206 63586 8258
rect 64990 8206 65042 8258
rect 66670 8206 66722 8258
rect 71150 8206 71202 8258
rect 71374 8206 71426 8258
rect 72046 8206 72098 8258
rect 72718 8206 72770 8258
rect 73166 8206 73218 8258
rect 73614 8206 73666 8258
rect 74622 8206 74674 8258
rect 74958 8206 75010 8258
rect 75518 8206 75570 8258
rect 75966 8206 76018 8258
rect 77310 8206 77362 8258
rect 77534 8206 77586 8258
rect 5854 8094 5906 8146
rect 10110 8094 10162 8146
rect 14254 8094 14306 8146
rect 19070 8094 19122 8146
rect 20190 8094 20242 8146
rect 26350 8094 26402 8146
rect 27022 8094 27074 8146
rect 27246 8094 27298 8146
rect 32286 8094 32338 8146
rect 38222 8094 38274 8146
rect 41582 8094 41634 8146
rect 43262 8094 43314 8146
rect 47630 8094 47682 8146
rect 48526 8094 48578 8146
rect 51886 8094 51938 8146
rect 62526 8094 62578 8146
rect 65326 8094 65378 8146
rect 66782 8094 66834 8146
rect 69806 8094 69858 8146
rect 70366 8094 70418 8146
rect 2494 7982 2546 8034
rect 3166 7982 3218 8034
rect 6190 7982 6242 8034
rect 6638 7982 6690 8034
rect 8206 7982 8258 8034
rect 9998 7982 10050 8034
rect 10670 7982 10722 8034
rect 11006 7982 11058 8034
rect 15822 7982 15874 8034
rect 17278 7982 17330 8034
rect 19966 7982 20018 8034
rect 21646 7982 21698 8034
rect 22206 7982 22258 8034
rect 22430 7982 22482 8034
rect 22542 7982 22594 8034
rect 24670 7982 24722 8034
rect 25118 7982 25170 8034
rect 29486 7982 29538 8034
rect 30718 7982 30770 8034
rect 37998 7982 38050 8034
rect 40686 7982 40738 8034
rect 48638 7982 48690 8034
rect 48862 7982 48914 8034
rect 49198 7982 49250 8034
rect 49646 7982 49698 8034
rect 50430 7982 50482 8034
rect 50654 7982 50706 8034
rect 51550 7982 51602 8034
rect 51774 7982 51826 8034
rect 52334 7982 52386 8034
rect 53342 7982 53394 8034
rect 53790 7982 53842 8034
rect 54238 7982 54290 8034
rect 56590 7982 56642 8034
rect 57374 7982 57426 8034
rect 57934 7982 57986 8034
rect 58830 7982 58882 8034
rect 64654 7982 64706 8034
rect 65214 7982 65266 8034
rect 67006 7982 67058 8034
rect 68014 7982 68066 8034
rect 68462 7982 68514 8034
rect 74174 7982 74226 8034
rect 74734 7982 74786 8034
rect 20534 7814 20586 7866
rect 20638 7814 20690 7866
rect 20742 7814 20794 7866
rect 39854 7814 39906 7866
rect 39958 7814 40010 7866
rect 40062 7814 40114 7866
rect 59174 7814 59226 7866
rect 59278 7814 59330 7866
rect 59382 7814 59434 7866
rect 78494 7814 78546 7866
rect 78598 7814 78650 7866
rect 78702 7814 78754 7866
rect 1822 7646 1874 7698
rect 2270 7646 2322 7698
rect 5518 7646 5570 7698
rect 6302 7646 6354 7698
rect 9886 7646 9938 7698
rect 10446 7646 10498 7698
rect 10894 7646 10946 7698
rect 12798 7646 12850 7698
rect 13582 7646 13634 7698
rect 13694 7646 13746 7698
rect 14590 7646 14642 7698
rect 14814 7646 14866 7698
rect 15374 7646 15426 7698
rect 15822 7646 15874 7698
rect 17614 7646 17666 7698
rect 23662 7646 23714 7698
rect 26686 7646 26738 7698
rect 27134 7646 27186 7698
rect 28702 7646 28754 7698
rect 28926 7646 28978 7698
rect 29598 7646 29650 7698
rect 29934 7646 29986 7698
rect 32734 7646 32786 7698
rect 40014 7646 40066 7698
rect 44382 7646 44434 7698
rect 48078 7646 48130 7698
rect 53566 7646 53618 7698
rect 59166 7646 59218 7698
rect 61070 7646 61122 7698
rect 63086 7646 63138 7698
rect 65550 7646 65602 7698
rect 65774 7646 65826 7698
rect 66558 7646 66610 7698
rect 67454 7646 67506 7698
rect 68462 7646 68514 7698
rect 69806 7646 69858 7698
rect 69918 7646 69970 7698
rect 73278 7646 73330 7698
rect 75518 7646 75570 7698
rect 2718 7534 2770 7586
rect 3054 7534 3106 7586
rect 6414 7534 6466 7586
rect 7870 7534 7922 7586
rect 9774 7534 9826 7586
rect 19182 7534 19234 7586
rect 23886 7534 23938 7586
rect 29038 7534 29090 7586
rect 31614 7534 31666 7586
rect 36542 7534 36594 7586
rect 48302 7534 48354 7586
rect 52446 7534 52498 7586
rect 56702 7534 56754 7586
rect 63310 7534 63362 7586
rect 68126 7534 68178 7586
rect 70590 7534 70642 7586
rect 75294 7534 75346 7586
rect 76974 7534 77026 7586
rect 77534 7534 77586 7586
rect 77870 7534 77922 7586
rect 4174 7422 4226 7474
rect 4510 7422 4562 7474
rect 5070 7422 5122 7474
rect 5630 7422 5682 7474
rect 5742 7422 5794 7474
rect 8430 7422 8482 7474
rect 13470 7422 13522 7474
rect 13806 7422 13858 7474
rect 14142 7422 14194 7474
rect 14926 7422 14978 7474
rect 18510 7422 18562 7474
rect 19070 7422 19122 7474
rect 22766 7422 22818 7474
rect 23998 7422 24050 7474
rect 28030 7422 28082 7474
rect 31502 7422 31554 7474
rect 31838 7422 31890 7474
rect 32174 7422 32226 7474
rect 32622 7422 32674 7474
rect 32846 7422 32898 7474
rect 37774 7422 37826 7474
rect 39902 7422 39954 7474
rect 40126 7422 40178 7474
rect 40574 7422 40626 7474
rect 44270 7422 44322 7474
rect 44494 7422 44546 7474
rect 44942 7422 44994 7474
rect 47406 7422 47458 7474
rect 48414 7422 48466 7474
rect 49870 7422 49922 7474
rect 51102 7422 51154 7474
rect 52670 7422 52722 7474
rect 52894 7422 52946 7474
rect 53006 7422 53058 7474
rect 54574 7422 54626 7474
rect 56142 7422 56194 7474
rect 62638 7422 62690 7474
rect 65438 7422 65490 7474
rect 66110 7422 66162 7474
rect 67342 7422 67394 7474
rect 67678 7422 67730 7474
rect 69358 7422 69410 7474
rect 70030 7422 70082 7474
rect 71710 7422 71762 7474
rect 75182 7422 75234 7474
rect 76302 7422 76354 7474
rect 76862 7422 76914 7474
rect 4622 7310 4674 7362
rect 8654 7310 8706 7362
rect 16270 7310 16322 7362
rect 16830 7310 16882 7362
rect 22318 7310 22370 7362
rect 24782 7310 24834 7362
rect 25566 7310 25618 7362
rect 26014 7310 26066 7362
rect 28254 7310 28306 7362
rect 30942 7310 30994 7362
rect 36318 7310 36370 7362
rect 38446 7310 38498 7362
rect 39342 7310 39394 7362
rect 45390 7310 45442 7362
rect 46622 7310 46674 7362
rect 47294 7310 47346 7362
rect 50094 7310 50146 7362
rect 52782 7310 52834 7362
rect 54686 7310 54738 7362
rect 57374 7310 57426 7362
rect 57822 7310 57874 7362
rect 58382 7310 58434 7362
rect 58718 7310 58770 7362
rect 59726 7310 59778 7362
rect 60062 7310 60114 7362
rect 60510 7310 60562 7362
rect 61406 7310 61458 7362
rect 61854 7310 61906 7362
rect 63198 7310 63250 7362
rect 63870 7310 63922 7362
rect 64318 7310 64370 7362
rect 64654 7310 64706 7362
rect 69582 7310 69634 7362
rect 71822 7310 71874 7362
rect 73838 7310 73890 7362
rect 74174 7310 74226 7362
rect 74734 7310 74786 7362
rect 9886 7198 9938 7250
rect 22654 7198 22706 7250
rect 27694 7198 27746 7250
rect 51326 7198 51378 7250
rect 57934 7198 57986 7250
rect 58718 7198 58770 7250
rect 60510 7198 60562 7250
rect 61854 7198 61906 7250
rect 63982 7198 64034 7250
rect 64654 7198 64706 7250
rect 68014 7198 68066 7250
rect 68462 7198 68514 7250
rect 72270 7198 72322 7250
rect 73838 7198 73890 7250
rect 74174 7198 74226 7250
rect 10874 7030 10926 7082
rect 10978 7030 11030 7082
rect 11082 7030 11134 7082
rect 30194 7030 30246 7082
rect 30298 7030 30350 7082
rect 30402 7030 30454 7082
rect 49514 7030 49566 7082
rect 49618 7030 49670 7082
rect 49722 7030 49774 7082
rect 68834 7030 68886 7082
rect 68938 7030 68990 7082
rect 69042 7030 69094 7082
rect 18958 6862 19010 6914
rect 32510 6862 32562 6914
rect 35534 6862 35586 6914
rect 39902 6862 39954 6914
rect 50094 6862 50146 6914
rect 50878 6862 50930 6914
rect 54686 6862 54738 6914
rect 55358 6862 55410 6914
rect 66446 6862 66498 6914
rect 8430 6750 8482 6802
rect 13694 6750 13746 6802
rect 15038 6750 15090 6802
rect 22206 6750 22258 6802
rect 27806 6750 27858 6802
rect 29486 6750 29538 6802
rect 32062 6750 32114 6802
rect 43486 6750 43538 6802
rect 49534 6750 49586 6802
rect 55918 6750 55970 6802
rect 60622 6750 60674 6802
rect 62190 6750 62242 6802
rect 65774 6750 65826 6802
rect 3054 6638 3106 6690
rect 4734 6638 4786 6690
rect 9326 6638 9378 6690
rect 9662 6638 9714 6690
rect 10446 6638 10498 6690
rect 10894 6638 10946 6690
rect 12574 6638 12626 6690
rect 12910 6638 12962 6690
rect 13918 6638 13970 6690
rect 14142 6638 14194 6690
rect 15598 6638 15650 6690
rect 16606 6638 16658 6690
rect 17726 6638 17778 6690
rect 18062 6638 18114 6690
rect 19070 6638 19122 6690
rect 19966 6638 20018 6690
rect 21982 6638 22034 6690
rect 22654 6638 22706 6690
rect 23998 6638 24050 6690
rect 24334 6638 24386 6690
rect 26350 6638 26402 6690
rect 27134 6638 27186 6690
rect 27582 6638 27634 6690
rect 28254 6638 28306 6690
rect 31166 6638 31218 6690
rect 32398 6638 32450 6690
rect 34974 6638 35026 6690
rect 35310 6638 35362 6690
rect 39678 6638 39730 6690
rect 40350 6638 40402 6690
rect 41022 6638 41074 6690
rect 41358 6638 41410 6690
rect 42590 6638 42642 6690
rect 43038 6638 43090 6690
rect 45950 6638 46002 6690
rect 51214 6638 51266 6690
rect 51550 6638 51602 6690
rect 52558 6638 52610 6690
rect 54574 6638 54626 6690
rect 55582 6638 55634 6690
rect 55806 6638 55858 6690
rect 56030 6638 56082 6690
rect 59726 6638 59778 6690
rect 61294 6638 61346 6690
rect 62078 6638 62130 6690
rect 62974 6638 63026 6690
rect 64766 6638 64818 6690
rect 65662 6638 65714 6690
rect 67790 6638 67842 6690
rect 68014 6638 68066 6690
rect 68350 6638 68402 6690
rect 70030 6638 70082 6690
rect 70926 6638 70978 6690
rect 72158 6638 72210 6690
rect 72606 6638 72658 6690
rect 73166 6638 73218 6690
rect 76078 6638 76130 6690
rect 77422 6638 77474 6690
rect 1934 6526 1986 6578
rect 4398 6526 4450 6578
rect 24110 6526 24162 6578
rect 25230 6526 25282 6578
rect 26798 6526 26850 6578
rect 28142 6526 28194 6578
rect 31054 6526 31106 6578
rect 34862 6526 34914 6578
rect 36094 6526 36146 6578
rect 36430 6526 36482 6578
rect 49982 6526 50034 6578
rect 51438 6526 51490 6578
rect 56702 6526 56754 6578
rect 56814 6526 56866 6578
rect 59166 6526 59218 6578
rect 64430 6526 64482 6578
rect 69694 6526 69746 6578
rect 75070 6526 75122 6578
rect 77310 6526 77362 6578
rect 3726 6414 3778 6466
rect 4510 6414 4562 6466
rect 5630 6414 5682 6466
rect 6078 6414 6130 6466
rect 8878 6414 8930 6466
rect 9550 6414 9602 6466
rect 10110 6414 10162 6466
rect 10334 6414 10386 6466
rect 11342 6414 11394 6466
rect 12014 6414 12066 6466
rect 12686 6414 12738 6466
rect 14254 6414 14306 6466
rect 14366 6414 14418 6466
rect 16270 6414 16322 6466
rect 16494 6414 16546 6466
rect 23214 6414 23266 6466
rect 23774 6414 23826 6466
rect 23886 6414 23938 6466
rect 24894 6414 24946 6466
rect 25118 6414 25170 6466
rect 25790 6414 25842 6466
rect 26910 6414 26962 6466
rect 28030 6414 28082 6466
rect 28814 6414 28866 6466
rect 30046 6414 30098 6466
rect 30606 6414 30658 6466
rect 34190 6414 34242 6466
rect 35086 6414 35138 6466
rect 36206 6414 36258 6466
rect 36766 6414 36818 6466
rect 37438 6414 37490 6466
rect 37886 6414 37938 6466
rect 41246 6414 41298 6466
rect 42142 6414 42194 6466
rect 44382 6414 44434 6466
rect 44718 6414 44770 6466
rect 45390 6414 45442 6466
rect 46510 6414 46562 6466
rect 47070 6414 47122 6466
rect 47406 6414 47458 6466
rect 47854 6414 47906 6466
rect 48302 6414 48354 6466
rect 48750 6414 48802 6466
rect 50094 6414 50146 6466
rect 51326 6414 51378 6466
rect 52110 6414 52162 6466
rect 53342 6414 53394 6466
rect 53902 6414 53954 6466
rect 54686 6414 54738 6466
rect 57038 6414 57090 6466
rect 57374 6414 57426 6466
rect 57822 6414 57874 6466
rect 58382 6414 58434 6466
rect 60174 6414 60226 6466
rect 63422 6414 63474 6466
rect 63870 6414 63922 6466
rect 64542 6414 64594 6466
rect 67006 6414 67058 6466
rect 67678 6414 67730 6466
rect 67902 6414 67954 6466
rect 71486 6414 71538 6466
rect 72494 6414 72546 6466
rect 72718 6414 72770 6466
rect 73614 6414 73666 6466
rect 74062 6414 74114 6466
rect 77534 6414 77586 6466
rect 77758 6414 77810 6466
rect 20534 6246 20586 6298
rect 20638 6246 20690 6298
rect 20742 6246 20794 6298
rect 39854 6246 39906 6298
rect 39958 6246 40010 6298
rect 40062 6246 40114 6298
rect 59174 6246 59226 6298
rect 59278 6246 59330 6298
rect 59382 6246 59434 6298
rect 78494 6246 78546 6298
rect 78598 6246 78650 6298
rect 78702 6246 78754 6298
rect 2494 6078 2546 6130
rect 10222 6078 10274 6130
rect 10446 6078 10498 6130
rect 11118 6078 11170 6130
rect 15486 6078 15538 6130
rect 16046 6078 16098 6130
rect 16830 6078 16882 6130
rect 22094 6078 22146 6130
rect 23326 6078 23378 6130
rect 35422 6078 35474 6130
rect 37326 6078 37378 6130
rect 45950 6078 46002 6130
rect 46174 6078 46226 6130
rect 48526 6078 48578 6130
rect 48638 6078 48690 6130
rect 51662 6078 51714 6130
rect 52446 6078 52498 6130
rect 53342 6078 53394 6130
rect 55806 6078 55858 6130
rect 56030 6078 56082 6130
rect 58942 6078 58994 6130
rect 59054 6078 59106 6130
rect 62638 6078 62690 6130
rect 62862 6078 62914 6130
rect 66670 6078 66722 6130
rect 67566 6078 67618 6130
rect 68574 6078 68626 6130
rect 69806 6078 69858 6130
rect 70254 6078 70306 6130
rect 70702 6078 70754 6130
rect 73278 6078 73330 6130
rect 74286 6078 74338 6130
rect 74510 6078 74562 6130
rect 77982 6078 78034 6130
rect 4622 5966 4674 6018
rect 7422 5966 7474 6018
rect 12798 5966 12850 6018
rect 16158 5966 16210 6018
rect 18510 5966 18562 6018
rect 21758 5966 21810 6018
rect 36318 5966 36370 6018
rect 36542 5966 36594 6018
rect 39118 5966 39170 6018
rect 49646 5966 49698 6018
rect 49758 5966 49810 6018
rect 51438 5966 51490 6018
rect 57710 5966 57762 6018
rect 57822 5966 57874 6018
rect 62190 5966 62242 6018
rect 62974 5966 63026 6018
rect 63646 5966 63698 6018
rect 63758 5966 63810 6018
rect 66558 5966 66610 6018
rect 68798 5966 68850 6018
rect 68910 5966 68962 6018
rect 75966 5966 76018 6018
rect 76526 5966 76578 6018
rect 3502 5854 3554 5906
rect 3838 5854 3890 5906
rect 5406 5854 5458 5906
rect 6750 5854 6802 5906
rect 8430 5854 8482 5906
rect 8654 5854 8706 5906
rect 13134 5854 13186 5906
rect 14030 5854 14082 5906
rect 15822 5854 15874 5906
rect 18286 5854 18338 5906
rect 18622 5854 18674 5906
rect 21982 5854 22034 5906
rect 22206 5854 22258 5906
rect 22878 5854 22930 5906
rect 23214 5854 23266 5906
rect 23550 5854 23602 5906
rect 24446 5854 24498 5906
rect 27134 5854 27186 5906
rect 28142 5854 28194 5906
rect 28814 5854 28866 5906
rect 30046 5854 30098 5906
rect 30942 5854 30994 5906
rect 32062 5854 32114 5906
rect 32510 5854 32562 5906
rect 32734 5854 32786 5906
rect 35086 5854 35138 5906
rect 36206 5854 36258 5906
rect 38670 5854 38722 5906
rect 39566 5854 39618 5906
rect 40798 5854 40850 5906
rect 42142 5854 42194 5906
rect 42590 5854 42642 5906
rect 44942 5854 44994 5906
rect 45838 5854 45890 5906
rect 46286 5854 46338 5906
rect 48414 5854 48466 5906
rect 51326 5854 51378 5906
rect 51998 5854 52050 5906
rect 54910 5854 54962 5906
rect 55582 5854 55634 5906
rect 55918 5854 55970 5906
rect 56142 5854 56194 5906
rect 58046 5854 58098 5906
rect 58830 5854 58882 5906
rect 59166 5854 59218 5906
rect 60062 5854 60114 5906
rect 61518 5854 61570 5906
rect 65886 5854 65938 5906
rect 66894 5854 66946 5906
rect 67902 5854 67954 5906
rect 68126 5854 68178 5906
rect 72046 5854 72098 5906
rect 72382 5854 72434 5906
rect 74174 5854 74226 5906
rect 75294 5854 75346 5906
rect 76974 5854 77026 5906
rect 6638 5742 6690 5794
rect 8990 5742 9042 5794
rect 9998 5742 10050 5794
rect 10334 5742 10386 5794
rect 11566 5742 11618 5794
rect 12014 5742 12066 5794
rect 14702 5742 14754 5794
rect 17614 5742 17666 5794
rect 19070 5742 19122 5794
rect 19518 5742 19570 5794
rect 19966 5742 20018 5794
rect 23438 5742 23490 5794
rect 24894 5742 24946 5794
rect 25678 5742 25730 5794
rect 26238 5742 26290 5794
rect 26686 5742 26738 5794
rect 30382 5742 30434 5794
rect 33854 5742 33906 5794
rect 34414 5742 34466 5794
rect 34862 5742 34914 5794
rect 36878 5742 36930 5794
rect 37774 5742 37826 5794
rect 39454 5742 39506 5794
rect 41694 5742 41746 5794
rect 43150 5742 43202 5794
rect 43486 5742 43538 5794
rect 44158 5742 44210 5794
rect 44830 5742 44882 5794
rect 46062 5742 46114 5794
rect 46846 5742 46898 5794
rect 47294 5742 47346 5794
rect 48190 5742 48242 5794
rect 50206 5742 50258 5794
rect 50654 5742 50706 5794
rect 52894 5742 52946 5794
rect 53790 5742 53842 5794
rect 54462 5742 54514 5794
rect 56702 5742 56754 5794
rect 58494 5742 58546 5794
rect 59950 5742 60002 5794
rect 64206 5742 64258 5794
rect 64654 5742 64706 5794
rect 65550 5742 65602 5794
rect 69358 5742 69410 5794
rect 72606 5742 72658 5794
rect 75070 5742 75122 5794
rect 77310 5742 77362 5794
rect 3614 5630 3666 5682
rect 9774 5630 9826 5682
rect 25566 5630 25618 5682
rect 26462 5630 26514 5682
rect 47966 5630 48018 5682
rect 49646 5630 49698 5682
rect 63646 5630 63698 5682
rect 10874 5462 10926 5514
rect 10978 5462 11030 5514
rect 11082 5462 11134 5514
rect 30194 5462 30246 5514
rect 30298 5462 30350 5514
rect 30402 5462 30454 5514
rect 49514 5462 49566 5514
rect 49618 5462 49670 5514
rect 49722 5462 49774 5514
rect 68834 5462 68886 5514
rect 68938 5462 68990 5514
rect 69042 5462 69094 5514
rect 8654 5294 8706 5346
rect 13694 5294 13746 5346
rect 14030 5294 14082 5346
rect 22206 5294 22258 5346
rect 25454 5294 25506 5346
rect 27470 5294 27522 5346
rect 28814 5294 28866 5346
rect 39790 5294 39842 5346
rect 46398 5294 46450 5346
rect 49198 5294 49250 5346
rect 53566 5294 53618 5346
rect 56590 5294 56642 5346
rect 59054 5294 59106 5346
rect 59278 5294 59330 5346
rect 60174 5294 60226 5346
rect 72494 5294 72546 5346
rect 76302 5294 76354 5346
rect 4510 5182 4562 5234
rect 7646 5182 7698 5234
rect 7982 5182 8034 5234
rect 9326 5182 9378 5234
rect 9886 5182 9938 5234
rect 10558 5182 10610 5234
rect 13022 5182 13074 5234
rect 14254 5182 14306 5234
rect 14926 5182 14978 5234
rect 21982 5182 22034 5234
rect 27470 5182 27522 5234
rect 27918 5182 27970 5234
rect 32286 5182 32338 5234
rect 34078 5182 34130 5234
rect 39118 5182 39170 5234
rect 42478 5182 42530 5234
rect 42926 5182 42978 5234
rect 47742 5182 47794 5234
rect 50430 5182 50482 5234
rect 57598 5182 57650 5234
rect 59278 5182 59330 5234
rect 61966 5182 62018 5234
rect 64318 5182 64370 5234
rect 64878 5182 64930 5234
rect 69246 5182 69298 5234
rect 69694 5182 69746 5234
rect 70590 5182 70642 5234
rect 71710 5182 71762 5234
rect 73502 5182 73554 5234
rect 75630 5182 75682 5234
rect 77198 5182 77250 5234
rect 2942 5070 2994 5122
rect 3838 5070 3890 5122
rect 4846 5070 4898 5122
rect 10670 5070 10722 5122
rect 12126 5070 12178 5122
rect 15150 5070 15202 5122
rect 17054 5070 17106 5122
rect 17502 5070 17554 5122
rect 18846 5070 18898 5122
rect 19182 5070 19234 5122
rect 20526 5070 20578 5122
rect 22542 5070 22594 5122
rect 23886 5070 23938 5122
rect 24558 5070 24610 5122
rect 25566 5070 25618 5122
rect 26462 5070 26514 5122
rect 28366 5070 28418 5122
rect 28926 5070 28978 5122
rect 29710 5070 29762 5122
rect 30046 5070 30098 5122
rect 30494 5070 30546 5122
rect 33518 5070 33570 5122
rect 35198 5070 35250 5122
rect 38110 5070 38162 5122
rect 38558 5070 38610 5122
rect 40126 5070 40178 5122
rect 41022 5070 41074 5122
rect 41470 5070 41522 5122
rect 43374 5070 43426 5122
rect 44494 5070 44546 5122
rect 45390 5070 45442 5122
rect 47630 5070 47682 5122
rect 49310 5070 49362 5122
rect 51102 5070 51154 5122
rect 51774 5070 51826 5122
rect 52110 5070 52162 5122
rect 55358 5070 55410 5122
rect 57150 5070 57202 5122
rect 60734 5070 60786 5122
rect 62526 5070 62578 5122
rect 63422 5070 63474 5122
rect 65774 5070 65826 5122
rect 66558 5070 66610 5122
rect 67678 5070 67730 5122
rect 67902 5070 67954 5122
rect 70254 5070 70306 5122
rect 72046 5070 72098 5122
rect 73950 5070 74002 5122
rect 75518 5070 75570 5122
rect 77646 5070 77698 5122
rect 78094 5070 78146 5122
rect 1934 4958 1986 5010
rect 8654 4958 8706 5010
rect 8766 4958 8818 5010
rect 11342 4958 11394 5010
rect 16494 4958 16546 5010
rect 16606 4958 16658 5010
rect 18510 4958 18562 5010
rect 29822 4958 29874 5010
rect 30830 4958 30882 5010
rect 32958 4958 33010 5010
rect 34862 4958 34914 5010
rect 36542 4958 36594 5010
rect 36766 4958 36818 5010
rect 39006 4958 39058 5010
rect 40462 4958 40514 5010
rect 44718 4958 44770 5010
rect 45614 4958 45666 5010
rect 45726 4958 45778 5010
rect 46510 4958 46562 5010
rect 53678 4958 53730 5010
rect 54798 4958 54850 5010
rect 56590 4958 56642 5010
rect 56702 4958 56754 5010
rect 58606 4958 58658 5010
rect 60398 4958 60450 5010
rect 60510 4958 60562 5010
rect 63086 4958 63138 5010
rect 65438 4958 65490 5010
rect 65550 4958 65602 5010
rect 66222 4958 66274 5010
rect 68238 4958 68290 5010
rect 3614 4846 3666 4898
rect 11790 4846 11842 4898
rect 12014 4846 12066 4898
rect 15486 4846 15538 4898
rect 16270 4846 16322 4898
rect 17950 4846 18002 4898
rect 18622 4846 18674 4898
rect 19854 4846 19906 4898
rect 19966 4846 20018 4898
rect 20078 4846 20130 4898
rect 20974 4846 21026 4898
rect 27022 4846 27074 4898
rect 30718 4846 30770 4898
rect 31278 4846 31330 4898
rect 31950 4846 32002 4898
rect 32846 4846 32898 4898
rect 33070 4846 33122 4898
rect 37774 4846 37826 4898
rect 39230 4846 39282 4898
rect 40238 4846 40290 4898
rect 40350 4846 40402 4898
rect 41918 4846 41970 4898
rect 44158 4846 44210 4898
rect 44270 4846 44322 4898
rect 44382 4846 44434 4898
rect 46398 4846 46450 4898
rect 53566 4846 53618 4898
rect 54462 4846 54514 4898
rect 54686 4846 54738 4898
rect 55918 4846 55970 4898
rect 58046 4846 58098 4898
rect 58718 4846 58770 4898
rect 58942 4846 58994 4898
rect 59726 4846 59778 4898
rect 61294 4846 61346 4898
rect 63198 4846 63250 4898
rect 63870 4846 63922 4898
rect 66334 4846 66386 4898
rect 66894 4846 66946 4898
rect 68126 4846 68178 4898
rect 68350 4846 68402 4898
rect 73054 4846 73106 4898
rect 74398 4846 74450 4898
rect 20534 4678 20586 4730
rect 20638 4678 20690 4730
rect 20742 4678 20794 4730
rect 39854 4678 39906 4730
rect 39958 4678 40010 4730
rect 40062 4678 40114 4730
rect 59174 4678 59226 4730
rect 59278 4678 59330 4730
rect 59382 4678 59434 4730
rect 78494 4678 78546 4730
rect 78598 4678 78650 4730
rect 78702 4678 78754 4730
rect 3614 4510 3666 4562
rect 13806 4510 13858 4562
rect 16382 4510 16434 4562
rect 17054 4510 17106 4562
rect 21086 4510 21138 4562
rect 22094 4510 22146 4562
rect 23438 4510 23490 4562
rect 23774 4510 23826 4562
rect 24558 4510 24610 4562
rect 26126 4510 26178 4562
rect 26350 4510 26402 4562
rect 27246 4510 27298 4562
rect 31278 4510 31330 4562
rect 35534 4510 35586 4562
rect 37886 4510 37938 4562
rect 38110 4510 38162 4562
rect 41694 4510 41746 4562
rect 41918 4510 41970 4562
rect 42702 4510 42754 4562
rect 46958 4510 47010 4562
rect 47518 4510 47570 4562
rect 48414 4510 48466 4562
rect 48638 4510 48690 4562
rect 50542 4510 50594 4562
rect 53006 4510 53058 4562
rect 53678 4510 53730 4562
rect 56478 4510 56530 4562
rect 57934 4510 57986 4562
rect 59614 4510 59666 4562
rect 61518 4510 61570 4562
rect 64430 4510 64482 4562
rect 3950 4398 4002 4450
rect 4510 4398 4562 4450
rect 9886 4398 9938 4450
rect 10558 4398 10610 4450
rect 12798 4398 12850 4450
rect 14814 4398 14866 4450
rect 16270 4398 16322 4450
rect 21310 4398 21362 4450
rect 21982 4398 22034 4450
rect 23998 4398 24050 4450
rect 24110 4398 24162 4450
rect 24782 4398 24834 4450
rect 24894 4398 24946 4450
rect 27694 4398 27746 4450
rect 32846 4398 32898 4450
rect 35646 4398 35698 4450
rect 40350 4398 40402 4450
rect 40462 4398 40514 4450
rect 42030 4398 42082 4450
rect 42254 4398 42306 4450
rect 43486 4398 43538 4450
rect 47406 4398 47458 4450
rect 49758 4398 49810 4450
rect 50094 4398 50146 4450
rect 50766 4398 50818 4450
rect 51550 4398 51602 4450
rect 51662 4398 51714 4450
rect 54798 4398 54850 4450
rect 57710 4398 57762 4450
rect 58942 4398 58994 4450
rect 59054 4398 59106 4450
rect 59838 4398 59890 4450
rect 59950 4398 60002 4450
rect 60398 4398 60450 4450
rect 63534 4398 63586 4450
rect 68238 4398 68290 4450
rect 71374 4398 71426 4450
rect 71934 4454 71986 4506
rect 72606 4510 72658 4562
rect 73278 4510 73330 4562
rect 74062 4510 74114 4562
rect 72046 4398 72098 4450
rect 76750 4398 76802 4450
rect 77086 4398 77138 4450
rect 77646 4398 77698 4450
rect 77982 4398 78034 4450
rect 3054 4286 3106 4338
rect 8654 4286 8706 4338
rect 11454 4286 11506 4338
rect 12238 4286 12290 4338
rect 14926 4286 14978 4338
rect 17950 4286 18002 4338
rect 20414 4286 20466 4338
rect 21422 4286 21474 4338
rect 25678 4286 25730 4338
rect 26014 4286 26066 4338
rect 27022 4286 27074 4338
rect 27358 4286 27410 4338
rect 27470 4286 27522 4338
rect 29150 4286 29202 4338
rect 30158 4286 30210 4338
rect 32174 4286 32226 4338
rect 32734 4286 32786 4338
rect 33630 4286 33682 4338
rect 34078 4286 34130 4338
rect 35310 4286 35362 4338
rect 36766 4286 36818 4338
rect 37774 4286 37826 4338
rect 39454 4286 39506 4338
rect 41806 4286 41858 4338
rect 48750 4286 48802 4338
rect 50878 4286 50930 4338
rect 51326 4286 51378 4338
rect 52446 4286 52498 4338
rect 55134 4286 55186 4338
rect 56142 4286 56194 4338
rect 58046 4286 58098 4338
rect 58158 4286 58210 4338
rect 58382 4286 58434 4338
rect 61294 4286 61346 4338
rect 61630 4286 61682 4338
rect 61966 4286 62018 4338
rect 65662 4286 65714 4338
rect 67006 4286 67058 4338
rect 69582 4286 69634 4338
rect 70926 4286 70978 4338
rect 74398 4286 74450 4338
rect 76190 4286 76242 4338
rect 1934 4174 1986 4226
rect 9102 4174 9154 4226
rect 11118 4174 11170 4226
rect 13358 4174 13410 4226
rect 18286 4174 18338 4226
rect 18958 4174 19010 4226
rect 20302 4174 20354 4226
rect 22878 4174 22930 4226
rect 26238 4174 26290 4226
rect 30606 4174 30658 4226
rect 34414 4174 34466 4226
rect 36206 4174 36258 4226
rect 37102 4174 37154 4226
rect 38670 4174 38722 4226
rect 38894 4174 38946 4226
rect 54126 4174 54178 4226
rect 55582 4174 55634 4226
rect 61406 4174 61458 4226
rect 62526 4174 62578 4226
rect 65886 4174 65938 4226
rect 69134 4174 69186 4226
rect 75518 4174 75570 4226
rect 9998 4062 10050 4114
rect 20078 4062 20130 4114
rect 22094 4062 22146 4114
rect 28478 4062 28530 4114
rect 40350 4062 40402 4114
rect 47518 4062 47570 4114
rect 59054 4062 59106 4114
rect 67678 4062 67730 4114
rect 72046 4062 72098 4114
rect 10874 3894 10926 3946
rect 10978 3894 11030 3946
rect 11082 3894 11134 3946
rect 30194 3894 30246 3946
rect 30298 3894 30350 3946
rect 30402 3894 30454 3946
rect 49514 3894 49566 3946
rect 49618 3894 49670 3946
rect 49722 3894 49774 3946
rect 68834 3894 68886 3946
rect 68938 3894 68990 3946
rect 69042 3894 69094 3946
rect 34190 3726 34242 3778
rect 42926 3726 42978 3778
rect 59614 3726 59666 3778
rect 67342 3726 67394 3778
rect 67678 3726 67730 3778
rect 4958 3614 5010 3666
rect 7198 3614 7250 3666
rect 10334 3614 10386 3666
rect 14030 3614 14082 3666
rect 15486 3614 15538 3666
rect 18510 3614 18562 3666
rect 20078 3614 20130 3666
rect 20526 3614 20578 3666
rect 21646 3614 21698 3666
rect 22654 3614 22706 3666
rect 24110 3614 24162 3666
rect 25454 3614 25506 3666
rect 27246 3614 27298 3666
rect 27694 3614 27746 3666
rect 28142 3614 28194 3666
rect 30158 3614 30210 3666
rect 31950 3614 32002 3666
rect 38670 3614 38722 3666
rect 45166 3614 45218 3666
rect 45502 3614 45554 3666
rect 46846 3614 46898 3666
rect 47406 3614 47458 3666
rect 53342 3614 53394 3666
rect 53902 3614 53954 3666
rect 55022 3614 55074 3666
rect 63534 3614 63586 3666
rect 65102 3614 65154 3666
rect 67118 3614 67170 3666
rect 68910 3614 68962 3666
rect 72382 3614 72434 3666
rect 74846 3614 74898 3666
rect 76302 3614 76354 3666
rect 77310 3614 77362 3666
rect 2158 3502 2210 3554
rect 5630 3502 5682 3554
rect 9662 3502 9714 3554
rect 11454 3502 11506 3554
rect 11678 3502 11730 3554
rect 13582 3502 13634 3554
rect 15262 3502 15314 3554
rect 15710 3502 15762 3554
rect 16606 3502 16658 3554
rect 17502 3502 17554 3554
rect 17950 3502 18002 3554
rect 18846 3502 18898 3554
rect 19854 3502 19906 3554
rect 22094 3502 22146 3554
rect 24558 3502 24610 3554
rect 25902 3502 25954 3554
rect 29262 3502 29314 3554
rect 32510 3502 32562 3554
rect 34302 3502 34354 3554
rect 34862 3502 34914 3554
rect 35982 3502 36034 3554
rect 37102 3502 37154 3554
rect 38222 3502 38274 3554
rect 39118 3502 39170 3554
rect 39902 3502 39954 3554
rect 40238 3502 40290 3554
rect 42814 3502 42866 3554
rect 43598 3502 43650 3554
rect 44046 3502 44098 3554
rect 44942 3502 44994 3554
rect 45390 3502 45442 3554
rect 52782 3502 52834 3554
rect 54462 3502 54514 3554
rect 55470 3502 55522 3554
rect 56926 3502 56978 3554
rect 57486 3502 57538 3554
rect 59502 3502 59554 3554
rect 64766 3502 64818 3554
rect 66558 3502 66610 3554
rect 68350 3502 68402 3554
rect 73390 3502 73442 3554
rect 75518 3502 75570 3554
rect 76750 3502 76802 3554
rect 2830 3390 2882 3442
rect 6750 3390 6802 3442
rect 8206 3390 8258 3442
rect 11566 3390 11618 3442
rect 11902 3390 11954 3442
rect 12910 3390 12962 3442
rect 15038 3390 15090 3442
rect 23550 3390 23602 3442
rect 26350 3390 26402 3442
rect 28590 3390 28642 3442
rect 30606 3390 30658 3442
rect 30942 3390 30994 3442
rect 31614 3390 31666 3442
rect 33182 3390 33234 3442
rect 34190 3390 34242 3442
rect 36430 3390 36482 3442
rect 39454 3390 39506 3442
rect 41246 3390 41298 3442
rect 42030 3390 42082 3442
rect 46286 3390 46338 3442
rect 47966 3390 48018 3442
rect 48750 3390 48802 3442
rect 50990 3390 51042 3442
rect 51774 3390 51826 3442
rect 58046 3390 58098 3442
rect 58606 3390 58658 3442
rect 58942 3390 58994 3442
rect 62974 3390 63026 3442
rect 65662 3390 65714 3442
rect 66222 3390 66274 3442
rect 70254 3390 70306 3442
rect 71374 3390 71426 3442
rect 77758 3390 77810 3442
rect 15150 3278 15202 3330
rect 16270 3278 16322 3330
rect 26686 3278 26738 3330
rect 29598 3278 29650 3330
rect 33518 3278 33570 3330
rect 35198 3278 35250 3330
rect 37438 3278 37490 3330
rect 40126 3278 40178 3330
rect 41582 3278 41634 3330
rect 42926 3278 42978 3330
rect 45614 3278 45666 3330
rect 56590 3278 56642 3330
rect 56814 3278 56866 3330
rect 59614 3278 59666 3330
rect 60510 3278 60562 3330
rect 71038 3278 71090 3330
rect 73166 3278 73218 3330
rect 20534 3110 20586 3162
rect 20638 3110 20690 3162
rect 20742 3110 20794 3162
rect 39854 3110 39906 3162
rect 39958 3110 40010 3162
rect 40062 3110 40114 3162
rect 59174 3110 59226 3162
rect 59278 3110 59330 3162
rect 59382 3110 59434 3162
rect 78494 3110 78546 3162
rect 78598 3110 78650 3162
rect 78702 3110 78754 3162
<< metal2 >>
rect 1680 39200 1792 40000
rect 4144 39200 4256 40000
rect 6608 39200 6720 40000
rect 9072 39200 9184 40000
rect 9436 39228 9828 39284
rect 1708 37940 1764 39200
rect 2156 38500 2212 38510
rect 1708 37884 2100 37940
rect 2044 36594 2100 37884
rect 2044 36542 2046 36594
rect 2098 36542 2100 36594
rect 2044 36530 2100 36542
rect 1932 36036 1988 36046
rect 1932 35810 1988 35980
rect 1932 35758 1934 35810
rect 1986 35758 1988 35810
rect 1932 35746 1988 35758
rect 2156 35026 2212 38444
rect 2492 37716 2548 37726
rect 2156 34974 2158 35026
rect 2210 34974 2212 35026
rect 2156 34962 2212 34974
rect 2268 37492 2324 37502
rect 1932 34018 1988 34030
rect 1932 33966 1934 34018
rect 1986 33966 1988 34018
rect 1932 33572 1988 33966
rect 1932 33506 1988 33516
rect 1932 31666 1988 31678
rect 1932 31614 1934 31666
rect 1986 31614 1988 31666
rect 1596 31220 1652 31230
rect 1484 29764 1540 29774
rect 1372 25732 1428 25742
rect 1372 7588 1428 25676
rect 1372 7522 1428 7532
rect 1484 5124 1540 29708
rect 1484 5058 1540 5068
rect 1596 4452 1652 31164
rect 1932 31108 1988 31614
rect 1932 31042 1988 31052
rect 1932 29314 1988 29326
rect 1932 29262 1934 29314
rect 1986 29262 1988 29314
rect 1932 28644 1988 29262
rect 1932 28578 1988 28588
rect 1932 26180 1988 26190
rect 1932 26086 1988 26124
rect 1932 23826 1988 23838
rect 1932 23774 1934 23826
rect 1986 23774 1988 23826
rect 1932 23716 1988 23774
rect 1932 23650 1988 23660
rect 2156 22146 2212 22158
rect 2156 22094 2158 22146
rect 2210 22094 2212 22146
rect 2044 21812 2100 21822
rect 2044 21476 2100 21756
rect 2156 21700 2212 22094
rect 2156 21634 2212 21644
rect 2156 21476 2212 21486
rect 2044 21474 2212 21476
rect 2044 21422 2158 21474
rect 2210 21422 2212 21474
rect 2044 21420 2212 21422
rect 2156 21410 2212 21420
rect 1932 21252 1988 21262
rect 1932 20914 1988 21196
rect 1932 20862 1934 20914
rect 1986 20862 1988 20914
rect 1932 20850 1988 20862
rect 2268 20188 2324 37436
rect 2380 29988 2436 29998
rect 2380 29894 2436 29932
rect 2492 26068 2548 37660
rect 4172 36594 4228 39200
rect 4172 36542 4174 36594
rect 4226 36542 4228 36594
rect 4172 36530 4228 36542
rect 5068 37156 5124 37166
rect 3164 36484 3220 36494
rect 3164 36390 3220 36428
rect 4956 36482 5012 36494
rect 4956 36430 4958 36482
rect 5010 36430 5012 36482
rect 4956 35924 5012 36430
rect 4956 35858 5012 35868
rect 3052 35812 3108 35822
rect 3052 35698 3108 35756
rect 3612 35812 3668 35822
rect 3612 35718 3668 35756
rect 4508 35810 4564 35822
rect 4508 35758 4510 35810
rect 4562 35758 4564 35810
rect 3052 35646 3054 35698
rect 3106 35646 3108 35698
rect 3052 35634 3108 35646
rect 3948 35698 4004 35710
rect 3948 35646 3950 35698
rect 4002 35646 4004 35698
rect 3948 35588 4004 35646
rect 3948 35522 4004 35532
rect 3052 35364 3108 35374
rect 3052 34914 3108 35308
rect 4508 35364 4564 35758
rect 4844 35812 4900 35822
rect 4844 35718 4900 35756
rect 4508 35298 4564 35308
rect 4844 35588 4900 35598
rect 5068 35588 5124 37100
rect 6636 36596 6692 39200
rect 9100 39060 9156 39200
rect 9436 39060 9492 39228
rect 9100 39004 9492 39060
rect 7084 37044 7140 37054
rect 6972 36596 7028 36606
rect 6636 36594 7028 36596
rect 6636 36542 6974 36594
rect 7026 36542 7028 36594
rect 6636 36540 7028 36542
rect 6972 36530 7028 36540
rect 6076 36484 6132 36494
rect 5292 36372 5348 36382
rect 5292 35922 5348 36316
rect 5292 35870 5294 35922
rect 5346 35870 5348 35922
rect 5292 35812 5348 35870
rect 5628 36258 5684 36270
rect 5628 36206 5630 36258
rect 5682 36206 5684 36258
rect 5628 35924 5684 36206
rect 5628 35858 5684 35868
rect 6076 36258 6132 36428
rect 6076 36206 6078 36258
rect 6130 36206 6132 36258
rect 5292 35746 5348 35756
rect 4900 35532 5124 35588
rect 3052 34862 3054 34914
rect 3106 34862 3108 34914
rect 3052 34850 3108 34862
rect 3948 35028 4004 35038
rect 3948 34914 4004 34972
rect 4396 35028 4452 35038
rect 4396 34934 4452 34972
rect 4844 35026 4900 35532
rect 4844 34974 4846 35026
rect 4898 34974 4900 35026
rect 4844 34962 4900 34974
rect 3948 34862 3950 34914
rect 4002 34862 4004 34914
rect 3948 34850 4004 34862
rect 3052 34692 3108 34702
rect 3052 34130 3108 34636
rect 3612 34692 3668 34702
rect 3612 34598 3668 34636
rect 3052 34078 3054 34130
rect 3106 34078 3108 34130
rect 3052 34066 3108 34078
rect 3724 33572 3780 33582
rect 3164 33460 3220 33470
rect 3164 33346 3220 33404
rect 3612 33460 3668 33470
rect 3612 33366 3668 33404
rect 3164 33294 3166 33346
rect 3218 33294 3220 33346
rect 3164 33282 3220 33294
rect 2828 33124 2884 33134
rect 2828 33122 2996 33124
rect 2828 33070 2830 33122
rect 2882 33070 2996 33122
rect 2828 33068 2996 33070
rect 2828 33058 2884 33068
rect 2828 32674 2884 32686
rect 2828 32622 2830 32674
rect 2882 32622 2884 32674
rect 2828 31948 2884 32622
rect 2604 31892 2884 31948
rect 2604 26292 2660 31892
rect 2940 31778 2996 33068
rect 3612 32788 3668 32798
rect 3724 32788 3780 33516
rect 3164 32786 3780 32788
rect 3164 32734 3614 32786
rect 3666 32734 3780 32786
rect 3164 32732 3780 32734
rect 3164 32674 3220 32732
rect 3612 32722 3668 32732
rect 3164 32622 3166 32674
rect 3218 32622 3220 32674
rect 3164 32610 3220 32622
rect 4172 32450 4228 32462
rect 4172 32398 4174 32450
rect 4226 32398 4228 32450
rect 4172 31948 4228 32398
rect 4396 32338 4452 32350
rect 4396 32286 4398 32338
rect 4450 32286 4452 32338
rect 4396 31948 4452 32286
rect 4732 32338 4788 32350
rect 4732 32286 4734 32338
rect 4786 32286 4788 32338
rect 4172 31892 4340 31948
rect 4396 31892 4564 31948
rect 2940 31726 2942 31778
rect 2994 31726 2996 31778
rect 2940 31714 2996 31726
rect 3052 31668 3108 31678
rect 2716 31106 2772 31118
rect 2716 31054 2718 31106
rect 2770 31054 2772 31106
rect 2716 27524 2772 31054
rect 3052 31106 3108 31612
rect 3500 31668 3556 31678
rect 4284 31668 4340 31892
rect 4508 31780 4564 31892
rect 4620 31780 4676 31790
rect 4508 31778 4676 31780
rect 4508 31726 4622 31778
rect 4674 31726 4676 31778
rect 4508 31724 4676 31726
rect 4396 31668 4452 31678
rect 4284 31666 4564 31668
rect 4284 31614 4398 31666
rect 4450 31614 4564 31666
rect 4284 31612 4564 31614
rect 3500 31574 3556 31612
rect 4396 31602 4452 31612
rect 3052 31054 3054 31106
rect 3106 31054 3108 31106
rect 3052 31042 3108 31054
rect 4172 31556 4228 31566
rect 4172 30994 4228 31500
rect 4172 30942 4174 30994
rect 4226 30942 4228 30994
rect 4172 30434 4228 30942
rect 4508 30996 4564 31612
rect 4620 30996 4676 31724
rect 4732 31444 4788 32286
rect 6076 31948 6132 36206
rect 7084 35028 7140 36988
rect 9772 36594 9828 39228
rect 11536 39200 11648 40000
rect 14000 39200 14112 40000
rect 16464 39200 16576 40000
rect 18928 39200 19040 40000
rect 21392 39200 21504 40000
rect 23856 39200 23968 40000
rect 26320 39200 26432 40000
rect 28784 39200 28896 40000
rect 31248 39200 31360 40000
rect 33712 39200 33824 40000
rect 36176 39200 36288 40000
rect 38640 39200 38752 40000
rect 41104 39200 41216 40000
rect 43568 39200 43680 40000
rect 46032 39200 46144 40000
rect 48496 39200 48608 40000
rect 50960 39200 51072 40000
rect 53424 39200 53536 40000
rect 55888 39200 56000 40000
rect 56252 39228 56868 39284
rect 9772 36542 9774 36594
rect 9826 36542 9828 36594
rect 9772 36530 9828 36542
rect 9996 37604 10052 37614
rect 8092 36482 8148 36494
rect 8092 36430 8094 36482
rect 8146 36430 8148 36482
rect 8092 36148 8148 36430
rect 9996 36372 10052 37548
rect 10872 36876 11136 36886
rect 10928 36820 10976 36876
rect 11032 36820 11080 36876
rect 10872 36810 11136 36820
rect 11564 36596 11620 39200
rect 11788 36596 11844 36606
rect 11564 36594 11844 36596
rect 11564 36542 11790 36594
rect 11842 36542 11844 36594
rect 11564 36540 11844 36542
rect 14028 36596 14084 39200
rect 15484 37268 15540 37278
rect 14364 36596 14420 36606
rect 14028 36594 14420 36596
rect 14028 36542 14366 36594
rect 14418 36542 14420 36594
rect 14028 36540 14420 36542
rect 11788 36530 11844 36540
rect 14364 36530 14420 36540
rect 10668 36484 10724 36494
rect 12572 36484 12628 36494
rect 9996 36306 10052 36316
rect 10444 36482 10724 36484
rect 10444 36430 10670 36482
rect 10722 36430 10724 36482
rect 10444 36428 10724 36430
rect 8092 36082 8148 36092
rect 8540 36258 8596 36270
rect 8540 36206 8542 36258
rect 8594 36206 8596 36258
rect 8540 36148 8596 36206
rect 8540 36082 8596 36092
rect 7084 34962 7140 34972
rect 10444 35586 10500 36428
rect 10668 36418 10724 36428
rect 12348 36482 12628 36484
rect 12348 36430 12574 36482
rect 12626 36430 12628 36482
rect 12348 36428 12628 36430
rect 11900 35812 11956 35822
rect 11004 35700 11060 35710
rect 11004 35606 11060 35644
rect 11452 35700 11508 35710
rect 11900 35700 11956 35756
rect 11452 35698 11956 35700
rect 11452 35646 11454 35698
rect 11506 35646 11902 35698
rect 11954 35646 11956 35698
rect 11452 35644 11956 35646
rect 11452 35634 11508 35644
rect 11900 35634 11956 35644
rect 12012 35810 12068 35822
rect 12012 35758 12014 35810
rect 12066 35758 12068 35810
rect 12012 35700 12068 35758
rect 12236 35700 12292 35710
rect 12068 35644 12180 35700
rect 12012 35634 12068 35644
rect 10444 35534 10446 35586
rect 10498 35534 10500 35586
rect 8988 34916 9044 34926
rect 8988 34242 9044 34860
rect 8988 34190 8990 34242
rect 9042 34190 9044 34242
rect 8988 34178 9044 34190
rect 9772 34692 9828 34702
rect 7196 34130 7252 34142
rect 7196 34078 7198 34130
rect 7250 34078 7252 34130
rect 6748 34018 6804 34030
rect 6748 33966 6750 34018
rect 6802 33966 6804 34018
rect 6748 33458 6804 33966
rect 6748 33406 6750 33458
rect 6802 33406 6804 33458
rect 6748 32788 6804 33406
rect 6748 32722 6804 32732
rect 7196 33234 7252 34078
rect 8204 34130 8260 34142
rect 8204 34078 8206 34130
rect 8258 34078 8260 34130
rect 8204 33348 8260 34078
rect 9660 34018 9716 34030
rect 9660 33966 9662 34018
rect 9714 33966 9716 34018
rect 8764 33908 8820 33918
rect 8764 33458 8820 33852
rect 8764 33406 8766 33458
rect 8818 33406 8820 33458
rect 8764 33394 8820 33406
rect 7196 33182 7198 33234
rect 7250 33182 7252 33234
rect 7196 32452 7252 33182
rect 8092 33346 8260 33348
rect 8092 33294 8206 33346
rect 8258 33294 8260 33346
rect 8092 33292 8260 33294
rect 7644 33124 7700 33134
rect 7420 32788 7476 32798
rect 7420 32694 7476 32732
rect 7644 32786 7700 33068
rect 7644 32734 7646 32786
rect 7698 32734 7700 32786
rect 7644 32722 7700 32734
rect 7308 32676 7364 32686
rect 7308 32582 7364 32620
rect 8092 32676 8148 33292
rect 8204 33282 8260 33292
rect 8988 33348 9044 33358
rect 8316 32900 8372 32910
rect 8204 32788 8260 32798
rect 8204 32694 8260 32732
rect 8316 32786 8372 32844
rect 8316 32734 8318 32786
rect 8370 32734 8372 32786
rect 7196 32386 7252 32396
rect 7644 32564 7700 32574
rect 8092 32544 8148 32620
rect 8316 32676 8372 32734
rect 8316 32610 8372 32620
rect 8988 32786 9044 33292
rect 9660 33348 9716 33966
rect 9772 33458 9828 34636
rect 10444 34580 10500 35534
rect 10872 35308 11136 35318
rect 10928 35252 10976 35308
rect 11032 35252 11080 35308
rect 10872 35242 11136 35252
rect 12124 35252 12180 35644
rect 12236 35606 12292 35644
rect 12124 35186 12180 35196
rect 12012 35140 12068 35150
rect 11676 35026 11732 35038
rect 11676 34974 11678 35026
rect 11730 34974 11732 35026
rect 11340 34916 11396 34926
rect 11340 34822 11396 34860
rect 10444 34514 10500 34524
rect 11676 34244 11732 34974
rect 12012 35026 12068 35084
rect 12012 34974 12014 35026
rect 12066 34974 12068 35026
rect 12012 34962 12068 34974
rect 11676 34178 11732 34188
rect 12348 34354 12404 36428
rect 12572 36418 12628 36428
rect 13692 36484 13748 36494
rect 12684 35698 12740 35710
rect 12684 35646 12686 35698
rect 12738 35646 12740 35698
rect 12684 34914 12740 35646
rect 12908 35700 12964 35710
rect 12908 35606 12964 35644
rect 13580 35698 13636 35710
rect 13580 35646 13582 35698
rect 13634 35646 13636 35698
rect 13244 35028 13300 35038
rect 12684 34862 12686 34914
rect 12738 34862 12740 34914
rect 12684 34850 12740 34862
rect 13020 34916 13076 34926
rect 12908 34804 12964 34814
rect 12908 34710 12964 34748
rect 12348 34302 12350 34354
rect 12402 34302 12404 34354
rect 10872 33740 11136 33750
rect 10928 33684 10976 33740
rect 11032 33684 11080 33740
rect 10872 33674 11136 33684
rect 9772 33406 9774 33458
rect 9826 33406 9828 33458
rect 9772 33394 9828 33406
rect 9660 33216 9716 33292
rect 10332 33348 10388 33358
rect 10332 33254 10388 33292
rect 11452 33348 11508 33358
rect 9436 33124 9492 33134
rect 9436 33030 9492 33068
rect 9884 33122 9940 33134
rect 9884 33070 9886 33122
rect 9938 33070 9940 33122
rect 8988 32734 8990 32786
rect 9042 32734 9044 32786
rect 4956 31892 5012 31902
rect 4956 31798 5012 31836
rect 5628 31892 5684 31902
rect 6076 31892 6468 31948
rect 5628 31778 5684 31836
rect 5628 31726 5630 31778
rect 5682 31726 5684 31778
rect 5628 31714 5684 31726
rect 6188 31668 6244 31678
rect 6188 31574 6244 31612
rect 6076 31556 6132 31566
rect 6076 31462 6132 31500
rect 6300 31554 6356 31566
rect 6300 31502 6302 31554
rect 6354 31502 6356 31554
rect 4732 31378 4788 31388
rect 6300 31444 6356 31502
rect 6300 31378 6356 31388
rect 5964 31332 6020 31342
rect 5964 31106 6020 31276
rect 5964 31054 5966 31106
rect 6018 31054 6020 31106
rect 5964 31042 6020 31054
rect 5180 30996 5236 31006
rect 4620 30994 5236 30996
rect 4620 30942 5182 30994
rect 5234 30942 5236 30994
rect 4620 30940 5236 30942
rect 4508 30902 4564 30940
rect 4172 30382 4174 30434
rect 4226 30382 4228 30434
rect 4172 30370 4228 30382
rect 4060 30212 4116 30222
rect 4060 30210 4564 30212
rect 4060 30158 4062 30210
rect 4114 30158 4564 30210
rect 4060 30156 4564 30158
rect 4060 30146 4116 30156
rect 3164 30098 3220 30110
rect 3164 30046 3166 30098
rect 3218 30046 3220 30098
rect 2828 29988 2884 29998
rect 3164 29988 3220 30046
rect 2828 29986 3108 29988
rect 2828 29934 2830 29986
rect 2882 29934 3108 29986
rect 2828 29932 3108 29934
rect 2828 29922 2884 29932
rect 2828 29426 2884 29438
rect 2828 29374 2830 29426
rect 2882 29374 2884 29426
rect 2828 28530 2884 29374
rect 2828 28478 2830 28530
rect 2882 28478 2884 28530
rect 2828 28466 2884 28478
rect 2716 27468 2996 27524
rect 2828 26292 2884 26302
rect 2604 26290 2884 26292
rect 2604 26238 2830 26290
rect 2882 26238 2884 26290
rect 2604 26236 2884 26238
rect 2828 26226 2884 26236
rect 2940 26068 2996 27468
rect 2156 20132 2324 20188
rect 2380 26012 2548 26068
rect 2828 26012 2996 26068
rect 2380 20188 2436 26012
rect 2828 23938 2884 26012
rect 2828 23886 2830 23938
rect 2882 23886 2884 23938
rect 2828 23874 2884 23886
rect 2940 24722 2996 24734
rect 2940 24670 2942 24722
rect 2994 24670 2996 24722
rect 2940 23716 2996 24670
rect 2492 22596 2548 22606
rect 2492 22482 2548 22540
rect 2492 22430 2494 22482
rect 2546 22430 2548 22482
rect 2492 22418 2548 22430
rect 2828 22596 2884 22606
rect 2716 21812 2772 21822
rect 2716 21718 2772 21756
rect 2604 21700 2660 21710
rect 2380 20132 2548 20188
rect 1820 20020 1876 20030
rect 1820 19926 1876 19964
rect 1932 19122 1988 19134
rect 1932 19070 1934 19122
rect 1986 19070 1988 19122
rect 1932 18788 1988 19070
rect 1932 18722 1988 18732
rect 1932 18564 1988 18574
rect 1932 18470 1988 18508
rect 2156 17668 2212 20132
rect 2380 20020 2436 20030
rect 2380 19926 2436 19964
rect 2380 18676 2436 18686
rect 2380 18582 2436 18620
rect 2268 17668 2324 17678
rect 2156 17666 2324 17668
rect 2156 17614 2270 17666
rect 2322 17614 2324 17666
rect 2156 17612 2324 17614
rect 2044 17442 2100 17454
rect 2044 17390 2046 17442
rect 2098 17390 2100 17442
rect 2044 16882 2100 17390
rect 2044 16830 2046 16882
rect 2098 16830 2100 16882
rect 2044 16818 2100 16830
rect 2156 17444 2212 17454
rect 1932 14418 1988 14430
rect 1932 14366 1934 14418
rect 1986 14366 1988 14418
rect 1932 13860 1988 14366
rect 1932 13794 1988 13804
rect 1820 13636 1876 13646
rect 2156 13636 2212 17388
rect 2268 16210 2324 17612
rect 2492 16996 2548 20132
rect 2604 17444 2660 21644
rect 2828 21476 2884 22540
rect 2940 21810 2996 23660
rect 3052 22708 3108 29932
rect 3164 29922 3220 29932
rect 4172 29986 4228 29998
rect 4172 29934 4174 29986
rect 4226 29934 4228 29986
rect 4172 29428 4228 29934
rect 4172 29334 4228 29372
rect 4508 29426 4564 30156
rect 4620 29540 4676 29550
rect 4620 29446 4676 29484
rect 4508 29374 4510 29426
rect 4562 29374 4564 29426
rect 3612 28868 3668 28878
rect 3612 28754 3668 28812
rect 3612 28702 3614 28754
rect 3666 28702 3668 28754
rect 3164 28532 3220 28542
rect 3164 28438 3220 28476
rect 3612 28532 3668 28702
rect 3612 28466 3668 28476
rect 3388 28420 3444 28430
rect 3164 27970 3220 27982
rect 3164 27918 3166 27970
rect 3218 27918 3220 27970
rect 3164 27860 3220 27918
rect 3164 27794 3220 27804
rect 3388 27858 3444 28364
rect 3388 27806 3390 27858
rect 3442 27806 3444 27858
rect 3388 27794 3444 27806
rect 4172 27860 4228 27870
rect 4172 27186 4228 27804
rect 4284 27858 4340 27870
rect 4284 27806 4286 27858
rect 4338 27806 4340 27858
rect 4284 27748 4340 27806
rect 4284 27682 4340 27692
rect 4172 27134 4174 27186
rect 4226 27134 4228 27186
rect 4172 27122 4228 27134
rect 4508 27188 4564 29374
rect 4620 28530 4676 28542
rect 4620 28478 4622 28530
rect 4674 28478 4676 28530
rect 4620 27748 4676 28478
rect 4732 27970 4788 30940
rect 5180 30930 5236 30940
rect 4844 29986 4900 29998
rect 4844 29934 4846 29986
rect 4898 29934 4900 29986
rect 4844 29428 4900 29934
rect 4844 29316 4900 29372
rect 5404 29876 5460 29886
rect 5068 29316 5124 29326
rect 4844 29314 5124 29316
rect 4844 29262 5070 29314
rect 5122 29262 5124 29314
rect 4844 29260 5124 29262
rect 4956 28754 5012 28766
rect 4956 28702 4958 28754
rect 5010 28702 5012 28754
rect 4844 28420 4900 28430
rect 4844 28326 4900 28364
rect 4956 28196 5012 28702
rect 5068 28756 5124 29260
rect 5068 28690 5124 28700
rect 4956 28140 5348 28196
rect 5292 28082 5348 28140
rect 5292 28030 5294 28082
rect 5346 28030 5348 28082
rect 5292 28018 5348 28030
rect 5404 28082 5460 29820
rect 6412 29652 6468 31892
rect 6748 31164 7140 31220
rect 6636 30994 6692 31006
rect 6636 30942 6638 30994
rect 6690 30942 6692 30994
rect 6636 30100 6692 30942
rect 6636 30034 6692 30044
rect 6748 30210 6804 31164
rect 7084 31106 7140 31164
rect 7084 31054 7086 31106
rect 7138 31054 7140 31106
rect 7084 31042 7140 31054
rect 6860 30994 6916 31006
rect 6860 30942 6862 30994
rect 6914 30942 6916 30994
rect 6860 30660 6916 30942
rect 6972 30996 7028 31006
rect 6972 30902 7028 30940
rect 6860 30604 7252 30660
rect 6748 30158 6750 30210
rect 6802 30158 6804 30210
rect 6748 29876 6804 30158
rect 6972 30212 7028 30222
rect 7196 30212 7252 30604
rect 6972 30210 7252 30212
rect 6972 30158 6974 30210
rect 7026 30158 7252 30210
rect 6972 30156 7252 30158
rect 7644 30210 7700 32508
rect 8540 32452 8596 32462
rect 8204 31108 8260 31118
rect 8204 31014 8260 31052
rect 7644 30158 7646 30210
rect 7698 30158 7700 30210
rect 6412 29586 6468 29596
rect 6524 29820 6804 29876
rect 6860 30100 6916 30110
rect 6524 29538 6580 29820
rect 6860 29652 6916 30044
rect 6524 29486 6526 29538
rect 6578 29486 6580 29538
rect 6524 29474 6580 29486
rect 6748 29596 6916 29652
rect 6748 28866 6804 29596
rect 6972 29540 7028 30156
rect 7644 30146 7700 30158
rect 6972 29474 7028 29484
rect 7196 29428 7252 29438
rect 7196 29426 7364 29428
rect 7196 29374 7198 29426
rect 7250 29374 7364 29426
rect 7196 29372 7364 29374
rect 7196 29362 7252 29372
rect 6748 28814 6750 28866
rect 6802 28814 6804 28866
rect 6748 28802 6804 28814
rect 6860 29314 6916 29326
rect 6860 29262 6862 29314
rect 6914 29262 6916 29314
rect 6860 28644 6916 29262
rect 7084 28644 7140 28654
rect 6860 28642 7140 28644
rect 6860 28590 7086 28642
rect 7138 28590 7140 28642
rect 6860 28588 7140 28590
rect 5628 28420 5684 28430
rect 6524 28420 6580 28430
rect 5628 28418 5796 28420
rect 5628 28366 5630 28418
rect 5682 28366 5796 28418
rect 5628 28364 5796 28366
rect 5628 28354 5684 28364
rect 5404 28030 5406 28082
rect 5458 28030 5460 28082
rect 5404 28018 5460 28030
rect 5628 28084 5684 28094
rect 4732 27918 4734 27970
rect 4786 27918 4788 27970
rect 4732 27906 4788 27918
rect 5516 27860 5572 27870
rect 5516 27766 5572 27804
rect 4620 27682 4676 27692
rect 4956 27748 5012 27758
rect 4508 27122 4564 27132
rect 4956 27186 5012 27692
rect 4956 27134 4958 27186
rect 5010 27134 5012 27186
rect 4956 27122 5012 27134
rect 3724 27076 3780 27086
rect 3724 26982 3780 27020
rect 4060 27074 4116 27086
rect 4060 27022 4062 27074
rect 4114 27022 4116 27074
rect 3164 26292 3220 26302
rect 4060 26292 4116 27022
rect 3164 25506 3220 26236
rect 3724 26290 4116 26292
rect 3724 26238 4062 26290
rect 4114 26238 4116 26290
rect 3724 26236 4116 26238
rect 3612 26178 3668 26190
rect 3612 26126 3614 26178
rect 3666 26126 3668 26178
rect 3612 25956 3668 26126
rect 3612 25890 3668 25900
rect 3276 25620 3332 25630
rect 3276 25526 3332 25564
rect 3612 25620 3668 25630
rect 3164 25454 3166 25506
rect 3218 25454 3220 25506
rect 3164 25442 3220 25454
rect 3612 24834 3668 25564
rect 3724 25506 3780 26236
rect 4060 26226 4116 26236
rect 4396 27076 4452 27086
rect 3724 25454 3726 25506
rect 3778 25454 3780 25506
rect 3724 25442 3780 25454
rect 3836 26066 3892 26078
rect 3836 26014 3838 26066
rect 3890 26014 3892 26066
rect 3836 25396 3892 26014
rect 4396 25618 4452 27020
rect 5404 26516 5460 26526
rect 5628 26516 5684 28028
rect 5740 27748 5796 28364
rect 6524 28082 6580 28364
rect 6524 28030 6526 28082
rect 6578 28030 6580 28082
rect 5964 27860 6020 27870
rect 6300 27860 6356 27870
rect 5964 27858 6356 27860
rect 5964 27806 5966 27858
rect 6018 27806 6302 27858
rect 6354 27806 6356 27858
rect 5964 27804 6356 27806
rect 5964 27794 6020 27804
rect 6300 27794 6356 27804
rect 5740 27682 5796 27692
rect 5852 27188 5908 27198
rect 5852 27094 5908 27132
rect 5740 27076 5796 27086
rect 5740 26982 5796 27020
rect 6076 27076 6132 27086
rect 6076 26982 6132 27020
rect 6524 26740 6580 28030
rect 6636 27858 6692 27870
rect 6636 27806 6638 27858
rect 6690 27806 6692 27858
rect 6636 27748 6692 27806
rect 6636 27682 6692 27692
rect 5404 26514 5684 26516
rect 5404 26462 5406 26514
rect 5458 26462 5684 26514
rect 5404 26460 5684 26462
rect 6188 26684 6580 26740
rect 6188 26514 6244 26684
rect 6188 26462 6190 26514
rect 6242 26462 6244 26514
rect 5404 26450 5460 26460
rect 6188 26450 6244 26462
rect 6300 26572 6692 26628
rect 6300 26514 6356 26572
rect 6300 26462 6302 26514
rect 6354 26462 6356 26514
rect 6300 26450 6356 26462
rect 6524 26402 6580 26414
rect 6524 26350 6526 26402
rect 6578 26350 6580 26402
rect 4508 26292 4564 26302
rect 4844 26292 4900 26302
rect 4508 26290 4900 26292
rect 4508 26238 4510 26290
rect 4562 26238 4846 26290
rect 4898 26238 4900 26290
rect 4508 26236 4900 26238
rect 4508 26226 4564 26236
rect 4844 26226 4900 26236
rect 5292 26292 5348 26302
rect 5292 26198 5348 26236
rect 5516 26290 5572 26302
rect 5516 26238 5518 26290
rect 5570 26238 5572 26290
rect 4396 25566 4398 25618
rect 4450 25566 4452 25618
rect 4396 25554 4452 25566
rect 4620 25956 4676 25966
rect 4620 25506 4676 25900
rect 5516 25620 5572 26238
rect 6076 26290 6132 26302
rect 6076 26238 6078 26290
rect 6130 26238 6132 26290
rect 6076 25620 6132 26238
rect 6188 25620 6244 25630
rect 6076 25618 6468 25620
rect 6076 25566 6190 25618
rect 6242 25566 6468 25618
rect 6076 25564 6468 25566
rect 5516 25554 5572 25564
rect 6188 25554 6244 25564
rect 4620 25454 4622 25506
rect 4674 25454 4676 25506
rect 4620 25442 4676 25454
rect 4284 25396 4340 25406
rect 3836 25394 4340 25396
rect 3836 25342 4286 25394
rect 4338 25342 4340 25394
rect 3836 25340 4340 25342
rect 3612 24782 3614 24834
rect 3666 24782 3668 24834
rect 3612 24770 3668 24782
rect 4060 24722 4116 25340
rect 4284 25330 4340 25340
rect 5292 25172 5348 25182
rect 4284 25116 4900 25172
rect 4284 24946 4340 25116
rect 4284 24894 4286 24946
rect 4338 24894 4340 24946
rect 4284 24882 4340 24894
rect 4396 24948 4452 24958
rect 4060 24670 4062 24722
rect 4114 24670 4116 24722
rect 3164 24610 3220 24622
rect 3164 24558 3166 24610
rect 3218 24558 3220 24610
rect 3164 23828 3220 24558
rect 4060 24500 4116 24670
rect 3724 24444 4116 24500
rect 4396 24834 4452 24892
rect 4396 24782 4398 24834
rect 4450 24782 4452 24834
rect 3164 22930 3220 23772
rect 3612 23828 3668 23838
rect 3612 23734 3668 23772
rect 3500 23156 3556 23166
rect 3724 23156 3780 24444
rect 3948 24052 4004 24062
rect 3948 24050 4340 24052
rect 3948 23998 3950 24050
rect 4002 23998 4340 24050
rect 3948 23996 4340 23998
rect 3948 23986 4004 23996
rect 3836 23716 3892 23726
rect 3836 23622 3892 23660
rect 4284 23266 4340 23996
rect 4396 24050 4452 24782
rect 4396 23998 4398 24050
rect 4450 23998 4452 24050
rect 4396 23492 4452 23998
rect 4844 24610 4900 25116
rect 4844 24558 4846 24610
rect 4898 24558 4900 24610
rect 4396 23426 4452 23436
rect 4732 23492 4788 23502
rect 4508 23268 4564 23278
rect 4284 23214 4286 23266
rect 4338 23214 4340 23266
rect 4284 23202 4340 23214
rect 4396 23266 4564 23268
rect 4396 23214 4510 23266
rect 4562 23214 4564 23266
rect 4396 23212 4564 23214
rect 3500 23154 3780 23156
rect 3500 23102 3502 23154
rect 3554 23102 3780 23154
rect 3500 23100 3780 23102
rect 3500 23090 3556 23100
rect 3164 22878 3166 22930
rect 3218 22878 3220 22930
rect 3164 22866 3220 22878
rect 3388 23044 3444 23054
rect 3052 22652 3220 22708
rect 3052 22484 3108 22494
rect 3052 22390 3108 22428
rect 2940 21758 2942 21810
rect 2994 21758 2996 21810
rect 2940 21746 2996 21758
rect 2716 21420 2884 21476
rect 2716 19906 2772 21420
rect 3164 21364 3220 22652
rect 3388 22596 3444 22988
rect 3500 22596 3556 22606
rect 3388 22594 3556 22596
rect 3388 22542 3502 22594
rect 3554 22542 3556 22594
rect 3388 22540 3556 22542
rect 3388 22484 3444 22540
rect 3388 22418 3444 22428
rect 3052 21308 3220 21364
rect 3052 20916 3108 21308
rect 3052 20802 3108 20860
rect 3052 20750 3054 20802
rect 3106 20750 3108 20802
rect 3052 20738 3108 20750
rect 3164 21028 3220 21038
rect 2716 19854 2718 19906
rect 2770 19854 2772 19906
rect 2716 18676 2772 19854
rect 3052 19234 3108 19246
rect 3052 19182 3054 19234
rect 3106 19182 3108 19234
rect 3052 19124 3108 19182
rect 3052 19058 3108 19068
rect 2716 18610 2772 18620
rect 2604 17378 2660 17388
rect 2828 18562 2884 18574
rect 2828 18510 2830 18562
rect 2882 18510 2884 18562
rect 2268 16158 2270 16210
rect 2322 16158 2324 16210
rect 2268 16146 2324 16158
rect 2380 16940 2548 16996
rect 2380 15538 2436 16940
rect 2492 16770 2548 16782
rect 2492 16718 2494 16770
rect 2546 16718 2548 16770
rect 2492 16324 2548 16718
rect 2492 16258 2548 16268
rect 2828 15652 2884 18510
rect 3164 18564 3220 20972
rect 3500 20356 3556 22540
rect 3724 22258 3780 23100
rect 4396 22708 4452 23212
rect 4508 23202 4564 23212
rect 4620 22932 4676 22942
rect 4620 22838 4676 22876
rect 3836 22652 4452 22708
rect 3836 22594 3892 22652
rect 3836 22542 3838 22594
rect 3890 22542 3892 22594
rect 3836 22530 3892 22542
rect 4508 22596 4564 22606
rect 3724 22206 3726 22258
rect 3778 22206 3780 22258
rect 3724 22194 3780 22206
rect 4508 22258 4564 22540
rect 4620 22372 4676 22382
rect 4732 22372 4788 23436
rect 4620 22370 4788 22372
rect 4620 22318 4622 22370
rect 4674 22318 4788 22370
rect 4620 22316 4788 22318
rect 4620 22306 4676 22316
rect 4508 22206 4510 22258
rect 4562 22206 4564 22258
rect 4508 22194 4564 22206
rect 4284 22148 4340 22158
rect 4060 22146 4340 22148
rect 4060 22094 4286 22146
rect 4338 22094 4340 22146
rect 4060 22092 4340 22094
rect 3948 21700 4004 21710
rect 3948 21026 4004 21644
rect 3948 20974 3950 21026
rect 4002 20974 4004 21026
rect 3948 20962 4004 20974
rect 4060 21698 4116 22092
rect 4284 22082 4340 22092
rect 4060 21646 4062 21698
rect 4114 21646 4116 21698
rect 4060 20916 4116 21646
rect 4732 21700 4788 21710
rect 4284 21588 4340 21598
rect 4284 21586 4676 21588
rect 4284 21534 4286 21586
rect 4338 21534 4676 21586
rect 4284 21532 4676 21534
rect 4172 20916 4228 20926
rect 4060 20914 4228 20916
rect 4060 20862 4174 20914
rect 4226 20862 4228 20914
rect 4060 20860 4228 20862
rect 4172 20850 4228 20860
rect 3612 20580 3668 20590
rect 3612 20578 3892 20580
rect 3612 20526 3614 20578
rect 3666 20526 3892 20578
rect 3612 20524 3892 20526
rect 3612 20514 3668 20524
rect 3500 20300 3780 20356
rect 3500 20132 3556 20142
rect 3164 18432 3220 18508
rect 3388 20020 3444 20030
rect 3052 16884 3108 16894
rect 3052 16322 3108 16828
rect 3052 16270 3054 16322
rect 3106 16270 3108 16322
rect 3052 16258 3108 16270
rect 3164 16210 3220 16222
rect 3164 16158 3166 16210
rect 3218 16158 3220 16210
rect 2828 15596 2996 15652
rect 2380 15486 2382 15538
rect 2434 15486 2436 15538
rect 2380 15316 2436 15486
rect 2380 15250 2436 15260
rect 2828 15426 2884 15438
rect 2828 15374 2830 15426
rect 2882 15374 2884 15426
rect 2716 14644 2772 14654
rect 2380 13858 2436 13870
rect 2380 13806 2382 13858
rect 2434 13806 2436 13858
rect 2268 13746 2324 13758
rect 2268 13694 2270 13746
rect 2322 13694 2324 13746
rect 2268 13636 2324 13694
rect 1820 13634 2324 13636
rect 1820 13582 1822 13634
rect 1874 13582 2324 13634
rect 1820 13580 2324 13582
rect 1820 10500 1876 13580
rect 2380 13300 2436 13806
rect 2604 13748 2660 13758
rect 2604 13654 2660 13692
rect 2380 13234 2436 13244
rect 2604 13412 2660 13422
rect 2044 12740 2100 12750
rect 2492 12740 2548 12750
rect 2604 12740 2660 13356
rect 2044 12738 2212 12740
rect 2044 12686 2046 12738
rect 2098 12686 2212 12738
rect 2044 12684 2212 12686
rect 2044 12674 2100 12684
rect 1932 12066 1988 12078
rect 1932 12014 1934 12066
rect 1986 12014 1988 12066
rect 1932 11396 1988 12014
rect 2044 11732 2100 11742
rect 2044 11506 2100 11676
rect 2044 11454 2046 11506
rect 2098 11454 2100 11506
rect 2044 11442 2100 11454
rect 1932 11330 1988 11340
rect 2156 10612 2212 12684
rect 2492 12738 2660 12740
rect 2492 12686 2494 12738
rect 2546 12686 2660 12738
rect 2492 12684 2660 12686
rect 2492 12674 2548 12684
rect 2604 10724 2660 12684
rect 2604 10630 2660 10668
rect 2492 10612 2548 10622
rect 2156 10610 2548 10612
rect 2156 10558 2494 10610
rect 2546 10558 2548 10610
rect 2156 10556 2548 10558
rect 1932 10500 1988 10510
rect 1820 10498 1988 10500
rect 1820 10446 1934 10498
rect 1986 10446 1988 10498
rect 1820 10444 1988 10446
rect 1932 10388 1988 10444
rect 1932 10322 1988 10332
rect 2492 9828 2548 10556
rect 2716 10500 2772 14588
rect 2828 14530 2884 15374
rect 2828 14478 2830 14530
rect 2882 14478 2884 14530
rect 2828 14466 2884 14478
rect 2828 13300 2884 13310
rect 2828 13074 2884 13244
rect 2828 13022 2830 13074
rect 2882 13022 2884 13074
rect 2828 13010 2884 13022
rect 2940 12178 2996 15596
rect 3052 15316 3108 15326
rect 3052 15222 3108 15260
rect 3164 13972 3220 16158
rect 3388 14308 3444 19964
rect 3500 20018 3556 20076
rect 3500 19966 3502 20018
rect 3554 19966 3556 20018
rect 3500 16100 3556 19966
rect 3724 20020 3780 20300
rect 3612 19908 3668 19918
rect 3612 19814 3668 19852
rect 3612 19124 3668 19134
rect 3612 19030 3668 19068
rect 3612 17666 3668 17678
rect 3612 17614 3614 17666
rect 3666 17614 3668 17666
rect 3612 16884 3668 17614
rect 3612 16790 3668 16828
rect 3612 16100 3668 16110
rect 3500 16098 3668 16100
rect 3500 16046 3614 16098
rect 3666 16046 3668 16098
rect 3500 16044 3668 16046
rect 3612 15092 3668 16044
rect 3612 15026 3668 15036
rect 3724 14754 3780 19964
rect 3836 20018 3892 20524
rect 3836 19966 3838 20018
rect 3890 19966 3892 20018
rect 3836 19954 3892 19966
rect 4172 20020 4228 20030
rect 4284 20020 4340 21532
rect 4620 20802 4676 21532
rect 4620 20750 4622 20802
rect 4674 20750 4676 20802
rect 4620 20738 4676 20750
rect 4620 20132 4676 20142
rect 4620 20038 4676 20076
rect 4172 20018 4340 20020
rect 4172 19966 4174 20018
rect 4226 19966 4340 20018
rect 4172 19964 4340 19966
rect 4172 19954 4228 19964
rect 4396 19794 4452 19806
rect 4396 19742 4398 19794
rect 4450 19742 4452 19794
rect 3948 19348 4004 19358
rect 3948 19234 4004 19292
rect 3948 19182 3950 19234
rect 4002 19182 4004 19234
rect 3948 19170 4004 19182
rect 3836 18676 3892 18686
rect 3836 18582 3892 18620
rect 3948 18452 4004 18462
rect 4396 18452 4452 19742
rect 3948 18450 4452 18452
rect 3948 18398 3950 18450
rect 4002 18398 4452 18450
rect 3948 18396 4452 18398
rect 4620 19348 4676 19358
rect 3948 18386 4004 18396
rect 3836 18226 3892 18238
rect 3836 18174 3838 18226
rect 3890 18174 3892 18226
rect 3836 17778 3892 18174
rect 3948 17892 4004 17902
rect 3948 17798 4004 17836
rect 3836 17726 3838 17778
rect 3890 17726 3892 17778
rect 3836 16996 3892 17726
rect 4060 17444 4116 18396
rect 4620 17778 4676 19292
rect 4620 17726 4622 17778
rect 4674 17726 4676 17778
rect 4620 17714 4676 17726
rect 4060 17378 4116 17388
rect 4732 17220 4788 21644
rect 4844 20578 4900 24558
rect 5068 23044 5124 23054
rect 5068 22950 5124 22988
rect 5292 21812 5348 25116
rect 6412 24834 6468 25564
rect 6412 24782 6414 24834
rect 6466 24782 6468 24834
rect 6412 24770 6468 24782
rect 5628 23492 5684 23502
rect 5628 22482 5684 23436
rect 5628 22430 5630 22482
rect 5682 22430 5684 22482
rect 5292 21746 5348 21756
rect 5516 21812 5572 21822
rect 5516 21718 5572 21756
rect 5404 21700 5460 21710
rect 5404 21606 5460 21644
rect 5628 21588 5684 22430
rect 5516 21532 5684 21588
rect 5852 23380 5908 23390
rect 4844 20526 4846 20578
rect 4898 20526 4900 20578
rect 4844 20468 4900 20526
rect 4844 20402 4900 20412
rect 4956 20692 5012 20702
rect 4844 19908 4900 19918
rect 4844 19346 4900 19852
rect 4956 19794 5012 20636
rect 5068 20020 5124 20030
rect 5068 19926 5124 19964
rect 4956 19742 4958 19794
rect 5010 19742 5012 19794
rect 4956 19730 5012 19742
rect 4956 19460 5012 19470
rect 4956 19366 5012 19404
rect 4844 19294 4846 19346
rect 4898 19294 4900 19346
rect 4844 19236 4900 19294
rect 4844 19170 4900 19180
rect 5404 18452 5460 18462
rect 5404 18358 5460 18396
rect 4956 18338 5012 18350
rect 4956 18286 4958 18338
rect 5010 18286 5012 18338
rect 4956 17892 5012 18286
rect 4956 17826 5012 17836
rect 4956 17444 5012 17454
rect 4956 17350 5012 17388
rect 4620 17164 4788 17220
rect 3948 16996 4004 17006
rect 3836 16994 4004 16996
rect 3836 16942 3950 16994
rect 4002 16942 4004 16994
rect 3836 16940 4004 16942
rect 3948 16930 4004 16940
rect 4396 16884 4452 16894
rect 3836 16772 3892 16782
rect 3836 16678 3892 16716
rect 4060 16212 4116 16222
rect 3948 15316 4004 15326
rect 3948 15222 4004 15260
rect 3724 14702 3726 14754
rect 3778 14702 3780 14754
rect 3724 14690 3780 14702
rect 3388 14242 3444 14252
rect 3612 14532 3668 14542
rect 3164 13906 3220 13916
rect 3612 13860 3668 14476
rect 3836 14418 3892 14430
rect 3836 14366 3838 14418
rect 3890 14366 3892 14418
rect 3724 14308 3780 14318
rect 3724 14214 3780 14252
rect 3836 14196 3892 14366
rect 3836 14130 3892 14140
rect 3948 14420 4004 14430
rect 3836 13972 3892 13982
rect 3612 13804 3780 13860
rect 3388 13748 3444 13758
rect 3388 13186 3444 13692
rect 3388 13134 3390 13186
rect 3442 13134 3444 13186
rect 3388 13122 3444 13134
rect 3500 13636 3556 13646
rect 2940 12126 2942 12178
rect 2994 12126 2996 12178
rect 2940 12114 2996 12126
rect 3164 11732 3220 11742
rect 2828 11508 2884 11518
rect 2828 10834 2884 11452
rect 2828 10782 2830 10834
rect 2882 10782 2884 10834
rect 2828 10770 2884 10782
rect 3164 11394 3220 11676
rect 3276 11508 3332 11518
rect 3276 11414 3332 11452
rect 3164 11342 3166 11394
rect 3218 11342 3220 11394
rect 2492 9762 2548 9772
rect 2604 10444 2772 10500
rect 2380 9714 2436 9726
rect 2380 9662 2382 9714
rect 2434 9662 2436 9714
rect 1932 9604 1988 9614
rect 1932 9510 1988 9548
rect 2380 9604 2436 9662
rect 2604 9604 2660 10444
rect 3164 10388 3220 11342
rect 3276 10612 3332 10622
rect 3500 10612 3556 13580
rect 3612 13634 3668 13646
rect 3612 13582 3614 13634
rect 3666 13582 3668 13634
rect 3612 13074 3668 13582
rect 3612 13022 3614 13074
rect 3666 13022 3668 13074
rect 3612 11394 3668 13022
rect 3612 11342 3614 11394
rect 3666 11342 3668 11394
rect 3612 11330 3668 11342
rect 3276 10610 3668 10612
rect 3276 10558 3278 10610
rect 3330 10558 3668 10610
rect 3276 10556 3668 10558
rect 3276 10546 3332 10556
rect 3500 10388 3556 10398
rect 3164 10332 3444 10388
rect 2380 9548 2660 9604
rect 2716 9604 2772 9614
rect 2716 9602 2884 9604
rect 2716 9550 2718 9602
rect 2770 9550 2884 9602
rect 2716 9548 2884 9550
rect 1932 8932 1988 8942
rect 1932 8838 1988 8876
rect 2156 8372 2212 8382
rect 2156 8278 2212 8316
rect 1820 7924 1876 7934
rect 1820 7698 1876 7868
rect 1820 7646 1822 7698
rect 1874 7646 1876 7698
rect 1820 7634 1876 7646
rect 2268 7700 2324 7710
rect 2380 7700 2436 9548
rect 2716 9538 2772 9548
rect 2828 9042 2884 9548
rect 2828 8990 2830 9042
rect 2882 8990 2884 9042
rect 2828 8978 2884 8990
rect 3276 9602 3332 9614
rect 3276 9550 3278 9602
rect 3330 9550 3332 9602
rect 3052 8260 3108 8270
rect 3276 8260 3332 9550
rect 3052 8258 3332 8260
rect 3052 8206 3054 8258
rect 3106 8206 3332 8258
rect 3052 8204 3332 8206
rect 3052 8194 3108 8204
rect 2492 8034 2548 8046
rect 2492 7982 2494 8034
rect 2546 7982 2548 8034
rect 2492 7924 2548 7982
rect 3164 8036 3220 8046
rect 3164 7942 3220 7980
rect 2492 7858 2548 7868
rect 3276 7924 3332 8204
rect 3388 8258 3444 10332
rect 3500 10294 3556 10332
rect 3612 8932 3668 10556
rect 3724 9940 3780 13804
rect 3836 12962 3892 13916
rect 3948 13074 4004 14364
rect 4060 13858 4116 16156
rect 4396 16210 4452 16828
rect 4508 16772 4564 16782
rect 4508 16678 4564 16716
rect 4396 16158 4398 16210
rect 4450 16158 4452 16210
rect 4284 14308 4340 14318
rect 4060 13806 4062 13858
rect 4114 13806 4116 13858
rect 4060 13794 4116 13806
rect 4172 14306 4340 14308
rect 4172 14254 4286 14306
rect 4338 14254 4340 14306
rect 4172 14252 4340 14254
rect 3948 13022 3950 13074
rect 4002 13022 4004 13074
rect 3948 13010 4004 13022
rect 3836 12910 3838 12962
rect 3890 12910 3892 12962
rect 3836 12898 3892 12910
rect 4060 12964 4116 12974
rect 4172 12964 4228 14252
rect 4284 14242 4340 14252
rect 4060 12962 4228 12964
rect 4060 12910 4062 12962
rect 4114 12910 4228 12962
rect 4060 12908 4228 12910
rect 4060 12898 4116 12908
rect 4172 12852 4228 12908
rect 4172 12290 4228 12796
rect 4172 12238 4174 12290
rect 4226 12238 4228 12290
rect 4172 12226 4228 12238
rect 4396 11732 4452 16158
rect 4620 15986 4676 17164
rect 4732 16994 4788 17006
rect 4732 16942 4734 16994
rect 4786 16942 4788 16994
rect 4732 16322 4788 16942
rect 5292 16884 5348 16894
rect 5292 16790 5348 16828
rect 4844 16772 4900 16782
rect 4844 16678 4900 16716
rect 4732 16270 4734 16322
rect 4786 16270 4788 16322
rect 4732 16258 4788 16270
rect 4620 15934 4622 15986
rect 4674 15934 4676 15986
rect 4620 15922 4676 15934
rect 5516 15652 5572 21532
rect 5628 20578 5684 20590
rect 5628 20526 5630 20578
rect 5682 20526 5684 20578
rect 5628 20468 5684 20526
rect 5628 20402 5684 20412
rect 5852 20130 5908 23324
rect 6412 23044 6468 23054
rect 6412 22950 6468 22988
rect 6188 22484 6244 22494
rect 6188 22390 6244 22428
rect 6524 22370 6580 26350
rect 6636 25506 6692 26572
rect 6636 25454 6638 25506
rect 6690 25454 6692 25506
rect 6636 22930 6692 25454
rect 6860 26180 6916 26190
rect 6860 23940 6916 26124
rect 6972 25620 7028 28588
rect 7084 28578 7140 28588
rect 7308 28644 7364 29372
rect 7980 29314 8036 29326
rect 7980 29262 7982 29314
rect 8034 29262 8036 29314
rect 7308 28550 7364 28588
rect 7756 28644 7812 28654
rect 7756 28550 7812 28588
rect 7980 28644 8036 29262
rect 7980 28578 8036 28588
rect 8316 27858 8372 27870
rect 8316 27806 8318 27858
rect 8370 27806 8372 27858
rect 7084 27748 7140 27758
rect 7868 27748 7924 27758
rect 7084 27654 7140 27692
rect 7644 27746 7924 27748
rect 7644 27694 7870 27746
rect 7922 27694 7924 27746
rect 7644 27692 7924 27694
rect 7084 26852 7140 26862
rect 7084 26180 7140 26796
rect 7644 26514 7700 27692
rect 7868 27682 7924 27692
rect 8316 26964 8372 27806
rect 8540 27748 8596 32396
rect 8988 32452 9044 32734
rect 9884 32788 9940 33070
rect 9884 32722 9940 32732
rect 8988 32386 9044 32396
rect 10108 32676 10164 32686
rect 9212 31890 9268 31902
rect 9212 31838 9214 31890
rect 9266 31838 9268 31890
rect 8764 31780 8820 31790
rect 9212 31780 9268 31838
rect 8652 31108 8708 31118
rect 8652 30770 8708 31052
rect 8652 30718 8654 30770
rect 8706 30718 8708 30770
rect 8652 30436 8708 30718
rect 8652 30370 8708 30380
rect 8764 27970 8820 31724
rect 8876 31724 9268 31780
rect 9324 31780 9380 31790
rect 8876 31218 8932 31724
rect 9324 31686 9380 31724
rect 8876 31166 8878 31218
rect 8930 31166 8932 31218
rect 8876 30100 8932 31166
rect 9772 30994 9828 31006
rect 9772 30942 9774 30994
rect 9826 30942 9828 30994
rect 8988 30884 9044 30894
rect 8988 30790 9044 30828
rect 9436 30436 9492 30446
rect 9436 30210 9492 30380
rect 9436 30158 9438 30210
rect 9490 30158 9492 30210
rect 9436 30146 9492 30158
rect 9772 30210 9828 30942
rect 10108 30882 10164 32620
rect 10872 32172 11136 32182
rect 10928 32116 10976 32172
rect 11032 32116 11080 32172
rect 10872 32106 11136 32116
rect 11452 31890 11508 33292
rect 12012 33348 12068 33358
rect 12012 33254 12068 33292
rect 12348 33124 12404 34302
rect 13020 34132 13076 34860
rect 12908 34130 13076 34132
rect 12908 34078 13022 34130
rect 13074 34078 13076 34130
rect 12908 34076 13076 34078
rect 12348 33058 12404 33068
rect 12684 33346 12740 33358
rect 12684 33294 12686 33346
rect 12738 33294 12740 33346
rect 12684 32900 12740 33294
rect 12908 33346 12964 34076
rect 13020 34066 13076 34076
rect 13244 34130 13300 34972
rect 13580 35028 13636 35646
rect 13580 34962 13636 34972
rect 13692 34804 13748 36428
rect 15484 36484 15540 37212
rect 15484 36352 15540 36428
rect 15596 36372 15652 36382
rect 14364 36260 14420 36270
rect 14364 35922 14420 36204
rect 14364 35870 14366 35922
rect 14418 35870 14420 35922
rect 14364 35858 14420 35870
rect 15036 35812 15092 35822
rect 15036 35718 15092 35756
rect 15596 35812 15652 36316
rect 16380 36260 16436 36270
rect 16380 36166 16436 36204
rect 15148 35588 15204 35598
rect 15148 35494 15204 35532
rect 14812 35476 14868 35486
rect 14812 35474 14980 35476
rect 14812 35422 14814 35474
rect 14866 35422 14980 35474
rect 14812 35420 14980 35422
rect 14812 35410 14868 35420
rect 13692 34738 13748 34748
rect 13916 35252 13972 35262
rect 13916 35026 13972 35196
rect 13916 34974 13918 35026
rect 13970 34974 13972 35026
rect 13916 34468 13972 34974
rect 14140 35028 14196 35038
rect 14140 34934 14196 34972
rect 14924 35028 14980 35420
rect 15036 35252 15092 35262
rect 15036 35138 15092 35196
rect 15036 35086 15038 35138
rect 15090 35086 15092 35138
rect 15036 35074 15092 35086
rect 14364 34916 14420 34926
rect 14364 34822 14420 34860
rect 14588 34916 14644 34926
rect 14588 34914 14868 34916
rect 14588 34862 14590 34914
rect 14642 34862 14868 34914
rect 14588 34860 14868 34862
rect 14588 34850 14644 34860
rect 13692 34412 13972 34468
rect 13468 34244 13524 34254
rect 13468 34150 13524 34188
rect 13244 34078 13246 34130
rect 13298 34078 13300 34130
rect 13244 34066 13300 34078
rect 13692 34130 13748 34412
rect 13692 34078 13694 34130
rect 13746 34078 13748 34130
rect 13692 33684 13748 34078
rect 13692 33618 13748 33628
rect 13804 34244 13860 34254
rect 14588 34244 14644 34254
rect 13804 34242 14644 34244
rect 13804 34190 13806 34242
rect 13858 34190 14590 34242
rect 14642 34190 14644 34242
rect 13804 34188 14644 34190
rect 13804 33570 13860 34188
rect 14588 34178 14644 34188
rect 14700 34244 14756 34254
rect 14700 34018 14756 34188
rect 14700 33966 14702 34018
rect 14754 33966 14756 34018
rect 14700 33954 14756 33966
rect 14364 33908 14420 33918
rect 14364 33814 14420 33852
rect 14812 33908 14868 34860
rect 14812 33842 14868 33852
rect 13804 33518 13806 33570
rect 13858 33518 13860 33570
rect 13804 33506 13860 33518
rect 14364 33684 14420 33694
rect 14364 33458 14420 33628
rect 14364 33406 14366 33458
rect 14418 33406 14420 33458
rect 14364 33394 14420 33406
rect 12908 33294 12910 33346
rect 12962 33294 12964 33346
rect 12908 33282 12964 33294
rect 13804 33348 13860 33358
rect 13132 33236 13188 33246
rect 13132 32900 13188 33180
rect 13692 33236 13748 33246
rect 13692 33142 13748 33180
rect 13804 33234 13860 33292
rect 13804 33182 13806 33234
rect 13858 33182 13860 33234
rect 13804 33170 13860 33182
rect 12684 32844 13188 32900
rect 13132 32786 13188 32844
rect 13132 32734 13134 32786
rect 13186 32734 13188 32786
rect 13132 32722 13188 32734
rect 11452 31838 11454 31890
rect 11506 31838 11508 31890
rect 11452 31826 11508 31838
rect 12796 32674 12852 32686
rect 12796 32622 12798 32674
rect 12850 32622 12852 32674
rect 10444 31780 10500 31790
rect 10444 30994 10500 31724
rect 10444 30942 10446 30994
rect 10498 30942 10500 30994
rect 10444 30930 10500 30942
rect 10668 31778 10724 31790
rect 10668 31726 10670 31778
rect 10722 31726 10724 31778
rect 10108 30830 10110 30882
rect 10162 30830 10164 30882
rect 10108 30818 10164 30830
rect 10332 30884 10388 30894
rect 10332 30790 10388 30828
rect 10668 30548 10724 31726
rect 11900 31554 11956 31566
rect 11900 31502 11902 31554
rect 11954 31502 11956 31554
rect 10872 30604 11136 30614
rect 10928 30548 10976 30604
rect 11032 30548 11080 30604
rect 10872 30538 11136 30548
rect 10668 30482 10724 30492
rect 9772 30158 9774 30210
rect 9826 30158 9828 30210
rect 9772 30146 9828 30158
rect 9884 30436 9940 30446
rect 8876 30034 8932 30044
rect 9548 30100 9604 30110
rect 9548 30006 9604 30044
rect 9884 29650 9940 30380
rect 11900 30436 11956 31502
rect 12796 31220 12852 32622
rect 14924 32674 14980 34972
rect 15260 34580 15316 34590
rect 15148 34018 15204 34030
rect 15148 33966 15150 34018
rect 15202 33966 15204 34018
rect 15148 33684 15204 33966
rect 15148 33618 15204 33628
rect 14924 32622 14926 32674
rect 14978 32622 14980 32674
rect 14924 32610 14980 32622
rect 15260 32676 15316 34524
rect 15596 34356 15652 35756
rect 16492 35812 16548 39200
rect 18844 37380 18900 37390
rect 17500 36484 17556 36494
rect 17276 36482 17556 36484
rect 17276 36430 17502 36482
rect 17554 36430 17556 36482
rect 17276 36428 17556 36430
rect 16716 36370 16772 36382
rect 16716 36318 16718 36370
rect 16770 36318 16772 36370
rect 16492 35746 16548 35756
rect 16604 36148 16660 36158
rect 16380 35700 16436 35710
rect 16380 35606 16436 35644
rect 16044 35588 16100 35598
rect 16044 35494 16100 35532
rect 16380 34916 16436 34926
rect 16380 34822 16436 34860
rect 15820 34804 15876 34814
rect 15820 34710 15876 34748
rect 16492 34356 16548 34366
rect 15596 34354 16548 34356
rect 15596 34302 15598 34354
rect 15650 34302 16494 34354
rect 16546 34302 16548 34354
rect 15596 34300 16548 34302
rect 15596 34290 15652 34300
rect 16492 34290 16548 34300
rect 15260 32610 15316 32620
rect 13020 32564 13076 32574
rect 13020 32470 13076 32508
rect 13244 32562 13300 32574
rect 13244 32510 13246 32562
rect 13298 32510 13300 32562
rect 13244 32452 13300 32510
rect 14028 32564 14084 32574
rect 14028 32470 14084 32508
rect 14252 32564 14308 32574
rect 13244 32386 13300 32396
rect 14140 32452 14196 32462
rect 14140 32002 14196 32396
rect 14140 31950 14142 32002
rect 14194 31950 14196 32002
rect 13804 31892 14084 31948
rect 14140 31938 14196 31950
rect 12796 31154 12852 31164
rect 13468 31220 13524 31230
rect 13468 31126 13524 31164
rect 13692 31220 13748 31230
rect 13804 31220 13860 31892
rect 13692 31218 13860 31220
rect 13692 31166 13694 31218
rect 13746 31166 13860 31218
rect 13692 31164 13860 31166
rect 13916 31778 13972 31790
rect 13916 31726 13918 31778
rect 13970 31726 13972 31778
rect 13692 31154 13748 31164
rect 11900 30370 11956 30380
rect 12460 30996 12516 31006
rect 10332 30324 10388 30334
rect 10332 30210 10388 30268
rect 10668 30324 10724 30334
rect 10332 30158 10334 30210
rect 10386 30158 10388 30210
rect 10332 30146 10388 30158
rect 10556 30212 10612 30222
rect 10444 30100 10500 30110
rect 10444 30006 10500 30044
rect 9884 29598 9886 29650
rect 9938 29598 9940 29650
rect 9884 29586 9940 29598
rect 10556 28868 10612 30156
rect 10668 29314 10724 30268
rect 11564 30324 11620 30334
rect 11564 30230 11620 30268
rect 11004 30210 11060 30222
rect 11004 30158 11006 30210
rect 11058 30158 11060 30210
rect 11004 29652 11060 30158
rect 11788 30212 11844 30222
rect 11788 30118 11844 30156
rect 12460 30210 12516 30940
rect 13804 30996 13860 31006
rect 13916 30996 13972 31726
rect 14028 31780 14084 31892
rect 14140 31780 14196 31790
rect 14028 31724 14140 31780
rect 14140 31648 14196 31724
rect 13860 30940 13972 30996
rect 13804 30864 13860 30940
rect 12460 30158 12462 30210
rect 12514 30158 12516 30210
rect 12460 30146 12516 30158
rect 13692 30436 13748 30446
rect 12908 29986 12964 29998
rect 12908 29934 12910 29986
rect 12962 29934 12964 29986
rect 12908 29876 12964 29934
rect 12908 29810 12964 29820
rect 11004 29586 11060 29596
rect 12124 29652 12180 29662
rect 12124 29558 12180 29596
rect 12348 29538 12404 29550
rect 12348 29486 12350 29538
rect 12402 29486 12404 29538
rect 11452 29428 11508 29438
rect 11452 29334 11508 29372
rect 12348 29428 12404 29486
rect 10668 29262 10670 29314
rect 10722 29262 10724 29314
rect 10668 29250 10724 29262
rect 11340 29316 11396 29326
rect 11340 29222 11396 29260
rect 12124 29316 12180 29326
rect 10872 29036 11136 29046
rect 10928 28980 10976 29036
rect 11032 28980 11080 29036
rect 10872 28970 11136 28980
rect 10668 28868 10724 28878
rect 10556 28866 10724 28868
rect 10556 28814 10670 28866
rect 10722 28814 10724 28866
rect 10556 28812 10724 28814
rect 10668 28802 10724 28812
rect 10444 28754 10500 28766
rect 10444 28702 10446 28754
rect 10498 28702 10500 28754
rect 8764 27918 8766 27970
rect 8818 27918 8820 27970
rect 8764 27906 8820 27918
rect 9884 28644 9940 28654
rect 10332 28644 10388 28654
rect 8540 27692 8932 27748
rect 8764 27300 8820 27310
rect 8316 26898 8372 26908
rect 8652 26964 8708 26974
rect 8652 26870 8708 26908
rect 8204 26852 8260 26862
rect 8204 26758 8260 26796
rect 7644 26462 7646 26514
rect 7698 26462 7700 26514
rect 7420 26404 7476 26414
rect 7084 26114 7140 26124
rect 7308 26290 7364 26302
rect 7308 26238 7310 26290
rect 7362 26238 7364 26290
rect 7308 26180 7364 26238
rect 7308 26114 7364 26124
rect 7084 25620 7140 25630
rect 6972 25618 7140 25620
rect 6972 25566 7086 25618
rect 7138 25566 7140 25618
rect 6972 25564 7140 25566
rect 7084 25554 7140 25564
rect 7420 25620 7476 26348
rect 7644 25956 7700 26462
rect 8652 26516 8708 26526
rect 8764 26516 8820 27244
rect 8876 27186 8932 27692
rect 8876 27134 8878 27186
rect 8930 27134 8932 27186
rect 8876 27122 8932 27134
rect 9212 27188 9268 27198
rect 8876 26962 8932 26974
rect 8876 26910 8878 26962
rect 8930 26910 8932 26962
rect 8876 26852 8932 26910
rect 9100 26964 9156 26974
rect 9212 26964 9268 27132
rect 9548 27188 9604 27198
rect 9548 27094 9604 27132
rect 9100 26962 9268 26964
rect 9100 26910 9102 26962
rect 9154 26910 9268 26962
rect 9100 26908 9268 26910
rect 9100 26898 9156 26908
rect 8876 26786 8932 26796
rect 8652 26514 8820 26516
rect 8652 26462 8654 26514
rect 8706 26462 8820 26514
rect 8652 26460 8820 26462
rect 9548 26740 9604 26750
rect 8652 26450 8708 26460
rect 7980 26404 8036 26414
rect 7980 26310 8036 26348
rect 8876 26404 8932 26414
rect 7644 25890 7700 25900
rect 7756 26292 7812 26302
rect 7420 25554 7476 25564
rect 7756 25618 7812 26236
rect 8876 26068 8932 26348
rect 8876 26002 8932 26012
rect 8988 26290 9044 26302
rect 8988 26238 8990 26290
rect 9042 26238 9044 26290
rect 7756 25566 7758 25618
rect 7810 25566 7812 25618
rect 7756 25554 7812 25566
rect 7980 25506 8036 25518
rect 7980 25454 7982 25506
rect 8034 25454 8036 25506
rect 7644 25396 7700 25406
rect 7196 25394 7700 25396
rect 7196 25342 7646 25394
rect 7698 25342 7700 25394
rect 7196 25340 7700 25342
rect 7084 24724 7140 24734
rect 7084 24630 7140 24668
rect 7196 24164 7252 25340
rect 7644 25330 7700 25340
rect 7980 24836 8036 25454
rect 8652 25282 8708 25294
rect 8652 25230 8654 25282
rect 8706 25230 8708 25282
rect 8092 24836 8148 24846
rect 7980 24834 8148 24836
rect 7980 24782 8094 24834
rect 8146 24782 8148 24834
rect 7980 24780 8148 24782
rect 7308 24612 7364 24622
rect 7980 24612 8036 24622
rect 7308 24610 8036 24612
rect 7308 24558 7310 24610
rect 7362 24558 7982 24610
rect 8034 24558 8036 24610
rect 7308 24556 8036 24558
rect 7308 24546 7364 24556
rect 7980 24546 8036 24556
rect 7420 24388 7476 24398
rect 7308 24164 7364 24174
rect 7196 24162 7364 24164
rect 7196 24110 7310 24162
rect 7362 24110 7364 24162
rect 7196 24108 7364 24110
rect 7308 24098 7364 24108
rect 7420 24162 7476 24332
rect 7420 24110 7422 24162
rect 7474 24110 7476 24162
rect 7420 24098 7476 24110
rect 7644 24164 7700 24174
rect 7644 24070 7700 24108
rect 8092 24164 8148 24780
rect 8316 24500 8372 24510
rect 8652 24500 8708 25230
rect 8988 25284 9044 26238
rect 9212 25284 9268 25294
rect 8988 25282 9268 25284
rect 8988 25230 9214 25282
rect 9266 25230 9268 25282
rect 8988 25228 9268 25230
rect 8316 24498 8708 24500
rect 8316 24446 8318 24498
rect 8370 24446 8708 24498
rect 8316 24444 8708 24446
rect 9100 24610 9156 24622
rect 9100 24558 9102 24610
rect 9154 24558 9156 24610
rect 8316 24434 8372 24444
rect 8092 24098 8148 24108
rect 8428 24050 8484 24444
rect 9100 24162 9156 24558
rect 9100 24110 9102 24162
rect 9154 24110 9156 24162
rect 9100 24098 9156 24110
rect 8428 23998 8430 24050
rect 8482 23998 8484 24050
rect 7868 23940 7924 23950
rect 6860 23884 7364 23940
rect 6972 23156 7028 23166
rect 6636 22878 6638 22930
rect 6690 22878 6692 22930
rect 6636 22866 6692 22878
rect 6748 23100 6972 23156
rect 6524 22318 6526 22370
rect 6578 22318 6580 22370
rect 6524 22306 6580 22318
rect 6748 22484 6804 23100
rect 6972 23062 7028 23100
rect 7084 23044 7140 23054
rect 7084 22596 7140 22988
rect 6748 22258 6804 22428
rect 6860 22540 7140 22596
rect 6860 22370 6916 22540
rect 6860 22318 6862 22370
rect 6914 22318 6916 22370
rect 6860 22306 6916 22318
rect 6748 22206 6750 22258
rect 6802 22206 6804 22258
rect 6748 22194 6804 22206
rect 6972 21700 7028 21710
rect 6972 21606 7028 21644
rect 7196 21700 7252 21710
rect 7196 21606 7252 21644
rect 6636 21588 6692 21598
rect 6636 21494 6692 21532
rect 7308 21588 7364 23884
rect 7868 23846 7924 23884
rect 8428 23940 8484 23998
rect 8428 23874 8484 23884
rect 9212 23716 9268 25228
rect 9548 24162 9604 26684
rect 9660 26178 9716 26190
rect 9660 26126 9662 26178
rect 9714 26126 9716 26178
rect 9660 26068 9716 26126
rect 9660 26002 9716 26012
rect 9772 25282 9828 25294
rect 9772 25230 9774 25282
rect 9826 25230 9828 25282
rect 9660 24724 9716 24734
rect 9660 24630 9716 24668
rect 9548 24110 9550 24162
rect 9602 24110 9604 24162
rect 9548 24098 9604 24110
rect 8764 23604 8820 23614
rect 8204 23156 8260 23166
rect 8204 23062 8260 23100
rect 7756 23044 7812 23054
rect 7644 22370 7700 22382
rect 7644 22318 7646 22370
rect 7698 22318 7700 22370
rect 7644 21812 7700 22318
rect 7644 21746 7700 21756
rect 7756 21810 7812 22988
rect 8540 22484 8596 22494
rect 8540 22390 8596 22428
rect 8092 22370 8148 22382
rect 8092 22318 8094 22370
rect 8146 22318 8148 22370
rect 8092 22260 8148 22318
rect 8092 22194 8148 22204
rect 7756 21758 7758 21810
rect 7810 21758 7812 21810
rect 7756 21746 7812 21758
rect 8204 21700 8260 21710
rect 8204 21606 8260 21644
rect 8540 21700 8596 21710
rect 6524 20916 6580 20926
rect 6524 20822 6580 20860
rect 7196 20804 7252 20814
rect 6076 20692 6132 20702
rect 6076 20598 6132 20636
rect 5852 20078 5854 20130
rect 5906 20078 5908 20130
rect 5852 20066 5908 20078
rect 5740 20018 5796 20030
rect 5740 19966 5742 20018
rect 5794 19966 5796 20018
rect 5740 19348 5796 19966
rect 5964 20018 6020 20030
rect 5964 19966 5966 20018
rect 6018 19966 6020 20018
rect 5964 19460 6020 19966
rect 6412 20020 6468 20030
rect 6412 20018 6692 20020
rect 6412 19966 6414 20018
rect 6466 19966 6692 20018
rect 6412 19964 6692 19966
rect 6412 19954 6468 19964
rect 5964 19394 6020 19404
rect 5852 19348 5908 19358
rect 5740 19346 5908 19348
rect 5740 19294 5854 19346
rect 5906 19294 5908 19346
rect 5740 19292 5908 19294
rect 5852 18562 5908 19292
rect 6076 19236 6132 19246
rect 6076 19142 6132 19180
rect 5852 18510 5854 18562
rect 5906 18510 5908 18562
rect 5852 18498 5908 18510
rect 6524 18562 6580 18574
rect 6524 18510 6526 18562
rect 6578 18510 6580 18562
rect 6412 18452 6468 18462
rect 5964 18450 6468 18452
rect 5964 18398 6414 18450
rect 6466 18398 6468 18450
rect 5964 18396 6468 18398
rect 5740 17892 5796 17902
rect 5740 17778 5796 17836
rect 5852 17892 5908 17902
rect 5964 17892 6020 18396
rect 6412 18386 6468 18396
rect 6524 18452 6580 18510
rect 6524 18386 6580 18396
rect 6524 18228 6580 18238
rect 6636 18228 6692 19964
rect 6748 19796 6804 19806
rect 6748 19346 6804 19740
rect 6748 19294 6750 19346
rect 6802 19294 6804 19346
rect 6748 19282 6804 19294
rect 6524 18226 6692 18228
rect 6524 18174 6526 18226
rect 6578 18174 6692 18226
rect 6524 18172 6692 18174
rect 6524 18162 6580 18172
rect 5852 17890 6020 17892
rect 5852 17838 5854 17890
rect 5906 17838 6020 17890
rect 5852 17836 6020 17838
rect 5852 17826 5908 17836
rect 5740 17726 5742 17778
rect 5794 17726 5796 17778
rect 5740 17714 5796 17726
rect 6972 17668 7028 17678
rect 6972 17574 7028 17612
rect 6860 17442 6916 17454
rect 7084 17444 7140 17454
rect 6860 17390 6862 17442
rect 6914 17390 6916 17442
rect 6860 16548 6916 17390
rect 6972 17442 7140 17444
rect 6972 17390 7086 17442
rect 7138 17390 7140 17442
rect 6972 17388 7140 17390
rect 6972 16882 7028 17388
rect 7084 17378 7140 17388
rect 6972 16830 6974 16882
rect 7026 16830 7028 16882
rect 6972 16772 7028 16830
rect 6972 16706 7028 16716
rect 7084 16770 7140 16782
rect 7084 16718 7086 16770
rect 7138 16718 7140 16770
rect 7084 16548 7140 16718
rect 6860 16492 7140 16548
rect 6860 16322 6916 16492
rect 6860 16270 6862 16322
rect 6914 16270 6916 16322
rect 6860 16258 6916 16270
rect 6188 16212 6244 16222
rect 6188 16118 6244 16156
rect 6636 16100 6692 16110
rect 6636 16006 6692 16044
rect 5516 15596 5908 15652
rect 4844 15316 4900 15326
rect 4508 15204 4564 15214
rect 4508 14418 4564 15148
rect 4620 14532 4676 14542
rect 4620 14438 4676 14476
rect 4508 14366 4510 14418
rect 4562 14366 4564 14418
rect 4508 14354 4564 14366
rect 4844 14084 4900 15260
rect 5404 15316 5460 15326
rect 5404 15222 5460 15260
rect 4620 14028 4900 14084
rect 4956 15202 5012 15214
rect 4956 15150 4958 15202
rect 5010 15150 5012 15202
rect 4956 15092 5012 15150
rect 4508 13972 4564 13982
rect 4508 13878 4564 13916
rect 4620 13412 4676 14028
rect 4732 13858 4788 13870
rect 4732 13806 4734 13858
rect 4786 13806 4788 13858
rect 4732 13636 4788 13806
rect 4844 13748 4900 13758
rect 4844 13654 4900 13692
rect 4732 13570 4788 13580
rect 4956 13524 5012 15036
rect 5516 14532 5572 15596
rect 5852 15538 5908 15596
rect 5852 15486 5854 15538
rect 5906 15486 5908 15538
rect 5852 15474 5908 15486
rect 7196 15148 7252 20748
rect 5628 15092 5684 15102
rect 5628 14642 5684 15036
rect 5628 14590 5630 14642
rect 5682 14590 5684 14642
rect 5628 14578 5684 14590
rect 6860 15092 7252 15148
rect 5516 14466 5572 14476
rect 6076 14308 6132 14318
rect 6132 14252 6244 14308
rect 6076 14176 6132 14252
rect 5516 13748 5572 13758
rect 5740 13748 5796 13758
rect 5572 13746 5796 13748
rect 5572 13694 5742 13746
rect 5794 13694 5796 13746
rect 5572 13692 5796 13694
rect 5292 13636 5348 13646
rect 5292 13542 5348 13580
rect 4956 13458 5012 13468
rect 4620 13346 4676 13356
rect 4844 12852 4900 12862
rect 4844 12758 4900 12796
rect 4956 12850 5012 12862
rect 4956 12798 4958 12850
rect 5010 12798 5012 12850
rect 4620 12738 4676 12750
rect 4620 12686 4622 12738
rect 4674 12686 4676 12738
rect 4396 11666 4452 11676
rect 4508 12178 4564 12190
rect 4508 12126 4510 12178
rect 4562 12126 4564 12178
rect 4172 11396 4228 11406
rect 4508 11396 4564 12126
rect 4172 11302 4228 11340
rect 4284 11394 4564 11396
rect 4284 11342 4510 11394
rect 4562 11342 4564 11394
rect 4284 11340 4564 11342
rect 4620 11396 4676 12686
rect 4956 12292 5012 12798
rect 4956 12226 5012 12236
rect 4732 11396 4788 11406
rect 4620 11394 4788 11396
rect 4620 11342 4734 11394
rect 4786 11342 4788 11394
rect 4620 11340 4788 11342
rect 4284 11060 4340 11340
rect 4508 11330 4564 11340
rect 4732 11330 4788 11340
rect 4620 11172 4676 11182
rect 4620 11078 4676 11116
rect 3836 11004 4340 11060
rect 3836 10834 3892 11004
rect 3836 10782 3838 10834
rect 3890 10782 3892 10834
rect 3836 10770 3892 10782
rect 4396 10612 4452 10622
rect 4452 10556 4564 10612
rect 4396 10518 4452 10556
rect 4508 10050 4564 10556
rect 4620 10388 4676 10398
rect 4620 10386 4788 10388
rect 4620 10334 4622 10386
rect 4674 10334 4788 10386
rect 4620 10332 4788 10334
rect 4620 10322 4676 10332
rect 4508 9998 4510 10050
rect 4562 9998 4564 10050
rect 4508 9986 4564 9998
rect 4732 10164 4788 10332
rect 3724 9938 4452 9940
rect 3724 9886 3726 9938
rect 3778 9886 4452 9938
rect 3724 9884 4452 9886
rect 3724 9874 3780 9884
rect 3724 8932 3780 8942
rect 3612 8930 3780 8932
rect 3612 8878 3726 8930
rect 3778 8878 3780 8930
rect 3612 8876 3780 8878
rect 3388 8206 3390 8258
rect 3442 8206 3444 8258
rect 3388 8194 3444 8206
rect 3276 7858 3332 7868
rect 3724 8036 3780 8876
rect 3836 8372 3892 9884
rect 4396 9828 4452 9884
rect 4620 9828 4676 9838
rect 4396 9826 4676 9828
rect 4396 9774 4622 9826
rect 4674 9774 4676 9826
rect 4396 9772 4676 9774
rect 4620 9762 4676 9772
rect 4508 9604 4564 9614
rect 4508 9156 4564 9548
rect 4732 9266 4788 10108
rect 4956 10386 5012 10398
rect 4956 10334 4958 10386
rect 5010 10334 5012 10386
rect 4956 9940 5012 10334
rect 4956 9874 5012 9884
rect 5516 9828 5572 13692
rect 5740 13682 5796 13692
rect 6076 13636 6132 13646
rect 5516 9762 5572 9772
rect 5628 13524 5684 13534
rect 5628 9826 5684 13468
rect 5852 12292 5908 12302
rect 5852 12198 5908 12236
rect 6076 12290 6132 13580
rect 6076 12238 6078 12290
rect 6130 12238 6132 12290
rect 6076 12226 6132 12238
rect 6188 11956 6244 14252
rect 6636 14306 6692 14318
rect 6636 14254 6638 14306
rect 6690 14254 6692 14306
rect 6636 13748 6692 14254
rect 6636 13682 6692 13692
rect 6636 13300 6692 13310
rect 6860 13300 6916 15092
rect 7084 14420 7140 14430
rect 7084 14326 7140 14364
rect 7196 14308 7252 14318
rect 7196 14214 7252 14252
rect 6692 13244 6916 13300
rect 6636 13234 6692 13244
rect 6188 11890 6244 11900
rect 5740 11506 5796 11518
rect 5740 11454 5742 11506
rect 5794 11454 5796 11506
rect 5740 11396 5796 11454
rect 5740 11330 5796 11340
rect 5852 11508 5908 11518
rect 5852 11282 5908 11452
rect 5852 11230 5854 11282
rect 5906 11230 5908 11282
rect 5852 11218 5908 11230
rect 6076 11282 6132 11294
rect 6076 11230 6078 11282
rect 6130 11230 6132 11282
rect 6076 10612 6132 11230
rect 6076 10480 6132 10556
rect 6412 10610 6468 10622
rect 6412 10558 6414 10610
rect 6466 10558 6468 10610
rect 5628 9774 5630 9826
rect 5682 9774 5684 9826
rect 5628 9762 5684 9774
rect 5740 10388 5796 10398
rect 5740 9380 5796 10332
rect 6412 10052 6468 10558
rect 6412 9986 6468 9996
rect 5964 9714 6020 9726
rect 5964 9662 5966 9714
rect 6018 9662 6020 9714
rect 5852 9604 5908 9614
rect 5852 9510 5908 9548
rect 5740 9324 5908 9380
rect 4732 9214 4734 9266
rect 4786 9214 4788 9266
rect 4732 9202 4788 9214
rect 4508 9090 4564 9100
rect 5740 9156 5796 9166
rect 5740 9062 5796 9100
rect 3836 8306 3892 8316
rect 4284 9044 4340 9054
rect 4284 8258 4340 8988
rect 4284 8206 4286 8258
rect 4338 8206 4340 8258
rect 4284 8194 4340 8206
rect 4620 9042 4676 9054
rect 4620 8990 4622 9042
rect 4674 8990 4676 9042
rect 4620 8260 4676 8990
rect 4956 9042 5012 9054
rect 4956 8990 4958 9042
rect 5010 8990 5012 9042
rect 4844 8930 4900 8942
rect 4844 8878 4846 8930
rect 4898 8878 4900 8930
rect 4844 8484 4900 8878
rect 4956 8820 5012 8990
rect 5516 9044 5572 9054
rect 5516 8950 5572 8988
rect 5852 9042 5908 9324
rect 5852 8990 5854 9042
rect 5906 8990 5908 9042
rect 4956 8764 5124 8820
rect 4620 8166 4676 8204
rect 4732 8428 4900 8484
rect 4956 8596 5012 8606
rect 5068 8596 5124 8764
rect 5404 8708 5460 8718
rect 5068 8540 5236 8596
rect 2268 7698 2436 7700
rect 2268 7646 2270 7698
rect 2322 7646 2436 7698
rect 2268 7644 2436 7646
rect 2268 7634 2324 7644
rect 2492 7588 2548 7598
rect 1932 6578 1988 6590
rect 1932 6526 1934 6578
rect 1986 6526 1988 6578
rect 1932 6468 1988 6526
rect 1932 6402 1988 6412
rect 2492 6130 2548 7532
rect 2716 7588 2772 7598
rect 2716 7494 2772 7532
rect 3052 7586 3108 7598
rect 3052 7534 3054 7586
rect 3106 7534 3108 7586
rect 3052 6690 3108 7534
rect 3052 6638 3054 6690
rect 3106 6638 3108 6690
rect 3052 6626 3108 6638
rect 3612 7476 3668 7486
rect 2492 6078 2494 6130
rect 2546 6078 2548 6130
rect 2492 6066 2548 6078
rect 3500 6356 3556 6366
rect 3500 5906 3556 6300
rect 3500 5854 3502 5906
rect 3554 5854 3556 5906
rect 3500 5842 3556 5854
rect 3612 5682 3668 7420
rect 3724 6468 3780 7980
rect 4732 7700 4788 8428
rect 4844 8260 4900 8270
rect 4956 8260 5012 8540
rect 4844 8258 5012 8260
rect 4844 8206 4846 8258
rect 4898 8206 5012 8258
rect 4844 8204 5012 8206
rect 4844 8194 4900 8204
rect 4732 7634 4788 7644
rect 4172 7588 4228 7598
rect 4172 7474 4228 7532
rect 4172 7422 4174 7474
rect 4226 7422 4228 7474
rect 4172 7410 4228 7422
rect 4508 7476 4564 7486
rect 5068 7476 5124 7486
rect 4508 7382 4564 7420
rect 4732 7474 5124 7476
rect 4732 7422 5070 7474
rect 5122 7422 5124 7474
rect 4732 7420 5124 7422
rect 4620 7364 4676 7374
rect 4620 7270 4676 7308
rect 4732 6690 4788 7420
rect 5068 7410 5124 7420
rect 4732 6638 4734 6690
rect 4786 6638 4788 6690
rect 4732 6626 4788 6638
rect 3724 6374 3780 6412
rect 4396 6578 4452 6590
rect 4396 6526 4398 6578
rect 4450 6526 4452 6578
rect 4396 6020 4452 6526
rect 4508 6466 4564 6478
rect 4508 6414 4510 6466
rect 4562 6414 4564 6466
rect 4508 6356 4564 6414
rect 5068 6468 5124 6478
rect 5180 6468 5236 8540
rect 5404 7476 5460 8652
rect 5852 8148 5908 8990
rect 5852 8054 5908 8092
rect 5964 7924 6020 9662
rect 6412 9604 6468 9614
rect 6412 9510 6468 9548
rect 6860 9604 6916 13244
rect 7196 12740 7252 12750
rect 7308 12740 7364 21532
rect 7644 20916 7700 20926
rect 7644 20822 7700 20860
rect 8204 20804 8260 20814
rect 8204 20710 8260 20748
rect 8316 20132 8372 20142
rect 8316 19348 8372 20076
rect 8540 19460 8596 21644
rect 8764 21588 8820 23548
rect 8988 22708 9044 22718
rect 8876 21812 8932 21822
rect 8876 21698 8932 21756
rect 8988 21810 9044 22652
rect 8988 21758 8990 21810
rect 9042 21758 9044 21810
rect 8988 21746 9044 21758
rect 8876 21646 8878 21698
rect 8930 21646 8932 21698
rect 8876 21634 8932 21646
rect 8652 20916 8708 20926
rect 8764 20916 8820 21532
rect 8652 20914 8764 20916
rect 8652 20862 8654 20914
rect 8706 20862 8764 20914
rect 8652 20860 8764 20862
rect 8652 20850 8708 20860
rect 8764 20850 8820 20860
rect 9212 20692 9268 23660
rect 9660 23716 9716 23726
rect 9772 23716 9828 25230
rect 9884 25284 9940 28588
rect 10108 28642 10388 28644
rect 10108 28590 10334 28642
rect 10386 28590 10388 28642
rect 10108 28588 10388 28590
rect 10108 27300 10164 28588
rect 10332 28578 10388 28588
rect 10108 27168 10164 27244
rect 10332 28420 10388 28430
rect 9996 27076 10052 27086
rect 9996 26628 10052 27020
rect 9996 26562 10052 26572
rect 10332 26516 10388 28364
rect 10444 27746 10500 28702
rect 12124 28642 12180 29260
rect 12124 28590 12126 28642
rect 12178 28590 12180 28642
rect 10444 27694 10446 27746
rect 10498 27694 10500 27746
rect 10444 27074 10500 27694
rect 10444 27022 10446 27074
rect 10498 27022 10500 27074
rect 10444 27010 10500 27022
rect 10556 27860 10612 27870
rect 10556 27074 10612 27804
rect 11004 27858 11060 27870
rect 11004 27806 11006 27858
rect 11058 27806 11060 27858
rect 11004 27636 11060 27806
rect 11116 27746 11172 27758
rect 11116 27694 11118 27746
rect 11170 27694 11172 27746
rect 11116 27636 11172 27694
rect 12012 27746 12068 27758
rect 12012 27694 12014 27746
rect 12066 27694 12068 27746
rect 11116 27580 11396 27636
rect 11004 27570 11060 27580
rect 10872 27468 11136 27478
rect 10928 27412 10976 27468
rect 11032 27412 11080 27468
rect 10872 27402 11136 27412
rect 10556 27022 10558 27074
rect 10610 27022 10612 27074
rect 10556 27010 10612 27022
rect 11340 27074 11396 27580
rect 11340 27022 11342 27074
rect 11394 27022 11396 27074
rect 11340 27010 11396 27022
rect 10668 26964 10724 26974
rect 10668 26870 10724 26908
rect 11676 26964 11732 26974
rect 11676 26870 11732 26908
rect 10780 26850 10836 26862
rect 10780 26798 10782 26850
rect 10834 26798 10836 26850
rect 10444 26516 10500 26526
rect 10332 26514 10500 26516
rect 10332 26462 10446 26514
rect 10498 26462 10500 26514
rect 10332 26460 10500 26462
rect 10444 26450 10500 26460
rect 9884 25218 9940 25228
rect 10332 26290 10388 26302
rect 10332 26238 10334 26290
rect 10386 26238 10388 26290
rect 10332 25618 10388 26238
rect 10332 25566 10334 25618
rect 10386 25566 10388 25618
rect 9996 25172 10052 25182
rect 9884 24834 9940 24846
rect 9884 24782 9886 24834
rect 9938 24782 9940 24834
rect 9884 24162 9940 24782
rect 9884 24110 9886 24162
rect 9938 24110 9940 24162
rect 9884 24098 9940 24110
rect 9996 24722 10052 25116
rect 10332 24948 10388 25566
rect 10556 26292 10612 26302
rect 10780 26292 10836 26798
rect 11564 26850 11620 26862
rect 11564 26798 11566 26850
rect 11618 26798 11620 26850
rect 11564 26740 11620 26798
rect 11564 26674 11620 26684
rect 12012 26740 12068 27694
rect 12012 26674 12068 26684
rect 12012 26404 12068 26414
rect 12012 26310 12068 26348
rect 10556 26290 10836 26292
rect 10556 26238 10558 26290
rect 10610 26238 10836 26290
rect 10556 26236 10836 26238
rect 11004 26292 11060 26302
rect 10556 25508 10612 26236
rect 11004 26198 11060 26236
rect 11452 26290 11508 26302
rect 11452 26238 11454 26290
rect 11506 26238 11508 26290
rect 10872 25900 11136 25910
rect 10928 25844 10976 25900
rect 11032 25844 11080 25900
rect 10872 25834 11136 25844
rect 10780 25508 10836 25518
rect 10556 25506 10948 25508
rect 10556 25454 10782 25506
rect 10834 25454 10948 25506
rect 10556 25452 10948 25454
rect 10780 25442 10836 25452
rect 10780 25060 10836 25070
rect 10444 24948 10500 24958
rect 10332 24946 10500 24948
rect 10332 24894 10446 24946
rect 10498 24894 10500 24946
rect 10332 24892 10500 24894
rect 10444 24882 10500 24892
rect 9996 24670 9998 24722
rect 10050 24670 10052 24722
rect 9660 23714 9828 23716
rect 9660 23662 9662 23714
rect 9714 23662 9828 23714
rect 9660 23660 9828 23662
rect 9996 23716 10052 24670
rect 10668 24834 10724 24846
rect 10668 24782 10670 24834
rect 10722 24782 10724 24834
rect 10108 24164 10164 24174
rect 10668 24164 10724 24782
rect 10780 24834 10836 25004
rect 10780 24782 10782 24834
rect 10834 24782 10836 24834
rect 10780 24770 10836 24782
rect 10892 24500 10948 25452
rect 11228 25396 11284 25406
rect 11452 25396 11508 26238
rect 11676 26292 11732 26302
rect 11676 26178 11732 26236
rect 11788 26292 11844 26302
rect 11788 26290 11956 26292
rect 11788 26238 11790 26290
rect 11842 26238 11956 26290
rect 11788 26236 11956 26238
rect 11788 26226 11844 26236
rect 11676 26126 11678 26178
rect 11730 26126 11732 26178
rect 11676 26114 11732 26126
rect 11228 25394 11508 25396
rect 11228 25342 11230 25394
rect 11282 25342 11508 25394
rect 11228 25340 11508 25342
rect 11228 24724 11284 25340
rect 11788 25282 11844 25294
rect 11788 25230 11790 25282
rect 11842 25230 11844 25282
rect 11452 24948 11508 24958
rect 11788 24948 11844 25230
rect 11900 25172 11956 26236
rect 12124 25508 12180 28590
rect 12348 28644 12404 29372
rect 12460 29426 12516 29438
rect 12460 29374 12462 29426
rect 12514 29374 12516 29426
rect 12460 29316 12516 29374
rect 12460 29250 12516 29260
rect 12908 29316 12964 29326
rect 12908 29222 12964 29260
rect 13356 29314 13412 29326
rect 13356 29262 13358 29314
rect 13410 29262 13412 29314
rect 12572 28644 12628 28654
rect 12348 28642 12628 28644
rect 12348 28590 12574 28642
rect 12626 28590 12628 28642
rect 12348 28588 12628 28590
rect 12572 28420 12628 28588
rect 12572 28354 12628 28364
rect 13244 28532 13300 28542
rect 13244 27858 13300 28476
rect 13356 28420 13412 29262
rect 13356 28354 13412 28364
rect 13692 28196 13748 30380
rect 14028 30212 14084 30222
rect 14252 30212 14308 32508
rect 16044 32450 16100 32462
rect 16044 32398 16046 32450
rect 16098 32398 16100 32450
rect 16044 31892 16100 32398
rect 15484 31836 16100 31892
rect 14812 31780 14868 31790
rect 14028 30210 14308 30212
rect 14028 30158 14030 30210
rect 14082 30158 14308 30210
rect 14028 30156 14308 30158
rect 14028 30146 14084 30156
rect 14140 29986 14196 29998
rect 14140 29934 14142 29986
rect 14194 29934 14196 29986
rect 13916 29876 13972 29886
rect 13916 29650 13972 29820
rect 13916 29598 13918 29650
rect 13970 29598 13972 29650
rect 13916 29586 13972 29598
rect 13804 28532 13860 28542
rect 13804 28438 13860 28476
rect 14140 28420 14196 29934
rect 14252 28866 14308 30156
rect 14364 31332 14420 31342
rect 14364 30210 14420 31276
rect 14700 31220 14756 31230
rect 14700 31126 14756 31164
rect 14812 31218 14868 31724
rect 15484 31666 15540 31836
rect 15484 31614 15486 31666
rect 15538 31614 15540 31666
rect 15484 31602 15540 31614
rect 15708 31668 15764 31678
rect 15708 31574 15764 31612
rect 15596 31554 15652 31566
rect 15596 31502 15598 31554
rect 15650 31502 15652 31554
rect 14812 31166 14814 31218
rect 14866 31166 14868 31218
rect 14812 31154 14868 31166
rect 14924 31332 14980 31342
rect 14924 31218 14980 31276
rect 14924 31166 14926 31218
rect 14978 31166 14980 31218
rect 14924 31154 14980 31166
rect 15596 31220 15652 31502
rect 15596 31154 15652 31164
rect 14924 30996 14980 31006
rect 14364 30158 14366 30210
rect 14418 30158 14420 30210
rect 14364 30146 14420 30158
rect 14812 30210 14868 30222
rect 14812 30158 14814 30210
rect 14866 30158 14868 30210
rect 14812 29876 14868 30158
rect 14812 29426 14868 29820
rect 14812 29374 14814 29426
rect 14866 29374 14868 29426
rect 14812 29362 14868 29374
rect 14252 28814 14254 28866
rect 14306 28814 14308 28866
rect 14252 28802 14308 28814
rect 14812 28756 14868 28766
rect 14924 28756 14980 30940
rect 15372 30996 15428 31006
rect 15372 30994 15876 30996
rect 15372 30942 15374 30994
rect 15426 30942 15876 30994
rect 15372 30940 15876 30942
rect 15372 30930 15428 30940
rect 14812 28754 14980 28756
rect 14812 28702 14814 28754
rect 14866 28702 14980 28754
rect 14812 28700 14980 28702
rect 15036 30210 15092 30222
rect 15036 30158 15038 30210
rect 15090 30158 15092 30210
rect 15036 29314 15092 30158
rect 15820 30210 15876 30940
rect 15820 30158 15822 30210
rect 15874 30158 15876 30210
rect 15820 30146 15876 30158
rect 16044 30994 16100 31836
rect 16044 30942 16046 30994
rect 16098 30942 16100 30994
rect 15036 29262 15038 29314
rect 15090 29262 15092 29314
rect 13916 28364 14196 28420
rect 14588 28642 14644 28654
rect 14588 28590 14590 28642
rect 14642 28590 14644 28642
rect 13692 28140 13860 28196
rect 13244 27806 13246 27858
rect 13298 27806 13300 27858
rect 12124 25442 12180 25452
rect 12348 27748 12404 27758
rect 11900 25106 11956 25116
rect 12124 25282 12180 25294
rect 12124 25230 12126 25282
rect 12178 25230 12180 25282
rect 11452 24946 11844 24948
rect 11452 24894 11454 24946
rect 11506 24894 11844 24946
rect 11452 24892 11844 24894
rect 12124 25060 12180 25230
rect 11452 24882 11508 24892
rect 11228 24658 11284 24668
rect 11564 24722 11620 24734
rect 11564 24670 11566 24722
rect 11618 24670 11620 24722
rect 11564 24612 11620 24670
rect 11452 24500 11508 24510
rect 10892 24498 11508 24500
rect 10892 24446 11454 24498
rect 11506 24446 11508 24498
rect 10892 24444 11508 24446
rect 11452 24434 11508 24444
rect 10872 24332 11136 24342
rect 10928 24276 10976 24332
rect 11032 24276 11080 24332
rect 11564 24276 11620 24556
rect 10872 24266 11136 24276
rect 11340 24220 11620 24276
rect 10668 24108 11172 24164
rect 10108 24070 10164 24108
rect 10556 23938 10612 23950
rect 10556 23886 10558 23938
rect 10610 23886 10612 23938
rect 10556 23828 10612 23886
rect 11004 23940 11060 23950
rect 10556 23762 10612 23772
rect 10668 23826 10724 23838
rect 10668 23774 10670 23826
rect 10722 23774 10724 23826
rect 9660 23604 9716 23660
rect 9996 23650 10052 23660
rect 9660 23538 9716 23548
rect 9884 23268 9940 23278
rect 9884 23266 10052 23268
rect 9884 23214 9886 23266
rect 9938 23214 10052 23266
rect 9884 23212 10052 23214
rect 9884 23202 9940 23212
rect 9772 23154 9828 23166
rect 9772 23102 9774 23154
rect 9826 23102 9828 23154
rect 9324 22932 9380 22942
rect 9324 22370 9380 22876
rect 9772 22708 9828 23102
rect 9772 22642 9828 22652
rect 9884 22930 9940 22942
rect 9884 22878 9886 22930
rect 9938 22878 9940 22930
rect 9436 22484 9492 22494
rect 9436 22390 9492 22428
rect 9772 22484 9828 22494
rect 9324 22318 9326 22370
rect 9378 22318 9380 22370
rect 9324 21924 9380 22318
rect 9324 21858 9380 21868
rect 9436 22260 9492 22270
rect 9212 20188 9268 20636
rect 9324 20916 9380 20926
rect 9324 20690 9380 20860
rect 9324 20638 9326 20690
rect 9378 20638 9380 20690
rect 9324 20626 9380 20638
rect 9212 20132 9380 20188
rect 8540 19394 8596 19404
rect 8316 19346 8484 19348
rect 8316 19294 8318 19346
rect 8370 19294 8484 19346
rect 8316 19292 8484 19294
rect 8316 19216 8372 19292
rect 8316 18788 8372 18798
rect 8316 18450 8372 18732
rect 8316 18398 8318 18450
rect 8370 18398 8372 18450
rect 8316 18386 8372 18398
rect 8428 18452 8484 19292
rect 8540 19234 8596 19246
rect 8540 19182 8542 19234
rect 8594 19182 8596 19234
rect 8540 18676 8596 19182
rect 8876 19236 8932 19246
rect 8876 19142 8932 19180
rect 8876 18676 8932 18686
rect 8540 18620 8820 18676
rect 8652 18452 8708 18462
rect 8428 18450 8708 18452
rect 8428 18398 8654 18450
rect 8706 18398 8708 18450
rect 8428 18396 8708 18398
rect 8652 18386 8708 18396
rect 7868 18340 7924 18350
rect 7868 18246 7924 18284
rect 8764 17892 8820 18620
rect 9324 18676 9380 20132
rect 9436 19796 9492 22204
rect 9772 21810 9828 22428
rect 9884 22036 9940 22878
rect 9996 22260 10052 23212
rect 10108 23156 10164 23166
rect 10108 22594 10164 23100
rect 10108 22542 10110 22594
rect 10162 22542 10164 22594
rect 10108 22530 10164 22542
rect 9996 22194 10052 22204
rect 9884 21980 10052 22036
rect 9772 21758 9774 21810
rect 9826 21758 9828 21810
rect 9772 21746 9828 21758
rect 9884 21812 9940 21822
rect 9996 21812 10052 21980
rect 10220 21812 10276 21822
rect 9996 21810 10276 21812
rect 9996 21758 10222 21810
rect 10274 21758 10276 21810
rect 9996 21756 10276 21758
rect 9884 21700 9940 21756
rect 10220 21746 10276 21756
rect 9884 21644 10052 21700
rect 9996 21586 10052 21644
rect 9996 21534 9998 21586
rect 10050 21534 10052 21586
rect 9996 21522 10052 21534
rect 9884 21476 9940 21486
rect 9884 21382 9940 21420
rect 10668 20804 10724 23774
rect 11004 23826 11060 23884
rect 11004 23774 11006 23826
rect 11058 23774 11060 23826
rect 11004 23762 11060 23774
rect 11116 23938 11172 24108
rect 11116 23886 11118 23938
rect 11170 23886 11172 23938
rect 11116 23604 11172 23886
rect 11116 23538 11172 23548
rect 11228 23940 11284 23950
rect 10872 22764 11136 22774
rect 10928 22708 10976 22764
rect 11032 22708 11080 22764
rect 10872 22698 11136 22708
rect 10872 21196 11136 21206
rect 10928 21140 10976 21196
rect 11032 21140 11080 21196
rect 10872 21130 11136 21140
rect 9884 20692 9940 20702
rect 9884 20598 9940 20636
rect 10556 20692 10612 20702
rect 10668 20672 10724 20748
rect 10780 21028 10836 21038
rect 10556 20598 10612 20636
rect 9548 20578 9604 20590
rect 10332 20580 10388 20590
rect 9548 20526 9550 20578
rect 9602 20526 9604 20578
rect 9548 20188 9604 20526
rect 9996 20578 10388 20580
rect 9996 20526 10334 20578
rect 10386 20526 10388 20578
rect 9996 20524 10388 20526
rect 9548 20132 9940 20188
rect 9884 19906 9940 20132
rect 9884 19854 9886 19906
rect 9938 19854 9940 19906
rect 9436 19740 9828 19796
rect 9436 19460 9492 19470
rect 9436 19366 9492 19404
rect 9660 19236 9716 19246
rect 9660 19142 9716 19180
rect 9772 19012 9828 19740
rect 9884 19460 9940 19854
rect 9884 19394 9940 19404
rect 9884 19236 9940 19246
rect 9996 19236 10052 20524
rect 10332 20514 10388 20524
rect 10780 20468 10836 20972
rect 11116 20916 11172 20926
rect 11228 20916 11284 23884
rect 11340 23828 11396 24220
rect 11340 23378 11396 23772
rect 11340 23326 11342 23378
rect 11394 23326 11396 23378
rect 11340 23314 11396 23326
rect 11676 23828 11732 24892
rect 12012 24836 12068 24846
rect 12012 24612 12068 24780
rect 11900 24556 12012 24612
rect 11788 24052 11844 24062
rect 11788 23958 11844 23996
rect 11676 22596 11732 23772
rect 11676 22530 11732 22540
rect 11116 20914 11284 20916
rect 11116 20862 11118 20914
rect 11170 20862 11284 20914
rect 11116 20860 11284 20862
rect 11116 20692 11172 20860
rect 11564 20804 11620 20814
rect 11564 20710 11620 20748
rect 11116 20626 11172 20636
rect 10780 20188 10836 20412
rect 10108 20132 10164 20142
rect 10108 20038 10164 20076
rect 10668 20132 10836 20188
rect 9884 19234 10052 19236
rect 9884 19182 9886 19234
rect 9938 19182 10052 19234
rect 9884 19180 10052 19182
rect 9884 19170 9940 19180
rect 9996 19012 10052 19022
rect 9772 19010 10052 19012
rect 9772 18958 9998 19010
rect 10050 18958 10052 19010
rect 9772 18956 10052 18958
rect 9996 18946 10052 18956
rect 10108 19012 10164 19022
rect 10108 19010 10276 19012
rect 10108 18958 10110 19010
rect 10162 18958 10276 19010
rect 10108 18956 10276 18958
rect 10108 18946 10164 18956
rect 9884 18676 9940 18686
rect 9324 18620 9828 18676
rect 8876 18582 8932 18620
rect 9772 18562 9828 18620
rect 9884 18582 9940 18620
rect 9772 18510 9774 18562
rect 9826 18510 9828 18562
rect 8764 17826 8820 17836
rect 8988 18450 9044 18462
rect 8988 18398 8990 18450
rect 9042 18398 9044 18450
rect 8988 18340 9044 18398
rect 7980 17780 8036 17790
rect 7532 17666 7588 17678
rect 7532 17614 7534 17666
rect 7586 17614 7588 17666
rect 7532 16324 7588 17614
rect 7868 16882 7924 16894
rect 7868 16830 7870 16882
rect 7922 16830 7924 16882
rect 7756 16324 7812 16334
rect 7532 16322 7812 16324
rect 7532 16270 7758 16322
rect 7810 16270 7812 16322
rect 7532 16268 7812 16270
rect 7756 16258 7812 16268
rect 7420 16212 7476 16222
rect 7476 16156 7700 16212
rect 7420 16146 7476 16156
rect 7644 16098 7700 16156
rect 7644 16046 7646 16098
rect 7698 16046 7700 16098
rect 7644 16034 7700 16046
rect 7756 16100 7812 16110
rect 7756 15986 7812 16044
rect 7756 15934 7758 15986
rect 7810 15934 7812 15986
rect 7756 15922 7812 15934
rect 7756 13636 7812 13646
rect 7756 13542 7812 13580
rect 7868 13188 7924 16830
rect 7980 15204 8036 17724
rect 8428 17780 8484 17790
rect 8484 17724 8596 17780
rect 8428 17714 8484 17724
rect 8540 17556 8596 17724
rect 8876 17668 8932 17678
rect 8876 17574 8932 17612
rect 8540 17462 8596 17500
rect 8652 17442 8708 17454
rect 8652 17390 8654 17442
rect 8706 17390 8708 17442
rect 8652 16772 8708 17390
rect 8988 16772 9044 18284
rect 9548 18452 9604 18462
rect 9548 17778 9604 18396
rect 9772 18228 9828 18510
rect 9772 18162 9828 18172
rect 10108 18450 10164 18462
rect 10108 18398 10110 18450
rect 10162 18398 10164 18450
rect 10108 18340 10164 18398
rect 9548 17726 9550 17778
rect 9602 17726 9604 17778
rect 9548 17714 9604 17726
rect 9660 17892 9716 17902
rect 9660 17666 9716 17836
rect 10108 17890 10164 18284
rect 10108 17838 10110 17890
rect 10162 17838 10164 17890
rect 10108 17826 10164 17838
rect 10220 18452 10276 18956
rect 9660 17614 9662 17666
rect 9714 17614 9716 17666
rect 9660 17602 9716 17614
rect 9772 17666 9828 17678
rect 9772 17614 9774 17666
rect 9826 17614 9828 17666
rect 8652 16770 9044 16772
rect 8652 16718 8990 16770
rect 9042 16718 9044 16770
rect 8652 16716 9044 16718
rect 8988 15876 9044 16716
rect 9436 17442 9492 17454
rect 9436 17390 9438 17442
rect 9490 17390 9492 17442
rect 9436 16100 9492 17390
rect 9772 17106 9828 17614
rect 9772 17054 9774 17106
rect 9826 17054 9828 17106
rect 9772 17042 9828 17054
rect 10220 17668 10276 18396
rect 10556 18676 10612 18686
rect 10444 18338 10500 18350
rect 10444 18286 10446 18338
rect 10498 18286 10500 18338
rect 10444 18228 10500 18286
rect 10444 18162 10500 18172
rect 10556 17778 10612 18620
rect 10556 17726 10558 17778
rect 10610 17726 10612 17778
rect 10556 17714 10612 17726
rect 10220 16884 10276 17612
rect 10332 16884 10388 16894
rect 10220 16882 10388 16884
rect 10220 16830 10334 16882
rect 10386 16830 10388 16882
rect 10220 16828 10388 16830
rect 10332 16818 10388 16828
rect 10108 16660 10164 16670
rect 10108 16658 10276 16660
rect 10108 16606 10110 16658
rect 10162 16606 10276 16658
rect 10108 16604 10276 16606
rect 10108 16594 10164 16604
rect 10220 16322 10276 16604
rect 10220 16270 10222 16322
rect 10274 16270 10276 16322
rect 10220 16258 10276 16270
rect 9660 16100 9716 16110
rect 9436 16098 9716 16100
rect 9436 16046 9662 16098
rect 9714 16046 9716 16098
rect 9436 16044 9716 16046
rect 8988 15810 9044 15820
rect 9212 15988 9268 15998
rect 9212 15874 9268 15932
rect 9212 15822 9214 15874
rect 9266 15822 9268 15874
rect 7980 15138 8036 15148
rect 8540 15314 8596 15326
rect 8540 15262 8542 15314
rect 8594 15262 8596 15314
rect 8540 15204 8596 15262
rect 8540 15138 8596 15148
rect 8988 15204 9044 15214
rect 9212 15204 9268 15822
rect 9660 15428 9716 16044
rect 9996 15988 10052 15998
rect 9996 15894 10052 15932
rect 9884 15876 9940 15886
rect 9884 15782 9940 15820
rect 10444 15876 10500 15886
rect 9660 15362 9716 15372
rect 8988 15202 9268 15204
rect 8988 15150 8990 15202
rect 9042 15150 9268 15202
rect 8988 15148 9268 15150
rect 9660 15204 9716 15214
rect 8092 14530 8148 14542
rect 8092 14478 8094 14530
rect 8146 14478 8148 14530
rect 8092 14420 8148 14478
rect 8092 14354 8148 14364
rect 8652 14530 8708 14542
rect 8652 14478 8654 14530
rect 8706 14478 8708 14530
rect 8652 14420 8708 14478
rect 8764 14532 8820 14542
rect 8764 14438 8820 14476
rect 8652 13858 8708 14364
rect 8652 13806 8654 13858
rect 8706 13806 8708 13858
rect 8652 13794 8708 13806
rect 8204 13748 8260 13758
rect 8204 13654 8260 13692
rect 7868 13122 7924 13132
rect 8988 13076 9044 15148
rect 9660 15110 9716 15148
rect 9436 14756 9492 14766
rect 9436 14642 9492 14700
rect 9436 14590 9438 14642
rect 9490 14590 9492 14642
rect 9436 14578 9492 14590
rect 9996 14530 10052 14542
rect 9996 14478 9998 14530
rect 10050 14478 10052 14530
rect 9324 14420 9380 14430
rect 9324 14326 9380 14364
rect 9548 14308 9604 14318
rect 9548 14214 9604 14252
rect 9884 14308 9940 14318
rect 9884 13970 9940 14252
rect 9884 13918 9886 13970
rect 9938 13918 9940 13970
rect 9772 13746 9828 13758
rect 9772 13694 9774 13746
rect 9826 13694 9828 13746
rect 9772 13636 9828 13694
rect 9884 13748 9940 13918
rect 9884 13682 9940 13692
rect 9772 13570 9828 13580
rect 9884 13524 9940 13534
rect 9996 13524 10052 14478
rect 10444 13860 10500 15820
rect 10444 13794 10500 13804
rect 9884 13522 10052 13524
rect 9884 13470 9886 13522
rect 9938 13470 10052 13522
rect 9884 13468 10052 13470
rect 10220 13636 10276 13646
rect 9884 13458 9940 13468
rect 8428 13074 9044 13076
rect 8428 13022 8990 13074
rect 9042 13022 9044 13074
rect 8428 13020 9044 13022
rect 8428 12850 8484 13020
rect 8988 13010 9044 13020
rect 8428 12798 8430 12850
rect 8482 12798 8484 12850
rect 8428 12786 8484 12798
rect 8540 12850 8596 12862
rect 8540 12798 8542 12850
rect 8594 12798 8596 12850
rect 7252 12684 7364 12740
rect 7756 12740 7812 12750
rect 8204 12740 8260 12750
rect 6524 9156 6580 9166
rect 5964 7858 6020 7868
rect 6188 8034 6244 8046
rect 6188 7982 6190 8034
rect 6242 7982 6244 8034
rect 6188 7924 6244 7982
rect 6188 7858 6244 7868
rect 6524 8036 6580 9100
rect 6748 9044 6804 9054
rect 6748 8950 6804 8988
rect 6636 8036 6692 8046
rect 6524 8034 6692 8036
rect 6524 7982 6638 8034
rect 6690 7982 6692 8034
rect 6524 7980 6692 7982
rect 5516 7700 5572 7710
rect 6300 7700 6356 7710
rect 5516 7698 6356 7700
rect 5516 7646 5518 7698
rect 5570 7646 6302 7698
rect 6354 7646 6356 7698
rect 5516 7644 6356 7646
rect 5516 7634 5572 7644
rect 6300 7634 6356 7644
rect 6412 7588 6468 7598
rect 6412 7494 6468 7532
rect 5628 7476 5684 7486
rect 5404 7474 5684 7476
rect 5404 7422 5630 7474
rect 5682 7422 5684 7474
rect 5404 7420 5684 7422
rect 5628 7410 5684 7420
rect 5740 7476 5796 7486
rect 5740 7382 5796 7420
rect 5628 6468 5684 6478
rect 5180 6466 5684 6468
rect 5180 6414 5630 6466
rect 5682 6414 5684 6466
rect 5180 6412 5684 6414
rect 4508 6290 4564 6300
rect 4732 6356 4788 6366
rect 4620 6020 4676 6030
rect 3836 6018 4676 6020
rect 3836 5966 4622 6018
rect 4674 5966 4676 6018
rect 3836 5964 4676 5966
rect 3836 5906 3892 5964
rect 4620 5954 4676 5964
rect 3836 5854 3838 5906
rect 3890 5854 3892 5906
rect 3836 5842 3892 5854
rect 3612 5630 3614 5682
rect 3666 5630 3668 5682
rect 3612 5618 3668 5630
rect 4508 5236 4564 5246
rect 4732 5236 4788 6300
rect 4508 5234 4788 5236
rect 4508 5182 4510 5234
rect 4562 5182 4788 5234
rect 4508 5180 4788 5182
rect 4508 5170 4564 5180
rect 2940 5122 2996 5134
rect 2940 5070 2942 5122
rect 2994 5070 2996 5122
rect 1932 5012 1988 5022
rect 1596 4386 1652 4396
rect 1820 5010 1988 5012
rect 1820 4958 1934 5010
rect 1986 4958 1988 5010
rect 1820 4956 1988 4958
rect 1820 1540 1876 4956
rect 1932 4946 1988 4956
rect 2940 4564 2996 5070
rect 3836 5124 3892 5134
rect 3836 5030 3892 5068
rect 4844 5124 4900 5134
rect 4844 5030 4900 5068
rect 2940 4498 2996 4508
rect 3052 4900 3108 4910
rect 3052 4338 3108 4844
rect 3612 4900 3668 4910
rect 3612 4806 3668 4844
rect 5068 4788 5124 6412
rect 5628 6020 5684 6412
rect 6076 6466 6132 6478
rect 6076 6414 6078 6466
rect 6130 6414 6132 6466
rect 6076 6356 6132 6414
rect 6076 6290 6132 6300
rect 5628 5954 5684 5964
rect 5404 5908 5460 5918
rect 5404 5814 5460 5852
rect 5068 4722 5124 4732
rect 3612 4564 3668 4574
rect 3612 4470 3668 4508
rect 3948 4452 4004 4462
rect 3948 4358 4004 4396
rect 4508 4452 4564 4462
rect 4508 4358 4564 4396
rect 3052 4286 3054 4338
rect 3106 4286 3108 4338
rect 3052 4274 3108 4286
rect 1932 4226 1988 4238
rect 1932 4174 1934 4226
rect 1986 4174 1988 4226
rect 1932 4004 1988 4174
rect 1932 3938 1988 3948
rect 4956 3668 5012 3678
rect 4956 3574 5012 3612
rect 2156 3556 2212 3566
rect 2156 3462 2212 3500
rect 2716 3556 2772 3566
rect 1820 1474 1876 1484
rect 2716 800 2772 3500
rect 5628 3556 5684 3566
rect 5628 3462 5684 3500
rect 2828 3444 2884 3454
rect 2828 3350 2884 3388
rect 6524 2884 6580 7980
rect 6636 7970 6692 7980
rect 6748 6020 6804 6030
rect 6748 5906 6804 5964
rect 6748 5854 6750 5906
rect 6802 5854 6804 5906
rect 6748 5842 6804 5854
rect 6636 5794 6692 5806
rect 6636 5742 6638 5794
rect 6690 5742 6692 5794
rect 6636 5348 6692 5742
rect 6636 5282 6692 5292
rect 6860 4452 6916 9548
rect 7084 9828 7140 9838
rect 7084 9602 7140 9772
rect 7084 9550 7086 9602
rect 7138 9550 7140 9602
rect 7084 9044 7140 9550
rect 7084 8978 7140 8988
rect 7196 9268 7252 12684
rect 7756 12646 7812 12684
rect 8092 12738 8260 12740
rect 8092 12686 8206 12738
rect 8258 12686 8260 12738
rect 8092 12684 8260 12686
rect 8092 12292 8148 12684
rect 8204 12674 8260 12684
rect 8540 12740 8596 12798
rect 8540 12674 8596 12684
rect 8876 12516 8932 12526
rect 8876 12402 8932 12460
rect 8876 12350 8878 12402
rect 8930 12350 8932 12402
rect 8876 12338 8932 12350
rect 7532 11956 7588 11966
rect 7420 10610 7476 10622
rect 7420 10558 7422 10610
rect 7474 10558 7476 10610
rect 7420 10164 7476 10558
rect 7420 10098 7476 10108
rect 7196 9042 7252 9212
rect 7196 8990 7198 9042
rect 7250 8990 7252 9042
rect 7196 8978 7252 8990
rect 7196 8372 7252 8382
rect 7196 8278 7252 8316
rect 7420 6020 7476 6030
rect 7420 5926 7476 5964
rect 6860 4386 6916 4396
rect 7196 3666 7252 3678
rect 7196 3614 7198 3666
rect 7250 3614 7252 3666
rect 7196 3556 7252 3614
rect 7196 3490 7252 3500
rect 6748 3444 6804 3482
rect 6748 3378 6804 3388
rect 6972 3444 7028 3454
rect 6524 2818 6580 2828
rect 6972 800 7028 3388
rect 7532 3332 7588 11900
rect 7868 10724 7924 10734
rect 7868 10630 7924 10668
rect 7980 10612 8036 10622
rect 7644 10052 7700 10062
rect 7700 9996 7812 10052
rect 7644 9958 7700 9996
rect 7756 9268 7812 9996
rect 7868 9940 7924 9950
rect 7868 9846 7924 9884
rect 7980 9828 8036 10556
rect 7868 9268 7924 9278
rect 7756 9266 7924 9268
rect 7756 9214 7870 9266
rect 7922 9214 7924 9266
rect 7756 9212 7924 9214
rect 7980 9268 8036 9772
rect 8092 9826 8148 12236
rect 8540 12290 8596 12302
rect 8540 12238 8542 12290
rect 8594 12238 8596 12290
rect 8540 10388 8596 12238
rect 8764 12180 8820 12190
rect 8988 12180 9044 12190
rect 8764 12178 8932 12180
rect 8764 12126 8766 12178
rect 8818 12126 8932 12178
rect 8764 12124 8932 12126
rect 8764 12114 8820 12124
rect 8876 11732 8932 12124
rect 8652 11506 8708 11518
rect 8652 11454 8654 11506
rect 8706 11454 8708 11506
rect 8652 10724 8708 11454
rect 8764 11396 8820 11406
rect 8764 10834 8820 11340
rect 8876 11172 8932 11676
rect 8988 11618 9044 12124
rect 9996 12178 10052 12190
rect 9996 12126 9998 12178
rect 10050 12126 10052 12178
rect 8988 11566 8990 11618
rect 9042 11566 9044 11618
rect 8988 11554 9044 11566
rect 9884 12068 9940 12078
rect 8876 11106 8932 11116
rect 8764 10782 8766 10834
rect 8818 10782 8820 10834
rect 8764 10770 8820 10782
rect 8652 10630 8708 10668
rect 8764 10388 8820 10398
rect 8540 10386 8820 10388
rect 8540 10334 8766 10386
rect 8818 10334 8820 10386
rect 8540 10332 8820 10334
rect 8764 10322 8820 10332
rect 8652 10164 8708 10174
rect 8204 9940 8260 9950
rect 8204 9846 8260 9884
rect 8092 9774 8094 9826
rect 8146 9774 8148 9826
rect 8092 9762 8148 9774
rect 8316 9602 8372 9614
rect 8316 9550 8318 9602
rect 8370 9550 8372 9602
rect 8092 9268 8148 9278
rect 7980 9266 8148 9268
rect 7980 9214 8094 9266
rect 8146 9214 8148 9266
rect 7980 9212 8148 9214
rect 7868 9202 7924 9212
rect 8092 9202 8148 9212
rect 8204 9042 8260 9054
rect 8204 8990 8206 9042
rect 8258 8990 8260 9042
rect 8204 8484 8260 8990
rect 8204 8418 8260 8428
rect 7756 8372 7812 8382
rect 7756 8278 7812 8316
rect 7868 8260 7924 8270
rect 7868 7586 7924 8204
rect 8316 8260 8372 9550
rect 8652 9266 8708 10108
rect 8988 10164 9044 10174
rect 8876 9828 8932 9838
rect 8876 9734 8932 9772
rect 8652 9214 8654 9266
rect 8706 9214 8708 9266
rect 8652 9202 8708 9214
rect 8876 9268 8932 9278
rect 8876 9174 8932 9212
rect 8988 9154 9044 10108
rect 8988 9102 8990 9154
rect 9042 9102 9044 9154
rect 7868 7534 7870 7586
rect 7922 7534 7924 7586
rect 7868 7522 7924 7534
rect 8204 8036 8260 8046
rect 8204 6804 8260 7980
rect 8316 7476 8372 8204
rect 8540 9044 8596 9054
rect 8428 7476 8484 7486
rect 8316 7474 8484 7476
rect 8316 7422 8430 7474
rect 8482 7422 8484 7474
rect 8316 7420 8484 7422
rect 8428 7410 8484 7420
rect 8428 6804 8484 6814
rect 7980 6802 8484 6804
rect 7980 6750 8430 6802
rect 8482 6750 8484 6802
rect 7980 6748 8484 6750
rect 7644 5236 7700 5246
rect 7644 5142 7700 5180
rect 7980 5236 8036 6748
rect 8428 6738 8484 6748
rect 8540 6132 8596 8988
rect 8988 8596 9044 9102
rect 9436 9602 9492 9614
rect 9436 9550 9438 9602
rect 9490 9550 9492 9602
rect 9436 8932 9492 9550
rect 9772 9602 9828 9614
rect 9772 9550 9774 9602
rect 9826 9550 9828 9602
rect 9772 9268 9828 9550
rect 9772 9202 9828 9212
rect 9660 8932 9716 8942
rect 9436 8930 9716 8932
rect 9436 8878 9662 8930
rect 9714 8878 9716 8930
rect 9436 8876 9716 8878
rect 8652 8540 9044 8596
rect 8652 8372 8708 8540
rect 8652 8306 8708 8316
rect 8876 8372 8932 8382
rect 8876 8260 8932 8316
rect 9660 8372 9716 8876
rect 9884 8708 9940 12012
rect 9996 11732 10052 12126
rect 10108 12180 10164 12190
rect 10108 12066 10164 12124
rect 10108 12014 10110 12066
rect 10162 12014 10164 12066
rect 10108 12002 10164 12014
rect 9996 11666 10052 11676
rect 10220 10164 10276 13580
rect 10668 11060 10724 20132
rect 11676 20130 11732 20142
rect 11676 20078 11678 20130
rect 11730 20078 11732 20130
rect 10872 19628 11136 19638
rect 10928 19572 10976 19628
rect 11032 19572 11080 19628
rect 10872 19562 11136 19572
rect 11452 18564 11508 18574
rect 11340 18340 11396 18350
rect 11340 18246 11396 18284
rect 10872 18060 11136 18070
rect 10928 18004 10976 18060
rect 11032 18004 11080 18060
rect 10872 17994 11136 18004
rect 10872 16492 11136 16502
rect 10928 16436 10976 16492
rect 11032 16436 11080 16492
rect 10872 16426 11136 16436
rect 11004 16324 11060 16334
rect 11452 16324 11508 18508
rect 11564 18562 11620 18574
rect 11564 18510 11566 18562
rect 11618 18510 11620 18562
rect 11564 18452 11620 18510
rect 11564 18386 11620 18396
rect 11676 17892 11732 20078
rect 11676 17826 11732 17836
rect 11788 17556 11844 17566
rect 11788 17462 11844 17500
rect 11900 17108 11956 24556
rect 12012 24546 12068 24556
rect 12124 24052 12180 25004
rect 12124 23986 12180 23996
rect 12236 24276 12292 24286
rect 12236 24050 12292 24220
rect 12236 23998 12238 24050
rect 12290 23998 12292 24050
rect 12236 23986 12292 23998
rect 12124 22596 12180 22606
rect 12124 22482 12180 22540
rect 12124 22430 12126 22482
rect 12178 22430 12180 22482
rect 12124 22418 12180 22430
rect 12348 22260 12404 27692
rect 12684 27746 12740 27758
rect 12684 27694 12686 27746
rect 12738 27694 12740 27746
rect 12460 26852 12516 26862
rect 12684 26852 12740 27694
rect 13244 27748 13300 27806
rect 12908 26964 12964 26974
rect 12460 26850 12740 26852
rect 12460 26798 12462 26850
rect 12514 26798 12740 26850
rect 12460 26796 12740 26798
rect 12796 26852 12852 26862
rect 12460 26404 12516 26796
rect 12796 26516 12852 26796
rect 12908 26852 12964 26908
rect 13244 26852 13300 27692
rect 12908 26850 13300 26852
rect 12908 26798 12910 26850
rect 12962 26798 13300 26850
rect 12908 26796 13300 26798
rect 12908 26786 12964 26796
rect 12908 26516 12964 26526
rect 12796 26460 12908 26516
rect 12908 26384 12964 26460
rect 12460 26338 12516 26348
rect 12460 26180 12516 26190
rect 12460 24948 12516 26124
rect 12572 25282 12628 25294
rect 12572 25230 12574 25282
rect 12626 25230 12628 25282
rect 12572 25172 12628 25230
rect 12572 25106 12628 25116
rect 12908 25172 12964 25182
rect 12460 24882 12516 24892
rect 12908 24050 12964 25116
rect 13244 24948 13300 26796
rect 13356 27970 13412 27982
rect 13356 27918 13358 27970
rect 13410 27918 13412 27970
rect 13356 26404 13412 27918
rect 13580 27860 13636 27870
rect 13580 27766 13636 27804
rect 13692 26964 13748 26974
rect 13692 26870 13748 26908
rect 13804 26852 13860 28140
rect 13916 28082 13972 28364
rect 13916 28030 13918 28082
rect 13970 28030 13972 28082
rect 13916 28018 13972 28030
rect 14028 28196 14084 28206
rect 14028 27636 14084 28140
rect 14588 28196 14644 28590
rect 14588 28130 14644 28140
rect 14700 28084 14756 28094
rect 14812 28084 14868 28700
rect 14700 28082 14868 28084
rect 14700 28030 14702 28082
rect 14754 28030 14868 28082
rect 14700 28028 14868 28030
rect 15036 28084 15092 29262
rect 15372 29986 15428 29998
rect 15372 29934 15374 29986
rect 15426 29934 15428 29986
rect 15372 29092 15428 29934
rect 15484 29988 15540 29998
rect 15484 29538 15540 29932
rect 16044 29986 16100 30942
rect 16156 31668 16212 31678
rect 16156 31554 16212 31612
rect 16156 31502 16158 31554
rect 16210 31502 16212 31554
rect 16156 30324 16212 31502
rect 16604 31220 16660 36092
rect 16716 35586 16772 36318
rect 16716 35534 16718 35586
rect 16770 35534 16772 35586
rect 16716 35522 16772 35534
rect 17276 35700 17332 36428
rect 17500 36418 17556 36428
rect 17724 36482 17780 36494
rect 17724 36430 17726 36482
rect 17778 36430 17780 36482
rect 17276 35026 17332 35644
rect 17276 34974 17278 35026
rect 17330 34974 17332 35026
rect 17276 34962 17332 34974
rect 17724 35028 17780 36430
rect 17948 36482 18004 36494
rect 17948 36430 17950 36482
rect 18002 36430 18004 36482
rect 17948 36372 18004 36430
rect 17948 36306 18004 36316
rect 18060 36370 18116 36382
rect 18060 36318 18062 36370
rect 18114 36318 18116 36370
rect 17836 35812 17892 35822
rect 17836 35718 17892 35756
rect 18060 35700 18116 36318
rect 18060 35634 18116 35644
rect 18508 36372 18564 36382
rect 16828 34914 16884 34926
rect 16828 34862 16830 34914
rect 16882 34862 16884 34914
rect 16828 34356 16884 34862
rect 16828 34290 16884 34300
rect 16940 34244 16996 34254
rect 16940 34150 16996 34188
rect 17724 34242 17780 34972
rect 18172 34692 18228 34702
rect 17836 34356 17892 34366
rect 17836 34262 17892 34300
rect 17724 34190 17726 34242
rect 17778 34190 17780 34242
rect 17724 34178 17780 34190
rect 17948 34242 18004 34254
rect 17948 34190 17950 34242
rect 18002 34190 18004 34242
rect 17948 33796 18004 34190
rect 18172 33908 18228 34636
rect 18508 34356 18564 36316
rect 18732 36258 18788 36270
rect 18732 36206 18734 36258
rect 18786 36206 18788 36258
rect 18732 35140 18788 36206
rect 18844 36260 18900 37324
rect 18956 36596 19012 39200
rect 19292 36596 19348 36606
rect 18956 36594 19348 36596
rect 18956 36542 19294 36594
rect 19346 36542 19348 36594
rect 18956 36540 19348 36542
rect 21420 36596 21476 39200
rect 21644 36596 21700 36606
rect 21420 36594 21700 36596
rect 21420 36542 21646 36594
rect 21698 36542 21700 36594
rect 21420 36540 21700 36542
rect 19292 36530 19348 36540
rect 21644 36530 21700 36540
rect 21868 36596 21924 36606
rect 18844 35698 18900 36204
rect 20412 36482 20468 36494
rect 20412 36430 20414 36482
rect 20466 36430 20468 36482
rect 18844 35646 18846 35698
rect 18898 35646 18900 35698
rect 18844 35634 18900 35646
rect 19628 35700 19684 35710
rect 19516 35588 19572 35598
rect 18732 35074 18788 35084
rect 18956 35586 19572 35588
rect 18956 35534 19518 35586
rect 19570 35534 19572 35586
rect 18956 35532 19572 35534
rect 18956 34914 19012 35532
rect 19516 35522 19572 35532
rect 19516 35028 19572 35038
rect 19628 35028 19684 35644
rect 19516 35026 19684 35028
rect 19516 34974 19518 35026
rect 19570 34974 19684 35026
rect 19516 34972 19684 34974
rect 19740 35698 19796 35710
rect 19740 35646 19742 35698
rect 19794 35646 19796 35698
rect 19740 35140 19796 35646
rect 19964 35700 20020 35710
rect 19964 35606 20020 35644
rect 19516 34962 19572 34972
rect 18956 34862 18958 34914
rect 19010 34862 19012 34914
rect 18956 34850 19012 34862
rect 19740 34916 19796 35084
rect 20076 35140 20132 35150
rect 20076 35046 20132 35084
rect 20412 35028 20468 36430
rect 20532 36092 20796 36102
rect 20588 36036 20636 36092
rect 20692 36036 20740 36092
rect 20532 36026 20796 36036
rect 21532 35586 21588 35598
rect 21532 35534 21534 35586
rect 21586 35534 21588 35586
rect 21532 35252 21588 35534
rect 21532 35186 21588 35196
rect 20412 34962 20468 34972
rect 21868 35026 21924 36540
rect 22764 36596 22820 36606
rect 22764 36482 22820 36540
rect 23884 36594 23940 39200
rect 26348 37940 26404 39200
rect 28812 37940 28868 39200
rect 26348 37884 26740 37940
rect 28812 37884 29428 37940
rect 23884 36542 23886 36594
rect 23938 36542 23940 36594
rect 23884 36530 23940 36542
rect 24892 37828 24948 37838
rect 24892 36596 24948 37772
rect 22764 36430 22766 36482
rect 22818 36430 22820 36482
rect 22764 36418 22820 36430
rect 24556 36484 24612 36494
rect 24556 36390 24612 36428
rect 23884 36372 23940 36382
rect 23212 35924 23268 35934
rect 21868 34974 21870 35026
rect 21922 34974 21924 35026
rect 21868 34962 21924 34974
rect 21980 35698 22036 35710
rect 21980 35646 21982 35698
rect 22034 35646 22036 35698
rect 19740 34850 19796 34860
rect 20524 34916 20580 34926
rect 20524 34822 20580 34860
rect 18620 34804 18676 34814
rect 18620 34710 18676 34748
rect 20532 34524 20796 34534
rect 20588 34468 20636 34524
rect 20692 34468 20740 34524
rect 20532 34458 20796 34468
rect 18620 34356 18676 34366
rect 18508 34354 18676 34356
rect 18508 34302 18622 34354
rect 18674 34302 18676 34354
rect 18508 34300 18676 34302
rect 18620 34290 18676 34300
rect 18844 34356 18900 34366
rect 18844 34354 19124 34356
rect 18844 34302 18846 34354
rect 18898 34302 19124 34354
rect 18844 34300 19124 34302
rect 18844 34290 18900 34300
rect 18172 33842 18228 33852
rect 18956 34130 19012 34142
rect 18956 34078 18958 34130
rect 19010 34078 19012 34130
rect 17948 33730 18004 33740
rect 17276 33684 17332 33694
rect 17276 33458 17332 33628
rect 17276 33406 17278 33458
rect 17330 33406 17332 33458
rect 17276 33394 17332 33406
rect 17612 33684 17668 33694
rect 17612 32786 17668 33628
rect 17836 33516 18228 33572
rect 17836 32788 17892 33516
rect 17612 32734 17614 32786
rect 17666 32734 17668 32786
rect 17612 32722 17668 32734
rect 17724 32786 17892 32788
rect 17724 32734 17838 32786
rect 17890 32734 17892 32786
rect 17724 32732 17892 32734
rect 16604 31154 16660 31164
rect 16940 31890 16996 31902
rect 16940 31838 16942 31890
rect 16994 31838 16996 31890
rect 16940 31106 16996 31838
rect 17724 31890 17780 32732
rect 17836 32722 17892 32732
rect 17948 33346 18004 33358
rect 17948 33294 17950 33346
rect 18002 33294 18004 33346
rect 17948 32674 18004 33294
rect 18172 33346 18228 33516
rect 18172 33294 18174 33346
rect 18226 33294 18228 33346
rect 18172 33282 18228 33294
rect 17948 32622 17950 32674
rect 18002 32622 18004 32674
rect 17948 31948 18004 32622
rect 18844 33236 18900 33246
rect 18956 33236 19012 34078
rect 18844 33234 19012 33236
rect 18844 33182 18846 33234
rect 18898 33182 19012 33234
rect 18844 33180 19012 33182
rect 18844 32562 18900 33180
rect 18844 32510 18846 32562
rect 18898 32510 18900 32562
rect 18844 32498 18900 32510
rect 19068 32564 19124 34300
rect 21196 34244 21252 34254
rect 20076 34130 20132 34142
rect 20076 34078 20078 34130
rect 20130 34078 20132 34130
rect 20076 33684 20132 34078
rect 21196 34130 21252 34188
rect 21980 34244 22036 35646
rect 22428 35700 22484 35710
rect 22428 35606 22484 35644
rect 22988 35588 23044 35598
rect 22652 35252 22708 35262
rect 22652 35138 22708 35196
rect 22652 35086 22654 35138
rect 22706 35086 22708 35138
rect 22652 35074 22708 35086
rect 22988 35138 23044 35532
rect 22988 35086 22990 35138
rect 23042 35086 23044 35138
rect 22988 35074 23044 35086
rect 23100 35586 23156 35598
rect 23100 35534 23102 35586
rect 23154 35534 23156 35586
rect 23100 35140 23156 35534
rect 23100 35074 23156 35084
rect 22428 34802 22484 34814
rect 22428 34750 22430 34802
rect 22482 34750 22484 34802
rect 22428 34244 22484 34750
rect 21980 34242 22484 34244
rect 21980 34190 21982 34242
rect 22034 34190 22484 34242
rect 21980 34188 22484 34190
rect 21980 34178 22036 34188
rect 21196 34078 21198 34130
rect 21250 34078 21252 34130
rect 21196 34066 21252 34078
rect 20188 34018 20244 34030
rect 20188 33966 20190 34018
rect 20242 33966 20244 34018
rect 20188 33908 20244 33966
rect 22988 34018 23044 34030
rect 22988 33966 22990 34018
rect 23042 33966 23044 34018
rect 20188 33842 20244 33852
rect 21980 33908 22036 33918
rect 20188 33684 20244 33694
rect 20076 33628 20188 33684
rect 19740 33346 19796 33358
rect 19740 33294 19742 33346
rect 19794 33294 19796 33346
rect 19740 32674 19796 33294
rect 20188 33348 20244 33628
rect 21980 33460 22036 33852
rect 22988 33908 23044 33966
rect 22988 33842 23044 33852
rect 22764 33684 22820 33694
rect 22428 33460 22484 33470
rect 21980 33458 22484 33460
rect 21980 33406 21982 33458
rect 22034 33406 22430 33458
rect 22482 33406 22484 33458
rect 21980 33404 22484 33406
rect 21980 33394 22036 33404
rect 22428 33394 22484 33404
rect 22764 33458 22820 33628
rect 22764 33406 22766 33458
rect 22818 33406 22820 33458
rect 22764 33394 22820 33406
rect 20412 33348 20468 33358
rect 20188 33346 20468 33348
rect 20188 33294 20414 33346
rect 20466 33294 20468 33346
rect 20188 33292 20468 33294
rect 19964 33124 20020 33134
rect 19964 33030 20020 33068
rect 19740 32622 19742 32674
rect 19794 32622 19796 32674
rect 19740 32610 19796 32622
rect 19068 32432 19124 32508
rect 17948 31892 18676 31948
rect 17724 31838 17726 31890
rect 17778 31838 17780 31890
rect 17724 31826 17780 31838
rect 17052 31778 17108 31790
rect 17052 31726 17054 31778
rect 17106 31726 17108 31778
rect 17052 31332 17108 31726
rect 17052 31266 17108 31276
rect 18620 31218 18676 31892
rect 20188 31444 20244 33292
rect 20412 33282 20468 33292
rect 20532 32956 20796 32966
rect 20588 32900 20636 32956
rect 20692 32900 20740 32956
rect 20532 32890 20796 32900
rect 22652 32676 22708 32686
rect 22652 32582 22708 32620
rect 20300 32564 20356 32574
rect 20300 31890 20356 32508
rect 22428 32562 22484 32574
rect 22428 32510 22430 32562
rect 22482 32510 22484 32562
rect 22428 31948 22484 32510
rect 22428 31892 22596 31948
rect 22652 31892 22708 31902
rect 20300 31838 20302 31890
rect 20354 31838 20356 31890
rect 20300 31826 20356 31838
rect 22540 31890 22708 31892
rect 22540 31838 22654 31890
rect 22706 31838 22708 31890
rect 22540 31836 22708 31838
rect 22652 31826 22708 31836
rect 20636 31780 20692 31790
rect 20188 31378 20244 31388
rect 20412 31724 20636 31780
rect 18620 31166 18622 31218
rect 18674 31166 18676 31218
rect 18620 31154 18676 31166
rect 20412 31220 20468 31724
rect 20636 31686 20692 31724
rect 20860 31778 20916 31790
rect 20860 31726 20862 31778
rect 20914 31726 20916 31778
rect 20860 31668 20916 31726
rect 21756 31780 21812 31790
rect 21756 31686 21812 31724
rect 21980 31778 22036 31790
rect 21980 31726 21982 31778
rect 22034 31726 22036 31778
rect 20532 31388 20796 31398
rect 20588 31332 20636 31388
rect 20692 31332 20740 31388
rect 20532 31322 20796 31332
rect 20412 31164 20692 31220
rect 16940 31054 16942 31106
rect 16994 31054 16996 31106
rect 16940 31042 16996 31054
rect 20636 31106 20692 31164
rect 20636 31054 20638 31106
rect 20690 31054 20692 31106
rect 20636 31042 20692 31054
rect 18508 30996 18564 31006
rect 18732 30996 18788 31006
rect 18508 30994 18676 30996
rect 18508 30942 18510 30994
rect 18562 30942 18676 30994
rect 18508 30940 18676 30942
rect 18508 30930 18564 30940
rect 16716 30884 16772 30894
rect 16604 30324 16660 30334
rect 16716 30324 16772 30828
rect 17612 30884 17668 30894
rect 17612 30436 17668 30828
rect 18620 30660 18676 30940
rect 18732 30902 18788 30940
rect 19180 30996 19236 31006
rect 19964 30996 20020 31006
rect 19180 30994 19460 30996
rect 19180 30942 19182 30994
rect 19234 30942 19460 30994
rect 19180 30940 19460 30942
rect 19180 30930 19236 30940
rect 19180 30660 19236 30670
rect 18620 30604 19180 30660
rect 17612 30370 17668 30380
rect 18732 30436 18788 30446
rect 16156 30322 16772 30324
rect 16156 30270 16606 30322
rect 16658 30270 16772 30322
rect 16156 30268 16772 30270
rect 16156 30210 16212 30268
rect 16604 30258 16660 30268
rect 16156 30158 16158 30210
rect 16210 30158 16212 30210
rect 16156 30146 16212 30158
rect 16044 29934 16046 29986
rect 16098 29934 16100 29986
rect 16044 29652 16100 29934
rect 17164 29986 17220 29998
rect 17164 29934 17166 29986
rect 17218 29934 17220 29986
rect 16044 29586 16100 29596
rect 16380 29652 16436 29662
rect 16380 29558 16436 29596
rect 17164 29652 17220 29934
rect 15484 29486 15486 29538
rect 15538 29486 15540 29538
rect 15484 29474 15540 29486
rect 15372 29026 15428 29036
rect 15484 28980 15540 28990
rect 15372 28644 15428 28654
rect 15372 28550 15428 28588
rect 15036 28028 15204 28084
rect 14700 28018 14756 28028
rect 14140 27970 14196 27982
rect 14140 27918 14142 27970
rect 14194 27918 14196 27970
rect 14140 27860 14196 27918
rect 14924 27972 14980 27982
rect 14924 27878 14980 27916
rect 14140 27794 14196 27804
rect 14252 27860 14308 27870
rect 15036 27860 15092 27870
rect 14252 27858 14868 27860
rect 14252 27806 14254 27858
rect 14306 27806 14868 27858
rect 14252 27804 14868 27806
rect 14252 27794 14308 27804
rect 14028 27074 14084 27580
rect 14028 27022 14030 27074
rect 14082 27022 14084 27074
rect 14028 27010 14084 27022
rect 14252 27300 14308 27310
rect 13804 26796 14084 26852
rect 13804 26628 13860 26638
rect 13580 26516 13636 26526
rect 13580 26422 13636 26460
rect 13804 26514 13860 26572
rect 13804 26462 13806 26514
rect 13858 26462 13860 26514
rect 13804 26450 13860 26462
rect 13356 26338 13412 26348
rect 13692 26404 13748 26414
rect 13692 26310 13748 26348
rect 13916 26292 13972 26302
rect 13916 26198 13972 26236
rect 13244 24882 13300 24892
rect 14028 24836 14084 26796
rect 14252 26850 14308 27244
rect 14812 27074 14868 27804
rect 15036 27766 15092 27804
rect 15148 27300 15204 28028
rect 14812 27022 14814 27074
rect 14866 27022 14868 27074
rect 14812 27010 14868 27022
rect 14924 27244 15204 27300
rect 15260 27972 15316 27982
rect 14364 26964 14420 26974
rect 14364 26870 14420 26908
rect 14252 26798 14254 26850
rect 14306 26798 14308 26850
rect 14140 26290 14196 26302
rect 14140 26238 14142 26290
rect 14194 26238 14196 26290
rect 14140 26180 14196 26238
rect 14140 26114 14196 26124
rect 14252 25284 14308 26798
rect 14924 26628 14980 27244
rect 15148 26964 15204 26974
rect 15148 26870 15204 26908
rect 15036 26850 15092 26862
rect 15036 26798 15038 26850
rect 15090 26798 15092 26850
rect 15036 26740 15092 26798
rect 15260 26740 15316 27916
rect 15484 26908 15540 28924
rect 16940 28418 16996 28430
rect 16940 28366 16942 28418
rect 16994 28366 16996 28418
rect 15596 27746 15652 27758
rect 15596 27694 15598 27746
rect 15650 27694 15652 27746
rect 15596 27300 15652 27694
rect 15596 27234 15652 27244
rect 15932 27746 15988 27758
rect 15932 27694 15934 27746
rect 15986 27694 15988 27746
rect 15036 26684 15316 26740
rect 14924 26572 15092 26628
rect 14812 26290 14868 26302
rect 14812 26238 14814 26290
rect 14866 26238 14868 26290
rect 14700 26180 14756 26190
rect 14588 25956 14644 25966
rect 14252 25228 14532 25284
rect 14252 24836 14308 24846
rect 14028 24834 14308 24836
rect 14028 24782 14254 24834
rect 14306 24782 14308 24834
rect 14028 24780 14308 24782
rect 14252 24770 14308 24780
rect 13020 24724 13076 24734
rect 13020 24630 13076 24668
rect 13580 24722 13636 24734
rect 13580 24670 13582 24722
rect 13634 24670 13636 24722
rect 12908 23998 12910 24050
rect 12962 23998 12964 24050
rect 12908 23940 12964 23998
rect 13580 23940 13636 24670
rect 13692 24724 13748 24734
rect 13692 24630 13748 24668
rect 14364 24724 14420 24734
rect 14364 24630 14420 24668
rect 14476 24164 14532 25228
rect 13916 24108 14532 24164
rect 13692 23940 13748 23950
rect 13580 23938 13748 23940
rect 13580 23886 13694 23938
rect 13746 23886 13748 23938
rect 13580 23884 13748 23886
rect 12908 23874 12964 23884
rect 13692 23874 13748 23884
rect 13916 23826 13972 24108
rect 14476 24050 14532 24108
rect 14476 23998 14478 24050
rect 14530 23998 14532 24050
rect 14476 23986 14532 23998
rect 14028 23940 14084 23950
rect 14028 23846 14084 23884
rect 14588 23828 14644 25900
rect 14700 25618 14756 26124
rect 14812 25956 14868 26238
rect 14812 25890 14868 25900
rect 14700 25566 14702 25618
rect 14754 25566 14756 25618
rect 14700 25554 14756 25566
rect 14924 24722 14980 24734
rect 14924 24670 14926 24722
rect 14978 24670 14980 24722
rect 14924 24612 14980 24670
rect 14924 24546 14980 24556
rect 13916 23774 13918 23826
rect 13970 23774 13972 23826
rect 13916 23762 13972 23774
rect 14252 23772 14644 23828
rect 13468 23156 13524 23166
rect 13468 23062 13524 23100
rect 13916 23156 13972 23166
rect 13020 23044 13076 23054
rect 12796 23042 13076 23044
rect 12796 22990 13022 23042
rect 13074 22990 13076 23042
rect 12796 22988 13076 22990
rect 12684 22820 12740 22830
rect 12572 22596 12628 22606
rect 12572 22502 12628 22540
rect 12348 22204 12628 22260
rect 12572 21698 12628 22204
rect 12572 21646 12574 21698
rect 12626 21646 12628 21698
rect 12572 21634 12628 21646
rect 12012 20580 12068 20590
rect 12012 20130 12068 20524
rect 12012 20078 12014 20130
rect 12066 20078 12068 20130
rect 12012 20066 12068 20078
rect 12348 18228 12404 18238
rect 11900 17106 12180 17108
rect 11900 17054 11902 17106
rect 11954 17054 12180 17106
rect 11900 17052 12180 17054
rect 11900 17042 11956 17052
rect 12012 16658 12068 16670
rect 12012 16606 12014 16658
rect 12066 16606 12068 16658
rect 11004 16322 11508 16324
rect 11004 16270 11006 16322
rect 11058 16270 11508 16322
rect 11004 16268 11508 16270
rect 11004 16258 11060 16268
rect 11340 16100 11396 16110
rect 11340 16006 11396 16044
rect 11452 16098 11508 16268
rect 11900 16324 11956 16334
rect 12012 16324 12068 16606
rect 11900 16322 12068 16324
rect 11900 16270 11902 16322
rect 11954 16270 12068 16322
rect 11900 16268 12068 16270
rect 11900 16258 11956 16268
rect 11452 16046 11454 16098
rect 11506 16046 11508 16098
rect 11452 16034 11508 16046
rect 11564 16098 11620 16110
rect 11564 16046 11566 16098
rect 11618 16046 11620 16098
rect 11228 15876 11284 15886
rect 11228 15782 11284 15820
rect 11564 15538 11620 16046
rect 12124 15988 12180 17052
rect 12348 17106 12404 18172
rect 12460 17892 12516 17902
rect 12460 17798 12516 17836
rect 12572 17556 12628 17566
rect 12572 17462 12628 17500
rect 12460 17444 12516 17454
rect 12460 17350 12516 17388
rect 12348 17054 12350 17106
rect 12402 17054 12404 17106
rect 12348 16996 12404 17054
rect 12348 16930 12404 16940
rect 12684 16212 12740 22764
rect 12796 22260 12852 22988
rect 13020 22978 13076 22988
rect 13356 22708 13412 22718
rect 12908 22482 12964 22494
rect 12908 22430 12910 22482
rect 12962 22430 12964 22482
rect 12908 22372 12964 22430
rect 12908 22306 12964 22316
rect 12796 22128 12852 22204
rect 13020 21586 13076 21598
rect 13020 21534 13022 21586
rect 13074 21534 13076 21586
rect 13020 20580 13076 21534
rect 13356 20916 13412 22652
rect 13804 22484 13860 22494
rect 13804 22390 13860 22428
rect 13692 22372 13748 22382
rect 13692 22278 13748 22316
rect 13916 22370 13972 23100
rect 13916 22318 13918 22370
rect 13970 22318 13972 22370
rect 13916 22306 13972 22318
rect 13916 22148 13972 22158
rect 13468 21476 13524 21486
rect 13468 21474 13748 21476
rect 13468 21422 13470 21474
rect 13522 21422 13748 21474
rect 13468 21420 13748 21422
rect 13468 21410 13524 21420
rect 13356 20850 13412 20860
rect 13020 20514 13076 20524
rect 13692 20802 13748 21420
rect 13804 20916 13860 20926
rect 13916 20916 13972 22092
rect 13804 20914 13972 20916
rect 13804 20862 13806 20914
rect 13858 20862 13972 20914
rect 13804 20860 13972 20862
rect 13804 20850 13860 20860
rect 13692 20750 13694 20802
rect 13746 20750 13748 20802
rect 13020 20132 13076 20142
rect 12796 17444 12852 17454
rect 12796 17106 12852 17388
rect 12796 17054 12798 17106
rect 12850 17054 12852 17106
rect 12796 17042 12852 17054
rect 12124 15922 12180 15932
rect 12460 16156 12740 16212
rect 11564 15486 11566 15538
rect 11618 15486 11620 15538
rect 11564 15474 11620 15486
rect 11900 15876 11956 15886
rect 11004 15428 11060 15438
rect 11004 15314 11060 15372
rect 11004 15262 11006 15314
rect 11058 15262 11060 15314
rect 11004 15250 11060 15262
rect 11228 15204 11284 15214
rect 11228 15110 11284 15148
rect 10872 14924 11136 14934
rect 10928 14868 10976 14924
rect 11032 14868 11080 14924
rect 10872 14858 11136 14868
rect 11452 13748 11508 13758
rect 11452 13654 11508 13692
rect 11900 13748 11956 15820
rect 12348 15876 12404 15886
rect 12348 15782 12404 15820
rect 12348 15204 12404 15214
rect 12348 14532 12404 15148
rect 12460 14756 12516 16156
rect 12572 15988 12628 15998
rect 12572 15894 12628 15932
rect 12684 15986 12740 15998
rect 12684 15934 12686 15986
rect 12738 15934 12740 15986
rect 12684 15652 12740 15934
rect 12684 15586 12740 15596
rect 12908 15876 12964 15886
rect 12684 15428 12740 15466
rect 12684 15362 12740 15372
rect 12460 14690 12516 14700
rect 12460 14532 12516 14542
rect 12348 14530 12516 14532
rect 12348 14478 12462 14530
rect 12514 14478 12516 14530
rect 12348 14476 12516 14478
rect 12460 14466 12516 14476
rect 12572 14530 12628 14542
rect 12908 14532 12964 15820
rect 13020 15148 13076 20076
rect 13692 19794 13748 20750
rect 14028 20692 14084 20702
rect 13916 20580 13972 20590
rect 13916 20486 13972 20524
rect 13916 19908 13972 19918
rect 13916 19814 13972 19852
rect 13692 19742 13694 19794
rect 13746 19742 13748 19794
rect 13692 19730 13748 19742
rect 13804 19460 13860 19470
rect 13804 19234 13860 19404
rect 13804 19182 13806 19234
rect 13858 19182 13860 19234
rect 13804 19170 13860 19182
rect 13244 18564 13300 18574
rect 13300 18508 13636 18564
rect 13244 18432 13300 18508
rect 13468 18340 13524 18350
rect 13468 18246 13524 18284
rect 13580 17666 13636 18508
rect 14028 18450 14084 20636
rect 14252 20132 14308 23772
rect 15036 23266 15092 26572
rect 15260 26516 15316 26684
rect 15148 26404 15204 26414
rect 15148 25620 15204 26348
rect 15260 26290 15316 26460
rect 15260 26238 15262 26290
rect 15314 26238 15316 26290
rect 15260 26180 15316 26238
rect 15260 26114 15316 26124
rect 15372 26852 15540 26908
rect 15596 26852 15652 26862
rect 15932 26852 15988 27694
rect 16492 27746 16548 27758
rect 16492 27694 16494 27746
rect 16546 27694 16548 27746
rect 16492 27636 16548 27694
rect 16492 27188 16548 27580
rect 16940 27300 16996 28366
rect 16828 27298 16996 27300
rect 16828 27246 16942 27298
rect 16994 27246 16996 27298
rect 16828 27244 16996 27246
rect 16828 27188 16884 27244
rect 16940 27234 16996 27244
rect 17052 27746 17108 27758
rect 17052 27694 17054 27746
rect 17106 27694 17108 27746
rect 16492 27122 16548 27132
rect 16604 27132 16884 27188
rect 17052 27188 17108 27694
rect 15148 25526 15204 25564
rect 15036 23214 15038 23266
rect 15090 23214 15092 23266
rect 15036 23202 15092 23214
rect 14812 23154 14868 23166
rect 14812 23102 14814 23154
rect 14866 23102 14868 23154
rect 14812 22596 14868 23102
rect 14812 22484 14868 22540
rect 14812 22428 15092 22484
rect 14364 22372 14420 22382
rect 14700 22372 14756 22382
rect 14364 22370 14756 22372
rect 14364 22318 14366 22370
rect 14418 22318 14702 22370
rect 14754 22318 14756 22370
rect 14364 22316 14756 22318
rect 14364 22306 14420 22316
rect 14700 22306 14756 22316
rect 14924 22260 14980 22270
rect 14924 22166 14980 22204
rect 15036 22258 15092 22428
rect 15036 22206 15038 22258
rect 15090 22206 15092 22258
rect 15036 22148 15092 22206
rect 15036 22092 15316 22148
rect 15260 21474 15316 22092
rect 15260 21422 15262 21474
rect 15314 21422 15316 21474
rect 15260 21028 15316 21422
rect 15372 21476 15428 26852
rect 15596 26850 15988 26852
rect 15596 26798 15598 26850
rect 15650 26798 15988 26850
rect 16156 26964 16212 26974
rect 16212 26908 16324 26964
rect 16156 26832 16212 26908
rect 15596 26796 15988 26798
rect 15596 26786 15652 26796
rect 15932 26516 15988 26796
rect 15932 26450 15988 26460
rect 16156 26404 16212 26414
rect 16044 26292 16100 26302
rect 15708 26178 15764 26190
rect 15708 26126 15710 26178
rect 15762 26126 15764 26178
rect 15708 25956 15764 26126
rect 15708 25890 15764 25900
rect 16044 25396 16100 26236
rect 16156 26178 16212 26348
rect 16156 26126 16158 26178
rect 16210 26126 16212 26178
rect 16156 25620 16212 26126
rect 16156 25554 16212 25564
rect 16044 25340 16212 25396
rect 15932 25284 15988 25294
rect 15932 24946 15988 25228
rect 15932 24894 15934 24946
rect 15986 24894 15988 24946
rect 15932 24882 15988 24894
rect 15820 24724 15876 24734
rect 15820 24630 15876 24668
rect 16044 24722 16100 24734
rect 16044 24670 16046 24722
rect 16098 24670 16100 24722
rect 16044 24612 16100 24670
rect 15932 24500 15988 24510
rect 15372 21410 15428 21420
rect 15484 22146 15540 22158
rect 15484 22094 15486 22146
rect 15538 22094 15540 22146
rect 15484 21028 15540 22094
rect 15260 20972 15540 21028
rect 14364 20804 14420 20814
rect 14364 20802 14868 20804
rect 14364 20750 14366 20802
rect 14418 20750 14868 20802
rect 14364 20748 14868 20750
rect 14364 20738 14420 20748
rect 14812 20242 14868 20748
rect 14812 20190 14814 20242
rect 14866 20190 14868 20242
rect 14812 20178 14868 20190
rect 14252 20066 14308 20076
rect 15036 20130 15092 20142
rect 15036 20078 15038 20130
rect 15090 20078 15092 20130
rect 14140 20020 14196 20030
rect 14140 19926 14196 19964
rect 15036 20020 15092 20078
rect 14252 19572 14308 19582
rect 14252 19346 14308 19516
rect 14252 19294 14254 19346
rect 14306 19294 14308 19346
rect 14252 18676 14308 19294
rect 14700 19460 14756 19470
rect 14700 19346 14756 19404
rect 14700 19294 14702 19346
rect 14754 19294 14756 19346
rect 14700 19282 14756 19294
rect 15036 19348 15092 19964
rect 15036 19282 15092 19292
rect 15148 20018 15204 20030
rect 15148 19966 15150 20018
rect 15202 19966 15204 20018
rect 15148 19908 15204 19966
rect 15148 18788 15204 19852
rect 15148 18722 15204 18732
rect 14252 18610 14308 18620
rect 14028 18398 14030 18450
rect 14082 18398 14084 18450
rect 14028 18386 14084 18398
rect 14476 18450 14532 18462
rect 14476 18398 14478 18450
rect 14530 18398 14532 18450
rect 13580 17614 13582 17666
rect 13634 17614 13636 17666
rect 13580 17602 13636 17614
rect 14364 17668 14420 17678
rect 13916 17554 13972 17566
rect 13916 17502 13918 17554
rect 13970 17502 13972 17554
rect 13804 17444 13860 17454
rect 13916 17444 13972 17502
rect 14364 17444 14420 17612
rect 13916 17442 14420 17444
rect 13916 17390 14366 17442
rect 14418 17390 14420 17442
rect 13916 17388 14420 17390
rect 13468 17108 13524 17118
rect 13468 17014 13524 17052
rect 13580 16996 13636 17006
rect 13636 16940 13748 16996
rect 13580 16902 13636 16940
rect 13244 16882 13300 16894
rect 13244 16830 13246 16882
rect 13298 16830 13300 16882
rect 13132 16660 13188 16670
rect 13244 16660 13300 16830
rect 13132 16658 13300 16660
rect 13132 16606 13134 16658
rect 13186 16606 13300 16658
rect 13132 16604 13300 16606
rect 13132 16594 13188 16604
rect 13244 15314 13300 16604
rect 13692 16100 13748 16940
rect 13804 16884 13860 17388
rect 14140 16884 14196 16894
rect 13804 16882 14196 16884
rect 13804 16830 14142 16882
rect 14194 16830 14196 16882
rect 13804 16828 14196 16830
rect 13244 15262 13246 15314
rect 13298 15262 13300 15314
rect 13244 15250 13300 15262
rect 13356 16044 13748 16100
rect 13020 15092 13188 15148
rect 12572 14478 12574 14530
rect 12626 14478 12628 14530
rect 12236 14420 12292 14430
rect 12236 14326 12292 14364
rect 12348 14308 12404 14318
rect 12348 14214 12404 14252
rect 12572 14084 12628 14478
rect 12012 14028 12628 14084
rect 12796 14530 12964 14532
rect 12796 14478 12910 14530
rect 12962 14478 12964 14530
rect 12796 14476 12964 14478
rect 12012 13970 12068 14028
rect 12012 13918 12014 13970
rect 12066 13918 12068 13970
rect 12012 13906 12068 13918
rect 11900 13682 11956 13692
rect 12124 13860 12180 13870
rect 11676 13524 11732 13534
rect 11676 13430 11732 13468
rect 10872 13356 11136 13366
rect 10928 13300 10976 13356
rect 11032 13300 11080 13356
rect 10872 13290 11136 13300
rect 11788 12738 11844 12750
rect 11788 12686 11790 12738
rect 11842 12686 11844 12738
rect 11788 12292 11844 12686
rect 11788 12198 11844 12236
rect 10780 11956 10836 11994
rect 10780 11890 10836 11900
rect 10872 11788 11136 11798
rect 10928 11732 10976 11788
rect 11032 11732 11080 11788
rect 10872 11722 11136 11732
rect 12012 11172 12068 11182
rect 12124 11172 12180 13804
rect 12796 13634 12852 14476
rect 12908 14466 12964 14476
rect 12908 13858 12964 13870
rect 12908 13806 12910 13858
rect 12962 13806 12964 13858
rect 12908 13748 12964 13806
rect 12908 13682 12964 13692
rect 12796 13582 12798 13634
rect 12850 13582 12852 13634
rect 12796 13570 12852 13582
rect 12348 13076 12404 13086
rect 12348 12982 12404 13020
rect 12348 12852 12404 12862
rect 12348 12290 12404 12796
rect 13020 12852 13076 12862
rect 12796 12738 12852 12750
rect 12796 12686 12798 12738
rect 12850 12686 12852 12738
rect 12348 12238 12350 12290
rect 12402 12238 12404 12290
rect 12348 12226 12404 12238
rect 12460 12292 12516 12302
rect 12460 12198 12516 12236
rect 12796 12292 12852 12686
rect 12796 12226 12852 12236
rect 12684 12180 12740 12190
rect 12684 12086 12740 12124
rect 12908 11956 12964 11966
rect 12012 11170 12180 11172
rect 12012 11118 12014 11170
rect 12066 11118 12180 11170
rect 12012 11116 12180 11118
rect 12460 11170 12516 11182
rect 12460 11118 12462 11170
rect 12514 11118 12516 11170
rect 10668 11004 11508 11060
rect 10556 10836 10612 10846
rect 11340 10836 11396 10846
rect 10556 10834 11396 10836
rect 10556 10782 10558 10834
rect 10610 10782 11342 10834
rect 11394 10782 11396 10834
rect 10556 10780 11396 10782
rect 10556 10770 10612 10780
rect 11340 10770 11396 10780
rect 11116 10610 11172 10622
rect 11116 10558 11118 10610
rect 11170 10558 11172 10610
rect 10220 10098 10276 10108
rect 10444 10498 10500 10510
rect 10444 10446 10446 10498
rect 10498 10446 10500 10498
rect 10444 9940 10500 10446
rect 11116 10388 11172 10558
rect 11228 10612 11284 10650
rect 11228 10546 11284 10556
rect 11116 10332 11396 10388
rect 10872 10220 11136 10230
rect 10928 10164 10976 10220
rect 11032 10164 11080 10220
rect 10872 10154 11136 10164
rect 10444 9874 10500 9884
rect 11004 9940 11060 9950
rect 11004 9826 11060 9884
rect 11004 9774 11006 9826
rect 11058 9774 11060 9826
rect 11004 9762 11060 9774
rect 11340 9938 11396 10332
rect 11340 9886 11342 9938
rect 11394 9886 11396 9938
rect 10556 9492 10612 9502
rect 9884 8642 9940 8652
rect 10444 9044 10500 9054
rect 10444 8930 10500 8988
rect 10444 8878 10446 8930
rect 10498 8878 10500 8930
rect 10444 8596 10500 8878
rect 10444 8530 10500 8540
rect 9660 8306 9716 8316
rect 8764 8258 8932 8260
rect 8764 8206 8878 8258
rect 8930 8206 8932 8258
rect 8764 8204 8932 8206
rect 8652 7362 8708 7374
rect 8652 7310 8654 7362
rect 8706 7310 8708 7362
rect 8652 6692 8708 7310
rect 8652 6626 8708 6636
rect 8540 6066 8596 6076
rect 8652 6468 8708 6478
rect 8428 6020 8484 6030
rect 8428 5906 8484 5964
rect 8428 5854 8430 5906
rect 8482 5854 8484 5906
rect 8428 5842 8484 5854
rect 8652 5908 8708 6412
rect 8652 5776 8708 5852
rect 8652 5348 8708 5358
rect 8652 5254 8708 5292
rect 8764 5236 8820 8204
rect 8876 8194 8932 8204
rect 9324 8258 9380 8270
rect 9324 8206 9326 8258
rect 9378 8206 9380 8258
rect 9324 8148 9380 8206
rect 9772 8260 9828 8270
rect 9772 8166 9828 8204
rect 9324 6916 9380 8092
rect 10108 8146 10164 8158
rect 10108 8094 10110 8146
rect 10162 8094 10164 8146
rect 9996 8036 10052 8046
rect 9996 7942 10052 7980
rect 10108 7924 10164 8094
rect 10108 7858 10164 7868
rect 9884 7700 9940 7710
rect 10444 7700 10500 7710
rect 10556 7700 10612 9436
rect 10892 9156 10948 9166
rect 10892 9042 10948 9100
rect 11340 9154 11396 9886
rect 11340 9102 11342 9154
rect 11394 9102 11396 9154
rect 11340 9090 11396 9102
rect 10892 8990 10894 9042
rect 10946 8990 10948 9042
rect 10892 8978 10948 8990
rect 10872 8652 11136 8662
rect 10928 8596 10976 8652
rect 11032 8596 11080 8652
rect 10872 8586 11136 8596
rect 10668 8036 10724 8046
rect 11004 8036 11060 8046
rect 10668 7812 10724 7980
rect 10668 7746 10724 7756
rect 10892 8034 11060 8036
rect 10892 7982 11006 8034
rect 11058 7982 11060 8034
rect 10892 7980 11060 7982
rect 10892 7924 10948 7980
rect 11004 7970 11060 7980
rect 9884 7698 10612 7700
rect 9884 7646 9886 7698
rect 9938 7646 10446 7698
rect 10498 7646 10612 7698
rect 9884 7644 10612 7646
rect 10892 7698 10948 7868
rect 10892 7646 10894 7698
rect 10946 7646 10948 7698
rect 9884 7634 9940 7644
rect 9324 6850 9380 6860
rect 9772 7588 9828 7626
rect 9660 6804 9716 6814
rect 9324 6692 9380 6702
rect 9324 6598 9380 6636
rect 9660 6690 9716 6748
rect 9660 6638 9662 6690
rect 9714 6638 9716 6690
rect 9660 6626 9716 6638
rect 9436 6580 9492 6590
rect 8876 6466 8932 6478
rect 8876 6414 8878 6466
rect 8930 6414 8932 6466
rect 8876 6132 8932 6414
rect 8876 6066 8932 6076
rect 9436 6020 9492 6524
rect 8988 5796 9044 5806
rect 8988 5702 9044 5740
rect 7980 5234 8596 5236
rect 7980 5182 7982 5234
rect 8034 5182 8596 5234
rect 7980 5180 8596 5182
rect 7980 5170 8036 5180
rect 8540 5012 8596 5180
rect 8652 5012 8708 5022
rect 8540 5010 8708 5012
rect 8540 4958 8654 5010
rect 8706 4958 8708 5010
rect 8540 4956 8708 4958
rect 8652 4946 8708 4956
rect 8764 5010 8820 5180
rect 9324 5236 9380 5246
rect 9436 5236 9492 5964
rect 9324 5234 9492 5236
rect 9324 5182 9326 5234
rect 9378 5182 9492 5234
rect 9324 5180 9492 5182
rect 9548 6466 9604 6478
rect 9548 6414 9550 6466
rect 9602 6414 9604 6466
rect 9548 6132 9604 6414
rect 9324 5170 9380 5180
rect 8764 4958 8766 5010
rect 8818 4958 8820 5010
rect 8764 4946 8820 4958
rect 8652 4340 8708 4350
rect 8652 4246 8708 4284
rect 9100 4228 9156 4238
rect 9100 4134 9156 4172
rect 8204 3444 8260 3482
rect 8204 3378 8260 3388
rect 9100 3444 9156 3454
rect 7532 3266 7588 3276
rect 9100 800 9156 3388
rect 9548 1092 9604 6076
rect 9772 5908 9828 7532
rect 9884 7250 9940 7262
rect 9884 7198 9886 7250
rect 9938 7198 9940 7250
rect 9884 6580 9940 7198
rect 9884 6514 9940 6524
rect 9996 6804 10052 7644
rect 10444 7634 10500 7644
rect 10892 7634 10948 7646
rect 10872 7084 11136 7094
rect 10928 7028 10976 7084
rect 11032 7028 11080 7084
rect 10872 7018 11136 7028
rect 9996 6244 10052 6748
rect 10220 6692 10276 6702
rect 10108 6468 10164 6478
rect 10108 6374 10164 6412
rect 9996 6178 10052 6188
rect 9660 5852 9828 5908
rect 9884 6132 9940 6142
rect 9660 5124 9716 5852
rect 9772 5682 9828 5694
rect 9772 5630 9774 5682
rect 9826 5630 9828 5682
rect 9772 5348 9828 5630
rect 9772 5282 9828 5292
rect 9884 5234 9940 6076
rect 10220 6130 10276 6636
rect 10444 6692 10500 6702
rect 10444 6598 10500 6636
rect 10892 6692 10948 6702
rect 10892 6598 10948 6636
rect 10220 6078 10222 6130
rect 10274 6078 10276 6130
rect 10220 6066 10276 6078
rect 10332 6468 10388 6478
rect 10332 6020 10388 6412
rect 11340 6468 11396 6478
rect 11340 6374 11396 6412
rect 11116 6244 11172 6254
rect 10444 6132 10500 6142
rect 10444 6038 10500 6076
rect 11116 6130 11172 6188
rect 11116 6078 11118 6130
rect 11170 6078 11172 6130
rect 11116 6066 11172 6078
rect 10332 5954 10388 5964
rect 9996 5796 10052 5806
rect 9996 5702 10052 5740
rect 10332 5794 10388 5806
rect 10332 5742 10334 5794
rect 10386 5742 10388 5794
rect 9884 5182 9886 5234
rect 9938 5182 9940 5234
rect 9884 5170 9940 5182
rect 9996 5124 10052 5134
rect 9660 5068 9828 5124
rect 9660 3668 9716 3678
rect 9660 3554 9716 3612
rect 9660 3502 9662 3554
rect 9714 3502 9716 3554
rect 9660 3490 9716 3502
rect 9772 2660 9828 5068
rect 9884 4452 9940 4462
rect 9996 4452 10052 5068
rect 10332 5124 10388 5742
rect 10872 5516 11136 5526
rect 10928 5460 10976 5516
rect 11032 5460 11080 5516
rect 10872 5450 11136 5460
rect 10332 5058 10388 5068
rect 10556 5234 10612 5246
rect 10556 5182 10558 5234
rect 10610 5182 10612 5234
rect 9884 4450 10052 4452
rect 9884 4398 9886 4450
rect 9938 4398 10052 4450
rect 9884 4396 10052 4398
rect 10556 4450 10612 5182
rect 10668 5124 10724 5134
rect 10668 5030 10724 5068
rect 11340 5012 11396 5022
rect 10556 4398 10558 4450
rect 10610 4398 10612 4450
rect 9884 4386 9940 4396
rect 9996 4114 10052 4126
rect 9996 4062 9998 4114
rect 10050 4062 10052 4114
rect 9996 3556 10052 4062
rect 9996 3490 10052 3500
rect 10332 3666 10388 3678
rect 10332 3614 10334 3666
rect 10386 3614 10388 3666
rect 10332 3444 10388 3614
rect 10556 3668 10612 4398
rect 10780 5010 11396 5012
rect 10780 4958 11342 5010
rect 11394 4958 11396 5010
rect 10780 4956 11396 4958
rect 10780 4228 10836 4956
rect 11340 4946 11396 4956
rect 11452 4564 11508 11004
rect 11676 10610 11732 10622
rect 11676 10558 11678 10610
rect 11730 10558 11732 10610
rect 11676 10052 11732 10558
rect 12012 10500 12068 11116
rect 12460 10724 12516 11118
rect 12908 10948 12964 11900
rect 13020 11506 13076 12796
rect 13020 11454 13022 11506
rect 13074 11454 13076 11506
rect 13020 11442 13076 11454
rect 13132 10948 13188 15092
rect 13356 13076 13412 16044
rect 13692 15988 13748 16044
rect 13916 16212 13972 16222
rect 13916 16098 13972 16156
rect 13916 16046 13918 16098
rect 13970 16046 13972 16098
rect 13916 16034 13972 16046
rect 13804 15988 13860 15998
rect 13692 15986 13860 15988
rect 13692 15934 13806 15986
rect 13858 15934 13860 15986
rect 13692 15932 13860 15934
rect 13804 15922 13860 15932
rect 13580 15876 13636 15886
rect 13580 15782 13636 15820
rect 13580 15652 13636 15662
rect 13580 14532 13636 15596
rect 13916 15314 13972 15326
rect 13916 15262 13918 15314
rect 13970 15262 13972 15314
rect 13804 15204 13860 15214
rect 13916 15204 13972 15262
rect 13860 15148 13972 15204
rect 14140 15148 14196 16828
rect 14252 15316 14308 17388
rect 14364 17378 14420 17388
rect 14476 17444 14532 18398
rect 15260 18338 15316 18350
rect 15260 18286 15262 18338
rect 15314 18286 15316 18338
rect 14476 17378 14532 17388
rect 14588 18116 14644 18126
rect 14588 17108 14644 18060
rect 15260 18116 15316 18286
rect 15372 18228 15428 20972
rect 15820 18564 15876 18574
rect 15820 18470 15876 18508
rect 15372 18162 15428 18172
rect 14812 17444 14868 17454
rect 14812 17350 14868 17388
rect 14588 17014 14644 17052
rect 14812 16996 14868 17006
rect 14364 16212 14420 16222
rect 14364 16118 14420 16156
rect 14812 16210 14868 16940
rect 15260 16772 15316 18060
rect 15932 17780 15988 24444
rect 16044 22930 16100 24556
rect 16044 22878 16046 22930
rect 16098 22878 16100 22930
rect 16044 22866 16100 22878
rect 16156 22260 16212 25340
rect 16268 24836 16324 26908
rect 16604 26404 16660 27132
rect 17052 27122 17108 27132
rect 16716 26964 16772 26974
rect 17052 26964 17108 26974
rect 16716 26962 17108 26964
rect 16716 26910 16718 26962
rect 16770 26910 17054 26962
rect 17106 26910 17108 26962
rect 16716 26908 17108 26910
rect 16716 26898 16772 26908
rect 17052 26740 17108 26908
rect 17052 26674 17108 26684
rect 16716 26404 16772 26414
rect 16604 26402 16772 26404
rect 16604 26350 16718 26402
rect 16770 26350 16772 26402
rect 16604 26348 16772 26350
rect 16716 26338 16772 26348
rect 16828 26404 16884 26414
rect 16828 26310 16884 26348
rect 17052 26292 17108 26302
rect 17052 26198 17108 26236
rect 17164 26180 17220 29596
rect 18284 29540 18340 29550
rect 18284 29446 18340 29484
rect 18060 29428 18116 29438
rect 17724 29426 18116 29428
rect 17724 29374 18062 29426
rect 18114 29374 18116 29426
rect 17724 29372 18116 29374
rect 17724 28642 17780 29372
rect 18060 29362 18116 29372
rect 18396 29428 18452 29438
rect 18396 29426 18676 29428
rect 18396 29374 18398 29426
rect 18450 29374 18676 29426
rect 18396 29372 18676 29374
rect 18396 29362 18452 29372
rect 17836 28756 17892 28766
rect 17836 28662 17892 28700
rect 18620 28754 18676 29372
rect 18620 28702 18622 28754
rect 18674 28702 18676 28754
rect 17724 28590 17726 28642
rect 17778 28590 17780 28642
rect 17724 28578 17780 28590
rect 18620 28644 18676 28702
rect 18620 28578 18676 28588
rect 17388 28532 17444 28542
rect 17388 28438 17444 28476
rect 17948 28530 18004 28542
rect 17948 28478 17950 28530
rect 18002 28478 18004 28530
rect 17612 28420 17668 28430
rect 17164 26114 17220 26124
rect 17388 27298 17444 27310
rect 17388 27246 17390 27298
rect 17442 27246 17444 27298
rect 17388 25284 17444 27246
rect 17500 27076 17556 27086
rect 17500 26404 17556 27020
rect 17500 26338 17556 26348
rect 16268 24770 16324 24780
rect 17276 25282 17444 25284
rect 17276 25230 17390 25282
rect 17442 25230 17444 25282
rect 17276 25228 17444 25230
rect 16492 24722 16548 24734
rect 16492 24670 16494 24722
rect 16546 24670 16548 24722
rect 15932 17714 15988 17724
rect 16044 22204 16212 22260
rect 16380 23042 16436 23054
rect 16380 22990 16382 23042
rect 16434 22990 16436 23042
rect 16380 22370 16436 22990
rect 16492 22594 16548 24670
rect 17276 23714 17332 25228
rect 17388 25218 17444 25228
rect 17612 24276 17668 28364
rect 17948 28420 18004 28478
rect 17948 28354 18004 28364
rect 18284 28420 18340 28430
rect 18284 28082 18340 28364
rect 18284 28030 18286 28082
rect 18338 28030 18340 28082
rect 18284 28018 18340 28030
rect 17724 27746 17780 27758
rect 17724 27694 17726 27746
rect 17778 27694 17780 27746
rect 17724 27298 17780 27694
rect 17948 27636 18004 27646
rect 17948 27542 18004 27580
rect 17724 27246 17726 27298
rect 17778 27246 17780 27298
rect 17724 27234 17780 27246
rect 18060 26962 18116 26974
rect 18060 26910 18062 26962
rect 18114 26910 18116 26962
rect 18060 26740 18116 26910
rect 18732 26908 18788 30380
rect 19180 30434 19236 30604
rect 19180 30382 19182 30434
rect 19234 30382 19236 30434
rect 19180 30370 19236 30382
rect 19292 30322 19348 30334
rect 19292 30270 19294 30322
rect 19346 30270 19348 30322
rect 18956 30210 19012 30222
rect 18956 30158 18958 30210
rect 19010 30158 19012 30210
rect 18060 26674 18116 26684
rect 18172 26852 18228 26862
rect 18172 26404 18228 26796
rect 18172 26338 18228 26348
rect 18396 26850 18452 26862
rect 18396 26798 18398 26850
rect 18450 26798 18452 26850
rect 18396 26402 18452 26798
rect 18620 26852 18788 26908
rect 18844 29540 18900 29550
rect 18844 28642 18900 29484
rect 18956 29314 19012 30158
rect 18956 29262 18958 29314
rect 19010 29262 19012 29314
rect 18956 28756 19012 29262
rect 19180 29204 19236 29214
rect 19292 29204 19348 30270
rect 19404 29652 19460 30940
rect 19964 30902 20020 30940
rect 19740 30882 19796 30894
rect 19740 30830 19742 30882
rect 19794 30830 19796 30882
rect 19740 30660 19796 30830
rect 19740 30594 19796 30604
rect 20532 29820 20796 29830
rect 20588 29764 20636 29820
rect 20692 29764 20740 29820
rect 20532 29754 20796 29764
rect 19516 29652 19572 29662
rect 19404 29650 19572 29652
rect 19404 29598 19518 29650
rect 19570 29598 19572 29650
rect 19404 29596 19572 29598
rect 19516 29586 19572 29596
rect 20860 29316 20916 31612
rect 21980 31668 22036 31726
rect 21980 31602 22036 31612
rect 22876 30884 22932 30894
rect 22876 30882 23044 30884
rect 22876 30830 22878 30882
rect 22930 30830 23044 30882
rect 22876 30828 23044 30830
rect 22876 30818 22932 30828
rect 22988 29988 23044 30828
rect 22988 29894 23044 29932
rect 21308 29538 21364 29550
rect 21308 29486 21310 29538
rect 21362 29486 21364 29538
rect 21308 29428 21364 29486
rect 21196 29316 21252 29326
rect 20860 29314 21252 29316
rect 20860 29262 21198 29314
rect 21250 29262 21252 29314
rect 20860 29260 21252 29262
rect 21196 29250 21252 29260
rect 19180 29202 19348 29204
rect 19180 29150 19182 29202
rect 19234 29150 19348 29202
rect 19180 29148 19348 29150
rect 19180 29138 19236 29148
rect 18956 28690 19012 28700
rect 18844 28590 18846 28642
rect 18898 28590 18900 28642
rect 18844 27858 18900 28590
rect 19180 28644 19236 28654
rect 19068 28532 19124 28542
rect 19068 28082 19124 28476
rect 19068 28030 19070 28082
rect 19122 28030 19124 28082
rect 19068 28018 19124 28030
rect 18844 27806 18846 27858
rect 18898 27806 18900 27858
rect 18844 26852 18900 27806
rect 19180 27970 19236 28588
rect 19180 27918 19182 27970
rect 19234 27918 19236 27970
rect 19180 27524 19236 27918
rect 18956 27468 19236 27524
rect 18956 27298 19012 27468
rect 18956 27246 18958 27298
rect 19010 27246 19012 27298
rect 18956 27234 19012 27246
rect 19068 27076 19124 27086
rect 19068 26982 19124 27020
rect 19292 26908 19348 29148
rect 20860 28756 20916 28766
rect 21308 28756 21364 29372
rect 22428 29428 22484 29438
rect 22428 29334 22484 29372
rect 23100 29428 23156 29438
rect 23100 29334 23156 29372
rect 21532 29316 21588 29326
rect 21532 29222 21588 29260
rect 22204 29316 22260 29326
rect 22204 29222 22260 29260
rect 22876 29316 22932 29326
rect 20860 28754 21364 28756
rect 20860 28702 20862 28754
rect 20914 28702 21364 28754
rect 20860 28700 21364 28702
rect 21756 29204 21812 29214
rect 20860 28690 20916 28700
rect 20188 28642 20244 28654
rect 20188 28590 20190 28642
rect 20242 28590 20244 28642
rect 20188 28420 20244 28590
rect 20188 28354 20244 28364
rect 21196 28308 21252 28318
rect 20532 28252 20796 28262
rect 20588 28196 20636 28252
rect 20692 28196 20740 28252
rect 20532 28186 20796 28196
rect 19740 27746 19796 27758
rect 19740 27694 19742 27746
rect 19794 27694 19796 27746
rect 19740 26908 19796 27694
rect 20076 27746 20132 27758
rect 20076 27694 20078 27746
rect 20130 27694 20132 27746
rect 19964 27076 20020 27086
rect 20076 27076 20132 27694
rect 19964 27074 20132 27076
rect 19964 27022 19966 27074
rect 20018 27022 20132 27074
rect 19964 27020 20132 27022
rect 19964 27010 20020 27020
rect 20076 26964 20132 27020
rect 20524 27746 20580 27758
rect 20524 27694 20526 27746
rect 20578 27694 20580 27746
rect 18396 26350 18398 26402
rect 18450 26350 18452 26402
rect 18396 26338 18452 26350
rect 18508 26404 18564 26414
rect 17948 26292 18004 26302
rect 17948 26178 18004 26236
rect 17948 26126 17950 26178
rect 18002 26126 18004 26178
rect 17948 25506 18004 26126
rect 18284 26180 18340 26190
rect 18284 25730 18340 26124
rect 18284 25678 18286 25730
rect 18338 25678 18340 25730
rect 18284 25666 18340 25678
rect 17948 25454 17950 25506
rect 18002 25454 18004 25506
rect 17948 25442 18004 25454
rect 18396 25508 18452 25518
rect 18396 25414 18452 25452
rect 18508 25284 18564 26348
rect 17612 24210 17668 24220
rect 18396 25228 18564 25284
rect 17724 24052 17780 24062
rect 18396 24052 18452 25228
rect 18620 24834 18676 26852
rect 18844 26786 18900 26796
rect 18956 26850 19012 26862
rect 19292 26852 19572 26908
rect 18956 26798 18958 26850
rect 19010 26798 19012 26850
rect 18956 26740 19012 26798
rect 18956 26674 19012 26684
rect 19516 26516 19572 26852
rect 19628 26852 19684 26862
rect 19740 26852 19908 26908
rect 20076 26898 20132 26908
rect 20412 26964 20468 26974
rect 19628 26740 19684 26796
rect 19852 26850 19908 26852
rect 19852 26798 19854 26850
rect 19906 26798 19908 26850
rect 19628 26684 19796 26740
rect 19628 26516 19684 26526
rect 19516 26514 19684 26516
rect 19516 26462 19630 26514
rect 19682 26462 19684 26514
rect 19516 26460 19684 26462
rect 19628 26450 19684 26460
rect 19516 26292 19572 26302
rect 19516 26198 19572 26236
rect 19292 25620 19348 25630
rect 19292 25526 19348 25564
rect 19404 25508 19460 25518
rect 19740 25508 19796 26684
rect 19852 26404 19908 26798
rect 19852 26338 19908 26348
rect 20188 26292 20244 26302
rect 20188 25508 20244 26236
rect 19404 25506 19796 25508
rect 19404 25454 19406 25506
rect 19458 25454 19796 25506
rect 19404 25452 19796 25454
rect 19964 25506 20244 25508
rect 19964 25454 20190 25506
rect 20242 25454 20244 25506
rect 19964 25452 20244 25454
rect 19404 25442 19460 25452
rect 18620 24782 18622 24834
rect 18674 24782 18676 24834
rect 18620 24770 18676 24782
rect 17724 24050 18452 24052
rect 17724 23998 17726 24050
rect 17778 23998 18452 24050
rect 17724 23996 18452 23998
rect 17724 23986 17780 23996
rect 17276 23662 17278 23714
rect 17330 23662 17332 23714
rect 17276 23492 17332 23662
rect 18284 23826 18340 23838
rect 18284 23774 18286 23826
rect 18338 23774 18340 23826
rect 16492 22542 16494 22594
rect 16546 22542 16548 22594
rect 16492 22530 16548 22542
rect 16604 23154 16660 23166
rect 16604 23102 16606 23154
rect 16658 23102 16660 23154
rect 16380 22318 16382 22370
rect 16434 22318 16436 22370
rect 15260 16706 15316 16716
rect 15372 17332 15428 17342
rect 14812 16158 14814 16210
rect 14866 16158 14868 16210
rect 14812 16146 14868 16158
rect 15148 16324 15204 16334
rect 14588 15988 14644 15998
rect 14476 15540 14532 15550
rect 14476 15446 14532 15484
rect 14252 15250 14308 15260
rect 13804 14754 13860 15148
rect 13804 14702 13806 14754
rect 13858 14702 13860 14754
rect 13804 14690 13860 14702
rect 14028 15092 14196 15148
rect 13692 14532 13748 14542
rect 13580 14530 13748 14532
rect 13580 14478 13694 14530
rect 13746 14478 13748 14530
rect 13580 14476 13748 14478
rect 13356 13010 13412 13020
rect 13468 14420 13524 14430
rect 13468 12290 13524 14364
rect 13692 13076 13748 14476
rect 13804 14420 13860 14430
rect 14028 14420 14084 15092
rect 13804 14418 14084 14420
rect 13804 14366 13806 14418
rect 13858 14366 14084 14418
rect 13804 14364 14084 14366
rect 14364 14420 14420 14430
rect 13804 14354 13860 14364
rect 13804 13524 13860 13534
rect 13804 13186 13860 13468
rect 13804 13134 13806 13186
rect 13858 13134 13860 13186
rect 13804 13122 13860 13134
rect 13692 13010 13748 13020
rect 13692 12852 13748 12862
rect 13468 12238 13470 12290
rect 13522 12238 13524 12290
rect 13468 12226 13524 12238
rect 13580 12850 13748 12852
rect 13580 12798 13694 12850
rect 13746 12798 13748 12850
rect 13580 12796 13748 12798
rect 13580 11844 13636 12796
rect 13692 12786 13748 12796
rect 13804 12852 13860 12862
rect 13916 12852 13972 14364
rect 14364 14326 14420 14364
rect 14588 14420 14644 15932
rect 15148 15876 15204 16268
rect 15260 15876 15316 15886
rect 15148 15874 15316 15876
rect 15148 15822 15262 15874
rect 15314 15822 15316 15874
rect 15148 15820 15316 15822
rect 15148 15764 15204 15820
rect 15260 15810 15316 15820
rect 15148 15698 15204 15708
rect 15260 15540 15316 15550
rect 15372 15540 15428 17276
rect 15708 16882 15764 16894
rect 15708 16830 15710 16882
rect 15762 16830 15764 16882
rect 15708 16772 15764 16830
rect 15708 16100 15764 16716
rect 15708 16034 15764 16044
rect 15932 15876 15988 15886
rect 15260 15538 15372 15540
rect 15260 15486 15262 15538
rect 15314 15486 15372 15538
rect 15260 15484 15372 15486
rect 15260 15474 15316 15484
rect 15372 15408 15428 15484
rect 15708 15820 15932 15876
rect 15708 15538 15764 15820
rect 15932 15782 15988 15820
rect 15708 15486 15710 15538
rect 15762 15486 15764 15538
rect 14812 14868 14868 14878
rect 14588 14326 14644 14364
rect 14700 14418 14756 14430
rect 14700 14366 14702 14418
rect 14754 14366 14756 14418
rect 14700 14308 14756 14366
rect 14700 14242 14756 14252
rect 14812 13858 14868 14812
rect 15596 14420 15652 14430
rect 15596 14326 15652 14364
rect 15148 14308 15204 14318
rect 15204 14252 15316 14308
rect 15148 14176 15204 14252
rect 14812 13806 14814 13858
rect 14866 13806 14868 13858
rect 14812 13794 14868 13806
rect 15260 13860 15316 14252
rect 15708 13860 15764 15486
rect 16044 15092 16100 22204
rect 16156 21588 16212 21598
rect 16156 21474 16212 21532
rect 16156 21422 16158 21474
rect 16210 21422 16212 21474
rect 16156 19572 16212 21422
rect 16380 21026 16436 22318
rect 16492 22260 16548 22270
rect 16604 22260 16660 23102
rect 16548 22204 16660 22260
rect 16492 22166 16548 22204
rect 17164 22148 17220 22158
rect 17276 22148 17332 23436
rect 18060 23604 18116 23614
rect 18060 23378 18116 23548
rect 18284 23492 18340 23774
rect 18396 23826 18452 23996
rect 19180 24722 19236 24734
rect 19852 24724 19908 24734
rect 19180 24670 19182 24722
rect 19234 24670 19236 24722
rect 18620 23940 18676 23950
rect 18620 23846 18676 23884
rect 18396 23774 18398 23826
rect 18450 23774 18452 23826
rect 18396 23762 18452 23774
rect 19180 23492 19236 24670
rect 19292 24722 19908 24724
rect 19292 24670 19854 24722
rect 19906 24670 19908 24722
rect 19292 24668 19908 24670
rect 19292 24162 19348 24668
rect 19852 24658 19908 24668
rect 19964 24500 20020 25452
rect 20188 25442 20244 25452
rect 20300 25620 20356 25630
rect 19292 24110 19294 24162
rect 19346 24110 19348 24162
rect 19292 23940 19348 24110
rect 19740 24444 20020 24500
rect 20076 25284 20132 25294
rect 19516 24052 19572 24062
rect 19516 23958 19572 23996
rect 19292 23874 19348 23884
rect 19740 23938 19796 24444
rect 19852 24276 19908 24286
rect 19852 24050 19908 24220
rect 19852 23998 19854 24050
rect 19906 23998 19908 24050
rect 19852 23986 19908 23998
rect 19740 23886 19742 23938
rect 19794 23886 19796 23938
rect 19740 23874 19796 23886
rect 18340 23436 18564 23492
rect 18284 23426 18340 23436
rect 18060 23326 18062 23378
rect 18114 23326 18116 23378
rect 18060 23268 18116 23326
rect 18060 23202 18116 23212
rect 18508 23378 18564 23436
rect 19180 23426 19236 23436
rect 19964 23714 20020 23726
rect 19964 23662 19966 23714
rect 20018 23662 20020 23714
rect 18508 23326 18510 23378
rect 18562 23326 18564 23378
rect 18284 23044 18340 23054
rect 16828 22146 17332 22148
rect 16828 22094 17166 22146
rect 17218 22094 17332 22146
rect 16828 22092 17332 22094
rect 17836 22932 17892 22942
rect 16828 21698 16884 22092
rect 17164 22082 17220 22092
rect 16828 21646 16830 21698
rect 16882 21646 16884 21698
rect 16716 21588 16772 21598
rect 16716 21494 16772 21532
rect 16380 20974 16382 21026
rect 16434 20974 16436 21026
rect 16380 20962 16436 20974
rect 16156 19506 16212 19516
rect 16604 20802 16660 20814
rect 16604 20750 16606 20802
rect 16658 20750 16660 20802
rect 16604 19236 16660 20750
rect 16828 19236 16884 21646
rect 17052 21586 17108 21598
rect 17052 21534 17054 21586
rect 17106 21534 17108 21586
rect 17052 21364 17108 21534
rect 17724 21364 17780 21374
rect 17052 21362 17780 21364
rect 17052 21310 17726 21362
rect 17778 21310 17780 21362
rect 17052 21308 17780 21310
rect 17724 20914 17780 21308
rect 17724 20862 17726 20914
rect 17778 20862 17780 20914
rect 17724 20850 17780 20862
rect 17724 20580 17780 20590
rect 17500 20020 17556 20030
rect 17052 19908 17108 19918
rect 17052 19906 17220 19908
rect 17052 19854 17054 19906
rect 17106 19854 17220 19906
rect 17052 19852 17220 19854
rect 17052 19842 17108 19852
rect 16940 19348 16996 19358
rect 16940 19254 16996 19292
rect 16268 19012 16324 19022
rect 16492 19012 16548 19022
rect 16268 19010 16436 19012
rect 16268 18958 16270 19010
rect 16322 18958 16436 19010
rect 16268 18956 16436 18958
rect 16268 18946 16324 18956
rect 16268 18788 16324 18798
rect 16156 18338 16212 18350
rect 16156 18286 16158 18338
rect 16210 18286 16212 18338
rect 16156 17108 16212 18286
rect 16268 17890 16324 18732
rect 16380 18676 16436 18956
rect 16380 18610 16436 18620
rect 16268 17838 16270 17890
rect 16322 17838 16324 17890
rect 16268 17826 16324 17838
rect 16380 18452 16436 18462
rect 16156 17052 16324 17108
rect 16156 16884 16212 16894
rect 16156 16790 16212 16828
rect 16268 16324 16324 17052
rect 16380 16884 16436 18396
rect 16380 16818 16436 16828
rect 16268 16210 16324 16268
rect 16268 16158 16270 16210
rect 16322 16158 16324 16210
rect 16268 16146 16324 16158
rect 16492 16212 16548 18956
rect 16604 18674 16660 19180
rect 16604 18622 16606 18674
rect 16658 18622 16660 18674
rect 16604 18610 16660 18622
rect 16716 19180 16884 19236
rect 17052 19236 17108 19246
rect 16716 18452 16772 19180
rect 17052 19142 17108 19180
rect 16828 19012 16884 19022
rect 16828 19010 17108 19012
rect 16828 18958 16830 19010
rect 16882 18958 17108 19010
rect 16828 18956 17108 18958
rect 16828 18946 16884 18956
rect 16940 18788 16996 18798
rect 16716 18386 16772 18396
rect 16828 18676 16884 18686
rect 16828 17444 16884 18620
rect 16940 18562 16996 18732
rect 16940 18510 16942 18562
rect 16994 18510 16996 18562
rect 16940 18116 16996 18510
rect 17052 18452 17108 18956
rect 17164 18788 17220 19852
rect 17276 19348 17332 19358
rect 17276 19254 17332 19292
rect 17164 18722 17220 18732
rect 17500 19234 17556 19964
rect 17500 19182 17502 19234
rect 17554 19182 17556 19234
rect 17052 18386 17108 18396
rect 16940 18050 16996 18060
rect 16604 17388 16884 17444
rect 16940 17666 16996 17678
rect 16940 17614 16942 17666
rect 16994 17614 16996 17666
rect 16604 16212 16660 17388
rect 16828 16994 16884 17006
rect 16828 16942 16830 16994
rect 16882 16942 16884 16994
rect 16716 16882 16772 16894
rect 16716 16830 16718 16882
rect 16770 16830 16772 16882
rect 16716 16772 16772 16830
rect 16828 16884 16884 16942
rect 16940 16996 16996 17614
rect 17052 17108 17108 17118
rect 17052 17014 17108 17052
rect 16940 16930 16996 16940
rect 17500 16884 17556 19182
rect 17724 18562 17780 20524
rect 17836 20130 17892 22876
rect 18284 21810 18340 22988
rect 18508 22932 18564 23326
rect 19068 23268 19124 23278
rect 19068 23174 19124 23212
rect 19180 23266 19236 23278
rect 19180 23214 19182 23266
rect 19234 23214 19236 23266
rect 18508 22866 18564 22876
rect 19180 22932 19236 23214
rect 19964 23268 20020 23662
rect 19964 23202 20020 23212
rect 20076 23266 20132 25228
rect 20300 24722 20356 25564
rect 20412 25394 20468 26908
rect 20524 26852 20580 27694
rect 21084 27746 21140 27758
rect 21084 27694 21086 27746
rect 21138 27694 21140 27746
rect 20748 26964 20804 26974
rect 21084 26908 21140 27694
rect 20748 26870 20804 26908
rect 20524 26786 20580 26796
rect 20860 26852 21140 26908
rect 20532 26684 20796 26694
rect 20588 26628 20636 26684
rect 20692 26628 20740 26684
rect 20532 26618 20796 26628
rect 20636 26404 20692 26414
rect 20524 26348 20636 26404
rect 20524 25844 20580 26348
rect 20636 26272 20692 26348
rect 20748 26292 20804 26302
rect 20860 26292 20916 26852
rect 20748 26290 20916 26292
rect 20748 26238 20750 26290
rect 20802 26238 20916 26290
rect 20748 26236 20916 26238
rect 20748 26226 20804 26236
rect 20524 25778 20580 25788
rect 20636 26066 20692 26078
rect 20636 26014 20638 26066
rect 20690 26014 20692 26066
rect 20636 25620 20692 26014
rect 20636 25554 20692 25564
rect 20412 25342 20414 25394
rect 20466 25342 20468 25394
rect 20412 25330 20468 25342
rect 20524 25394 20580 25406
rect 20524 25342 20526 25394
rect 20578 25342 20580 25394
rect 20524 25284 20580 25342
rect 20524 25218 20580 25228
rect 20860 25284 20916 26236
rect 20532 25116 20796 25126
rect 20588 25060 20636 25116
rect 20692 25060 20740 25116
rect 20532 25050 20796 25060
rect 20300 24670 20302 24722
rect 20354 24670 20356 24722
rect 20300 24658 20356 24670
rect 20860 24050 20916 25228
rect 20860 23998 20862 24050
rect 20914 23998 20916 24050
rect 20860 23986 20916 23998
rect 20532 23548 20796 23558
rect 20076 23214 20078 23266
rect 20130 23214 20132 23266
rect 20076 23202 20132 23214
rect 20188 23492 20244 23502
rect 20588 23492 20636 23548
rect 20692 23492 20740 23548
rect 21196 23492 21252 28252
rect 21756 27860 21812 29148
rect 22876 28756 22932 29260
rect 22764 28754 22932 28756
rect 22764 28702 22878 28754
rect 22930 28702 22932 28754
rect 22764 28700 22932 28702
rect 22428 28420 22484 28430
rect 22428 28418 22596 28420
rect 22428 28366 22430 28418
rect 22482 28366 22596 28418
rect 22428 28364 22596 28366
rect 22428 28354 22484 28364
rect 22428 27970 22484 27982
rect 22428 27918 22430 27970
rect 22482 27918 22484 27970
rect 21868 27860 21924 27870
rect 21756 27804 21868 27860
rect 21868 27766 21924 27804
rect 21420 27748 21476 27758
rect 21420 27746 21588 27748
rect 21420 27694 21422 27746
rect 21474 27694 21588 27746
rect 21420 27692 21588 27694
rect 21420 27682 21476 27692
rect 21420 26964 21476 26974
rect 21420 26180 21476 26908
rect 21532 26852 21588 27692
rect 22428 26964 22484 27918
rect 22540 27860 22596 28364
rect 22652 27860 22708 27870
rect 22540 27858 22708 27860
rect 22540 27806 22654 27858
rect 22706 27806 22708 27858
rect 22540 27804 22708 27806
rect 22652 27076 22708 27804
rect 22764 27746 22820 28700
rect 22876 28690 22932 28700
rect 23212 28532 23268 35868
rect 23324 35700 23380 35710
rect 23324 35606 23380 35644
rect 23660 35700 23716 35710
rect 23548 35140 23604 35150
rect 23548 34914 23604 35084
rect 23548 34862 23550 34914
rect 23602 34862 23604 34914
rect 23548 34850 23604 34862
rect 23660 34802 23716 35644
rect 23884 34914 23940 36316
rect 24892 35922 24948 36540
rect 26684 36594 26740 37884
rect 26684 36542 26686 36594
rect 26738 36542 26740 36594
rect 26684 36530 26740 36542
rect 27804 36596 27860 36606
rect 24892 35870 24894 35922
rect 24946 35870 24948 35922
rect 24892 35858 24948 35870
rect 25228 36484 25284 36494
rect 25228 36258 25284 36428
rect 27804 36482 27860 36540
rect 29372 36594 29428 37884
rect 30192 36876 30456 36886
rect 30248 36820 30296 36876
rect 30352 36820 30400 36876
rect 30192 36810 30456 36820
rect 29372 36542 29374 36594
rect 29426 36542 29428 36594
rect 29372 36530 29428 36542
rect 31276 36594 31332 39200
rect 33740 38164 33796 39200
rect 33740 38108 34132 38164
rect 33964 37940 34020 37950
rect 33964 36708 34020 37884
rect 31276 36542 31278 36594
rect 31330 36542 31332 36594
rect 31276 36530 31332 36542
rect 33516 36596 33572 36606
rect 33516 36502 33572 36540
rect 27804 36430 27806 36482
rect 27858 36430 27860 36482
rect 25788 36372 25844 36382
rect 25788 36278 25844 36316
rect 27356 36372 27412 36382
rect 25228 36206 25230 36258
rect 25282 36206 25284 36258
rect 23996 35700 24052 35710
rect 24556 35700 24612 35710
rect 23996 35698 24612 35700
rect 23996 35646 23998 35698
rect 24050 35646 24558 35698
rect 24610 35646 24612 35698
rect 23996 35644 24612 35646
rect 25228 35700 25284 36206
rect 25900 36258 25956 36270
rect 25900 36206 25902 36258
rect 25954 36206 25956 36258
rect 25228 35644 25508 35700
rect 23996 35634 24052 35644
rect 24556 35634 24612 35644
rect 25340 34916 25396 34926
rect 23884 34862 23886 34914
rect 23938 34862 23940 34914
rect 23884 34850 23940 34862
rect 25116 34860 25340 34916
rect 23660 34750 23662 34802
rect 23714 34750 23716 34802
rect 23660 34738 23716 34750
rect 25004 34692 25060 34702
rect 24892 34636 25004 34692
rect 24780 34468 24836 34478
rect 23324 34130 23380 34142
rect 23324 34078 23326 34130
rect 23378 34078 23380 34130
rect 23324 33684 23380 34078
rect 23884 34132 23940 34142
rect 23884 34038 23940 34076
rect 24332 34018 24388 34030
rect 24332 33966 24334 34018
rect 24386 33966 24388 34018
rect 23324 33458 23380 33628
rect 23436 33908 23492 33918
rect 23436 33572 23492 33852
rect 23884 33908 23940 33918
rect 23548 33572 23604 33582
rect 23436 33570 23604 33572
rect 23436 33518 23550 33570
rect 23602 33518 23604 33570
rect 23436 33516 23604 33518
rect 23548 33506 23604 33516
rect 23884 33570 23940 33852
rect 24332 33684 24388 33966
rect 24332 33618 24388 33628
rect 23884 33518 23886 33570
rect 23938 33518 23940 33570
rect 23884 33506 23940 33518
rect 23324 33406 23326 33458
rect 23378 33406 23380 33458
rect 23324 33394 23380 33406
rect 24108 32564 24164 32574
rect 23436 32452 23492 32462
rect 23436 31948 23492 32396
rect 23996 32452 24052 32462
rect 23436 31892 23604 31948
rect 23548 31556 23604 31892
rect 23996 31890 24052 32396
rect 23996 31838 23998 31890
rect 24050 31838 24052 31890
rect 23996 31826 24052 31838
rect 23548 31490 23604 31500
rect 23884 30994 23940 31006
rect 23884 30942 23886 30994
rect 23938 30942 23940 30994
rect 23436 30882 23492 30894
rect 23436 30830 23438 30882
rect 23490 30830 23492 30882
rect 23436 29988 23492 30830
rect 23884 30210 23940 30942
rect 23996 30324 24052 30334
rect 24108 30324 24164 32508
rect 24444 32564 24500 32574
rect 24444 32562 24724 32564
rect 24444 32510 24446 32562
rect 24498 32510 24724 32562
rect 24444 32508 24724 32510
rect 24444 32498 24500 32508
rect 24556 31666 24612 31678
rect 24556 31614 24558 31666
rect 24610 31614 24612 31666
rect 24556 31556 24612 31614
rect 24556 31490 24612 31500
rect 24668 31554 24724 32508
rect 24780 31780 24836 34412
rect 24892 34244 24948 34636
rect 25004 34560 25060 34636
rect 24892 34150 24948 34188
rect 24892 32676 24948 32686
rect 25116 32676 25172 34860
rect 25340 34784 25396 34860
rect 25452 34804 25508 35644
rect 25900 35588 25956 36206
rect 26124 36260 26180 36270
rect 26124 36166 26180 36204
rect 26796 35924 26852 35934
rect 26796 35830 26852 35868
rect 25900 35522 25956 35532
rect 26012 35812 26068 35822
rect 26012 35138 26068 35756
rect 26460 35812 26516 35822
rect 26460 35698 26516 35756
rect 26460 35646 26462 35698
rect 26514 35646 26516 35698
rect 26460 35634 26516 35646
rect 27356 35698 27412 36316
rect 27468 35924 27524 35934
rect 27468 35830 27524 35868
rect 27356 35646 27358 35698
rect 27410 35646 27412 35698
rect 27356 35634 27412 35646
rect 27468 35700 27524 35710
rect 26236 35588 26292 35598
rect 26236 35494 26292 35532
rect 26012 35086 26014 35138
rect 26066 35086 26068 35138
rect 26012 35074 26068 35086
rect 27468 35026 27524 35644
rect 27468 34974 27470 35026
rect 27522 34974 27524 35026
rect 27468 34962 27524 34974
rect 27804 35028 27860 36430
rect 30492 36482 30548 36494
rect 30492 36430 30494 36482
rect 30546 36430 30548 36482
rect 28588 36372 28644 36382
rect 28588 36278 28644 36316
rect 30492 36372 30548 36430
rect 32396 36484 32452 36494
rect 32396 36482 32676 36484
rect 32396 36430 32398 36482
rect 32450 36430 32676 36482
rect 32396 36428 32676 36430
rect 32396 36418 32452 36428
rect 30492 36306 30548 36316
rect 29596 36260 29652 36270
rect 28476 35924 28532 35962
rect 28476 35858 28532 35868
rect 28588 35812 28644 35822
rect 28588 35718 28644 35756
rect 28476 35700 28532 35710
rect 29372 35700 29428 35710
rect 28476 35606 28532 35644
rect 28812 35698 29428 35700
rect 28812 35646 29374 35698
rect 29426 35646 29428 35698
rect 28812 35644 29428 35646
rect 27916 35028 27972 35038
rect 27804 35026 27972 35028
rect 27804 34974 27918 35026
rect 27970 34974 27972 35026
rect 27804 34972 27972 34974
rect 27916 34962 27972 34972
rect 26572 34916 26628 34926
rect 25452 34738 25508 34748
rect 26236 34914 26628 34916
rect 26236 34862 26574 34914
rect 26626 34862 26628 34914
rect 26236 34860 26628 34862
rect 25676 34692 25732 34702
rect 25676 34598 25732 34636
rect 25900 34690 25956 34702
rect 25900 34638 25902 34690
rect 25954 34638 25956 34690
rect 25900 34132 25956 34638
rect 26012 34692 26068 34702
rect 26012 34242 26068 34636
rect 26236 34354 26292 34860
rect 26572 34850 26628 34860
rect 26796 34916 26852 34926
rect 26796 34822 26852 34860
rect 27132 34916 27188 34926
rect 26236 34302 26238 34354
rect 26290 34302 26292 34354
rect 26236 34290 26292 34302
rect 26012 34190 26014 34242
rect 26066 34190 26068 34242
rect 26012 34178 26068 34190
rect 26460 34244 26516 34254
rect 25900 34066 25956 34076
rect 26236 34132 26292 34142
rect 26236 34038 26292 34076
rect 26460 34130 26516 34188
rect 27132 34242 27188 34860
rect 28364 34916 28420 34926
rect 27468 34356 27524 34366
rect 27468 34262 27524 34300
rect 27132 34190 27134 34242
rect 27186 34190 27188 34242
rect 27132 34178 27188 34190
rect 27244 34244 27300 34254
rect 27244 34150 27300 34188
rect 26460 34078 26462 34130
rect 26514 34078 26516 34130
rect 26460 33908 26516 34078
rect 26460 33842 26516 33852
rect 28364 33458 28420 34860
rect 28812 34914 28868 35644
rect 29372 35634 29428 35644
rect 29596 35698 29652 36204
rect 31164 35924 31220 35934
rect 32060 35924 32116 35934
rect 31164 35922 31556 35924
rect 31164 35870 31166 35922
rect 31218 35870 31556 35922
rect 31164 35868 31556 35870
rect 31164 35858 31220 35868
rect 29596 35646 29598 35698
rect 29650 35646 29652 35698
rect 29596 35634 29652 35646
rect 29820 35700 29876 35710
rect 29820 35606 29876 35644
rect 31052 35698 31108 35710
rect 31052 35646 31054 35698
rect 31106 35646 31108 35698
rect 30192 35308 30456 35318
rect 30248 35252 30296 35308
rect 30352 35252 30400 35308
rect 30192 35242 30456 35252
rect 28812 34862 28814 34914
rect 28866 34862 28868 34914
rect 28812 34850 28868 34862
rect 30268 35140 30324 35150
rect 28476 34804 28532 34814
rect 28476 34710 28532 34748
rect 29596 34690 29652 34702
rect 29596 34638 29598 34690
rect 29650 34638 29652 34690
rect 29596 34468 29652 34638
rect 29596 34402 29652 34412
rect 30268 34690 30324 35084
rect 31052 35140 31108 35646
rect 31052 35074 31108 35084
rect 31388 35698 31444 35710
rect 31388 35646 31390 35698
rect 31442 35646 31444 35698
rect 31388 35026 31444 35646
rect 31388 34974 31390 35026
rect 31442 34974 31444 35026
rect 31388 34962 31444 34974
rect 31276 34914 31332 34926
rect 31276 34862 31278 34914
rect 31330 34862 31332 34914
rect 30492 34804 30548 34814
rect 31276 34804 31332 34862
rect 30492 34802 31332 34804
rect 30492 34750 30494 34802
rect 30546 34750 31332 34802
rect 30492 34748 31332 34750
rect 30492 34738 30548 34748
rect 30268 34638 30270 34690
rect 30322 34638 30324 34690
rect 30268 34356 30324 34638
rect 30380 34692 30436 34702
rect 30380 34598 30436 34636
rect 30268 34290 30324 34300
rect 28364 33406 28366 33458
rect 28418 33406 28420 33458
rect 28364 33394 28420 33406
rect 28700 34020 28756 34030
rect 28252 33348 28308 33358
rect 24892 32674 25172 32676
rect 24892 32622 24894 32674
rect 24946 32622 25172 32674
rect 24892 32620 25172 32622
rect 27020 33124 27076 33134
rect 24892 32610 24948 32620
rect 26908 31890 26964 31902
rect 26908 31838 26910 31890
rect 26962 31838 26964 31890
rect 24892 31780 24948 31790
rect 24780 31778 24948 31780
rect 24780 31726 24894 31778
rect 24946 31726 24948 31778
rect 24780 31724 24948 31726
rect 24892 31714 24948 31724
rect 24668 31502 24670 31554
rect 24722 31502 24724 31554
rect 23996 30322 24164 30324
rect 23996 30270 23998 30322
rect 24050 30270 24164 30322
rect 23996 30268 24164 30270
rect 24220 31220 24276 31230
rect 23996 30258 24052 30268
rect 23884 30158 23886 30210
rect 23938 30158 23940 30210
rect 23436 29922 23492 29932
rect 23548 30098 23604 30110
rect 23548 30046 23550 30098
rect 23602 30046 23604 30098
rect 23548 29092 23604 30046
rect 23660 29428 23716 29438
rect 23660 29334 23716 29372
rect 23548 29026 23604 29036
rect 23884 28644 23940 30158
rect 24108 30098 24164 30110
rect 24108 30046 24110 30098
rect 24162 30046 24164 30098
rect 24108 29988 24164 30046
rect 24108 29922 24164 29932
rect 23996 29538 24052 29550
rect 23996 29486 23998 29538
rect 24050 29486 24052 29538
rect 23996 29428 24052 29486
rect 23996 29362 24052 29372
rect 24220 29428 24276 31164
rect 24332 31108 24388 31118
rect 24668 31108 24724 31502
rect 24332 31106 24724 31108
rect 24332 31054 24334 31106
rect 24386 31054 24724 31106
rect 24332 31052 24724 31054
rect 25340 31554 25396 31566
rect 25340 31502 25342 31554
rect 25394 31502 25396 31554
rect 24332 31042 24388 31052
rect 24892 30882 24948 30894
rect 24892 30830 24894 30882
rect 24946 30830 24948 30882
rect 24892 30772 24948 30830
rect 24892 30716 25284 30772
rect 25004 30324 25060 30334
rect 24892 29988 24948 29998
rect 25004 29988 25060 30268
rect 24892 29986 25060 29988
rect 24892 29934 24894 29986
rect 24946 29934 25060 29986
rect 24892 29932 25060 29934
rect 24892 29922 24948 29932
rect 24220 29362 24276 29372
rect 24556 29316 24612 29326
rect 24444 29260 24556 29316
rect 23996 28644 24052 28654
rect 23884 28642 24052 28644
rect 23884 28590 23998 28642
rect 24050 28590 24052 28642
rect 23884 28588 24052 28590
rect 23996 28578 24052 28588
rect 24444 28642 24500 29260
rect 24556 29184 24612 29260
rect 24780 28756 24836 28766
rect 24780 28662 24836 28700
rect 24444 28590 24446 28642
rect 24498 28590 24500 28642
rect 23212 28466 23268 28476
rect 23772 28532 23828 28542
rect 22988 28418 23044 28430
rect 22988 28366 22990 28418
rect 23042 28366 23044 28418
rect 22988 28084 23044 28366
rect 22988 28018 23044 28028
rect 23436 28418 23492 28430
rect 23436 28366 23438 28418
rect 23490 28366 23492 28418
rect 22876 27860 22932 27870
rect 23436 27860 23492 28366
rect 23660 28084 23716 28094
rect 23660 27990 23716 28028
rect 22876 27766 22932 27804
rect 22988 27804 23492 27860
rect 22764 27694 22766 27746
rect 22818 27694 22820 27746
rect 22764 27682 22820 27694
rect 22652 27010 22708 27020
rect 22764 27524 22820 27534
rect 22540 26964 22596 26974
rect 22428 26962 22596 26964
rect 22428 26910 22542 26962
rect 22594 26910 22596 26962
rect 22428 26908 22596 26910
rect 21980 26852 22036 26862
rect 21532 26404 21588 26796
rect 21532 26338 21588 26348
rect 21868 26850 22036 26852
rect 21868 26798 21982 26850
rect 22034 26798 22036 26850
rect 21868 26796 22036 26798
rect 21868 26404 21924 26796
rect 21980 26786 22036 26796
rect 22540 26852 22596 26908
rect 22764 26964 22820 27468
rect 22764 26870 22820 26908
rect 22540 26786 22596 26796
rect 22988 26852 23044 27804
rect 23436 27636 23492 27646
rect 23100 27634 23492 27636
rect 23100 27582 23438 27634
rect 23490 27582 23492 27634
rect 23100 27580 23492 27582
rect 23100 27186 23156 27580
rect 23436 27570 23492 27580
rect 23772 27634 23828 28476
rect 24444 28196 24500 28590
rect 24444 28130 24500 28140
rect 24892 28420 24948 28430
rect 24892 28084 24948 28364
rect 24556 28082 24948 28084
rect 24556 28030 24894 28082
rect 24946 28030 24948 28082
rect 24556 28028 24948 28030
rect 24220 27748 24276 27758
rect 24556 27748 24612 28028
rect 24892 28018 24948 28028
rect 24220 27746 24612 27748
rect 24220 27694 24222 27746
rect 24274 27694 24612 27746
rect 24220 27692 24612 27694
rect 24220 27682 24276 27692
rect 23772 27582 23774 27634
rect 23826 27582 23828 27634
rect 23772 27412 23828 27582
rect 23772 27346 23828 27356
rect 23100 27134 23102 27186
rect 23154 27134 23156 27186
rect 23100 27122 23156 27134
rect 23884 27188 23940 27198
rect 23212 27076 23268 27086
rect 23212 26982 23268 27020
rect 23884 27074 23940 27132
rect 23884 27022 23886 27074
rect 23938 27022 23940 27074
rect 23548 26964 23604 26974
rect 22988 26850 23156 26852
rect 22988 26798 22990 26850
rect 23042 26798 23156 26850
rect 22988 26796 23156 26798
rect 22988 26786 23044 26796
rect 22988 26516 23044 26526
rect 22988 26422 23044 26460
rect 21532 26180 21588 26190
rect 21420 26178 21588 26180
rect 21420 26126 21534 26178
rect 21586 26126 21588 26178
rect 21420 26124 21588 26126
rect 21532 26066 21588 26124
rect 21532 26014 21534 26066
rect 21586 26014 21588 26066
rect 21532 26002 21588 26014
rect 21756 25844 21812 25854
rect 21756 25282 21812 25788
rect 21868 25396 21924 26348
rect 21980 26178 22036 26190
rect 21980 26126 21982 26178
rect 22034 26126 22036 26178
rect 21980 26066 22036 26126
rect 21980 26014 21982 26066
rect 22034 26014 22036 26066
rect 21980 25956 22036 26014
rect 22428 26180 22484 26190
rect 21980 25900 22260 25956
rect 21980 25508 22036 25518
rect 21980 25414 22036 25452
rect 21868 25302 21924 25340
rect 21756 25230 21758 25282
rect 21810 25230 21812 25282
rect 21532 24610 21588 24622
rect 21532 24558 21534 24610
rect 21586 24558 21588 24610
rect 21532 24498 21588 24558
rect 21532 24446 21534 24498
rect 21586 24446 21588 24498
rect 21532 24434 21588 24446
rect 21756 24498 21812 25230
rect 22092 25284 22148 25294
rect 22092 25190 22148 25228
rect 22204 25060 22260 25900
rect 22316 25394 22372 25406
rect 22316 25342 22318 25394
rect 22370 25342 22372 25394
rect 22316 25060 22372 25342
rect 22428 25284 22484 26124
rect 22428 25218 22484 25228
rect 22652 25284 22708 25294
rect 22876 25284 22932 25294
rect 21980 25004 22316 25060
rect 21756 24446 21758 24498
rect 21810 24446 21812 24498
rect 21756 24434 21812 24446
rect 21868 24948 21924 24958
rect 21868 24050 21924 24892
rect 21868 23998 21870 24050
rect 21922 23998 21924 24050
rect 21868 23940 21924 23998
rect 21868 23874 21924 23884
rect 21980 24610 22036 25004
rect 22316 24928 22372 25004
rect 22652 24946 22708 25228
rect 22652 24894 22654 24946
rect 22706 24894 22708 24946
rect 22652 24882 22708 24894
rect 22764 25282 22932 25284
rect 22764 25230 22878 25282
rect 22930 25230 22932 25282
rect 22764 25228 22932 25230
rect 21980 24558 21982 24610
rect 22034 24558 22036 24610
rect 21868 23716 21924 23726
rect 21868 23604 21924 23660
rect 20532 23482 20796 23492
rect 19404 23156 19460 23166
rect 19404 23062 19460 23100
rect 19180 22866 19236 22876
rect 20188 22370 20244 23436
rect 21084 23436 21252 23492
rect 21756 23548 21924 23604
rect 20188 22318 20190 22370
rect 20242 22318 20244 22370
rect 20076 22260 20132 22270
rect 20076 22166 20132 22204
rect 19964 22148 20020 22158
rect 18284 21758 18286 21810
rect 18338 21758 18340 21810
rect 18284 21746 18340 21758
rect 19852 22146 20020 22148
rect 19852 22094 19966 22146
rect 20018 22094 20020 22146
rect 19852 22092 20020 22094
rect 18172 21700 18228 21710
rect 18172 21606 18228 21644
rect 18060 21586 18116 21598
rect 18060 21534 18062 21586
rect 18114 21534 18116 21586
rect 17948 20804 18004 20814
rect 17948 20710 18004 20748
rect 17836 20078 17838 20130
rect 17890 20078 17892 20130
rect 17836 20066 17892 20078
rect 18060 19348 18116 21534
rect 18396 21586 18452 21598
rect 18396 21534 18398 21586
rect 18450 21534 18452 21586
rect 18284 20356 18340 20366
rect 18172 19348 18228 19358
rect 18060 19346 18228 19348
rect 18060 19294 18174 19346
rect 18226 19294 18228 19346
rect 18060 19292 18228 19294
rect 18172 19282 18228 19292
rect 18284 19234 18340 20300
rect 18396 20244 18452 21534
rect 19516 21588 19572 21598
rect 19516 21494 19572 21532
rect 19852 20804 19908 22092
rect 19964 22082 20020 22092
rect 19964 21476 20020 21486
rect 19964 20916 20020 21420
rect 20188 21364 20244 22318
rect 20188 21298 20244 21308
rect 20300 23154 20356 23166
rect 20300 23102 20302 23154
rect 20354 23102 20356 23154
rect 20300 21700 20356 23102
rect 20636 23156 20692 23166
rect 20636 22594 20692 23100
rect 20636 22542 20638 22594
rect 20690 22542 20692 22594
rect 20636 22530 20692 22542
rect 19964 20850 20020 20860
rect 18396 20178 18452 20188
rect 18620 20692 18676 20702
rect 18284 19182 18286 19234
rect 18338 19182 18340 19234
rect 18284 19170 18340 19182
rect 18396 20018 18452 20030
rect 18396 19966 18398 20018
rect 18450 19966 18452 20018
rect 18172 19124 18228 19134
rect 18172 19030 18228 19068
rect 18060 18676 18116 18686
rect 18396 18676 18452 19966
rect 18620 19124 18676 20636
rect 19628 20692 19684 20702
rect 19628 20598 19684 20636
rect 18732 20580 18788 20590
rect 19180 20580 19236 20590
rect 18732 20486 18788 20524
rect 19068 20578 19236 20580
rect 19068 20526 19182 20578
rect 19234 20526 19236 20578
rect 19068 20524 19236 20526
rect 18844 19460 18900 19470
rect 18508 19010 18564 19022
rect 18508 18958 18510 19010
rect 18562 18958 18564 19010
rect 18508 18900 18564 18958
rect 18508 18834 18564 18844
rect 18620 18788 18676 19068
rect 18732 19124 18788 19134
rect 18844 19124 18900 19404
rect 19068 19460 19124 20524
rect 19180 20514 19236 20524
rect 19404 20244 19460 20254
rect 19180 20020 19236 20030
rect 19180 19926 19236 19964
rect 19068 19394 19124 19404
rect 18732 19122 18900 19124
rect 18732 19070 18734 19122
rect 18786 19070 18900 19122
rect 18732 19068 18900 19070
rect 18732 19058 18788 19068
rect 18732 18788 18788 18798
rect 18620 18732 18732 18788
rect 18732 18722 18788 18732
rect 18396 18620 18564 18676
rect 18060 18582 18116 18620
rect 17724 18510 17726 18562
rect 17778 18510 17780 18562
rect 16828 16772 16884 16828
rect 17052 16828 17556 16884
rect 17612 17666 17668 17678
rect 17612 17614 17614 17666
rect 17666 17614 17668 17666
rect 17612 17108 17668 17614
rect 17724 17668 17780 18510
rect 17836 18564 17892 18574
rect 17836 18470 17892 18508
rect 18396 18452 18452 18462
rect 17724 17602 17780 17612
rect 18172 17892 18228 17902
rect 17612 16884 17668 17052
rect 18172 17106 18228 17836
rect 18284 17668 18340 17678
rect 18396 17668 18452 18396
rect 18508 17892 18564 18620
rect 18620 18564 18676 18574
rect 18620 18470 18676 18508
rect 18508 17826 18564 17836
rect 18732 18450 18788 18462
rect 18732 18398 18734 18450
rect 18786 18398 18788 18450
rect 18284 17666 18452 17668
rect 18284 17614 18286 17666
rect 18338 17614 18452 17666
rect 18284 17612 18452 17614
rect 18732 17780 18788 18398
rect 18284 17602 18340 17612
rect 18172 17054 18174 17106
rect 18226 17054 18228 17106
rect 18172 17042 18228 17054
rect 17724 16884 17780 16894
rect 17612 16882 17780 16884
rect 17612 16830 17726 16882
rect 17778 16830 17780 16882
rect 17612 16828 17780 16830
rect 16828 16716 16996 16772
rect 16716 16706 16772 16716
rect 16716 16212 16772 16222
rect 16604 16210 16772 16212
rect 16604 16158 16718 16210
rect 16770 16158 16772 16210
rect 16604 16156 16772 16158
rect 16492 16146 16548 16156
rect 16716 15988 16772 16156
rect 16716 15922 16772 15932
rect 16716 15540 16772 15550
rect 16716 15426 16772 15484
rect 16716 15374 16718 15426
rect 16770 15374 16772 15426
rect 16716 15362 16772 15374
rect 16828 15426 16884 15438
rect 16828 15374 16830 15426
rect 16882 15374 16884 15426
rect 16268 15204 16324 15242
rect 16268 15138 16324 15148
rect 16044 15026 16100 15036
rect 15316 13804 15428 13860
rect 15260 13794 15316 13804
rect 14140 13746 14196 13758
rect 14140 13694 14142 13746
rect 14194 13694 14196 13746
rect 14140 13524 14196 13694
rect 15260 13634 15316 13646
rect 15260 13582 15262 13634
rect 15314 13582 15316 13634
rect 15260 13524 15316 13582
rect 13804 12850 14084 12852
rect 13804 12798 13806 12850
rect 13858 12798 14084 12850
rect 13804 12796 14084 12798
rect 13804 12786 13860 12796
rect 12908 10882 12964 10892
rect 13020 10892 13188 10948
rect 13356 11788 13636 11844
rect 13804 12180 13860 12190
rect 12796 10836 12852 10846
rect 12796 10742 12852 10780
rect 12460 10630 12516 10668
rect 12572 10722 12628 10734
rect 12572 10670 12574 10722
rect 12626 10670 12628 10722
rect 12012 10434 12068 10444
rect 12572 10500 12628 10670
rect 12572 10434 12628 10444
rect 12684 10724 12740 10734
rect 11676 9996 11844 10052
rect 11676 9828 11732 9838
rect 11676 9734 11732 9772
rect 11788 8820 11844 9996
rect 12572 9940 12628 9950
rect 12572 9846 12628 9884
rect 12012 9156 12068 9166
rect 12012 9062 12068 9100
rect 11900 9044 11956 9054
rect 11900 8950 11956 8988
rect 12012 8820 12068 8830
rect 11788 8818 12068 8820
rect 11788 8766 12014 8818
rect 12066 8766 12068 8818
rect 11788 8764 12068 8766
rect 12012 8754 12068 8764
rect 12684 7700 12740 10668
rect 12908 10500 12964 10510
rect 12908 9602 12964 10444
rect 12908 9550 12910 9602
rect 12962 9550 12964 9602
rect 12908 9380 12964 9550
rect 12908 9314 12964 9324
rect 12796 7700 12852 7710
rect 12684 7698 12852 7700
rect 12684 7646 12798 7698
rect 12850 7646 12852 7698
rect 12684 7644 12852 7646
rect 12572 6692 12628 6702
rect 12684 6692 12740 7644
rect 12796 7634 12852 7644
rect 12628 6636 12740 6692
rect 12908 6804 12964 6814
rect 12908 6690 12964 6748
rect 12908 6638 12910 6690
rect 12962 6638 12964 6690
rect 12572 6560 12628 6636
rect 12908 6626 12964 6638
rect 12012 6468 12068 6478
rect 12012 6374 12068 6412
rect 12684 6468 12740 6478
rect 13020 6468 13076 10892
rect 13244 10836 13300 10846
rect 13244 10276 13300 10780
rect 13244 9042 13300 10220
rect 13356 10834 13412 11788
rect 13692 11620 13748 11630
rect 13804 11620 13860 12124
rect 13692 11618 13860 11620
rect 13692 11566 13694 11618
rect 13746 11566 13860 11618
rect 13692 11564 13860 11566
rect 13692 11554 13748 11564
rect 13916 11394 13972 11406
rect 13916 11342 13918 11394
rect 13970 11342 13972 11394
rect 13356 10782 13358 10834
rect 13410 10782 13412 10834
rect 13356 9940 13412 10782
rect 13580 10836 13636 10846
rect 13916 10836 13972 11342
rect 13580 10834 13972 10836
rect 13580 10782 13582 10834
rect 13634 10782 13972 10834
rect 13580 10780 13972 10782
rect 13580 10770 13636 10780
rect 13468 10610 13524 10622
rect 13468 10558 13470 10610
rect 13522 10558 13524 10610
rect 13468 10500 13524 10558
rect 13468 10434 13524 10444
rect 13692 10610 13748 10622
rect 13692 10558 13694 10610
rect 13746 10558 13748 10610
rect 13692 10164 13748 10558
rect 13916 10612 13972 10622
rect 14028 10612 14084 12796
rect 14140 11394 14196 13468
rect 15036 13468 15316 13524
rect 14364 13076 14420 13086
rect 14364 12982 14420 13020
rect 14812 12738 14868 12750
rect 14812 12686 14814 12738
rect 14866 12686 14868 12738
rect 14812 12516 14868 12686
rect 15036 12516 15092 13468
rect 14812 12460 15092 12516
rect 14476 12292 14532 12302
rect 14140 11342 14142 11394
rect 14194 11342 14196 11394
rect 14140 11330 14196 11342
rect 14252 11396 14308 11406
rect 14252 11302 14308 11340
rect 14364 11170 14420 11182
rect 14364 11118 14366 11170
rect 14418 11118 14420 11170
rect 14364 10836 14420 11118
rect 14364 10770 14420 10780
rect 14364 10612 14420 10622
rect 13916 10610 14420 10612
rect 13916 10558 13918 10610
rect 13970 10558 14366 10610
rect 14418 10558 14420 10610
rect 13916 10556 14420 10558
rect 13916 10546 13972 10556
rect 14364 10500 14420 10556
rect 14364 10434 14420 10444
rect 14140 10388 14196 10398
rect 13692 10098 13748 10108
rect 13916 10386 14196 10388
rect 13916 10334 14142 10386
rect 14194 10334 14196 10386
rect 13916 10332 14196 10334
rect 13412 9884 13748 9940
rect 13356 9808 13412 9884
rect 13692 9826 13748 9884
rect 13692 9774 13694 9826
rect 13746 9774 13748 9826
rect 13692 9762 13748 9774
rect 13804 9604 13860 9614
rect 13804 9510 13860 9548
rect 13916 9380 13972 10332
rect 14140 10322 14196 10332
rect 14252 10276 14308 10286
rect 13692 9324 13972 9380
rect 14028 9602 14084 9614
rect 14028 9550 14030 9602
rect 14082 9550 14084 9602
rect 13244 8990 13246 9042
rect 13298 8990 13300 9042
rect 13244 8978 13300 8990
rect 13580 9156 13636 9166
rect 13468 8818 13524 8830
rect 13468 8766 13470 8818
rect 13522 8766 13524 8818
rect 13468 7700 13524 8766
rect 13468 7634 13524 7644
rect 13580 7698 13636 9100
rect 13580 7646 13582 7698
rect 13634 7646 13636 7698
rect 13580 7634 13636 7646
rect 13692 7698 13748 9324
rect 13692 7646 13694 7698
rect 13746 7646 13748 7698
rect 13692 7634 13748 7646
rect 13804 8818 13860 8830
rect 13804 8766 13806 8818
rect 13858 8766 13860 8818
rect 13468 7474 13524 7486
rect 13468 7422 13470 7474
rect 13522 7422 13524 7474
rect 12684 6374 12740 6412
rect 12908 6412 13076 6468
rect 13132 6804 13188 6814
rect 12796 6018 12852 6030
rect 12796 5966 12798 6018
rect 12850 5966 12852 6018
rect 11452 4498 11508 4508
rect 11564 5794 11620 5806
rect 11564 5742 11566 5794
rect 11618 5742 11620 5794
rect 11228 4340 11284 4350
rect 10556 3602 10612 3612
rect 10668 4172 10836 4228
rect 11116 4228 11172 4238
rect 10332 3378 10388 3388
rect 9772 2594 9828 2604
rect 10668 2436 10724 4172
rect 11116 4134 11172 4172
rect 10872 3948 11136 3958
rect 10928 3892 10976 3948
rect 11032 3892 11080 3948
rect 10872 3882 11136 3892
rect 10668 2370 10724 2380
rect 9548 1026 9604 1036
rect 11228 800 11284 4284
rect 11452 4338 11508 4350
rect 11452 4286 11454 4338
rect 11506 4286 11508 4338
rect 11452 4116 11508 4286
rect 11452 4050 11508 4060
rect 11564 3780 11620 5742
rect 12012 5796 12068 5806
rect 12012 5794 12180 5796
rect 12012 5742 12014 5794
rect 12066 5742 12180 5794
rect 12012 5740 12180 5742
rect 12012 5730 12068 5740
rect 12124 5460 12180 5740
rect 12124 5122 12180 5404
rect 12796 5236 12852 5966
rect 12796 5170 12852 5180
rect 12124 5070 12126 5122
rect 12178 5070 12180 5122
rect 11564 3714 11620 3724
rect 11788 4898 11844 4910
rect 11788 4846 11790 4898
rect 11842 4846 11844 4898
rect 11452 3668 11508 3678
rect 11452 3554 11508 3612
rect 11452 3502 11454 3554
rect 11506 3502 11508 3554
rect 11452 3490 11508 3502
rect 11676 3556 11732 3566
rect 11676 3462 11732 3500
rect 11564 3442 11620 3454
rect 11564 3390 11566 3442
rect 11618 3390 11620 3442
rect 11564 3332 11620 3390
rect 11788 3444 11844 4846
rect 12012 4898 12068 4910
rect 12012 4846 12014 4898
rect 12066 4846 12068 4898
rect 12012 4116 12068 4846
rect 12124 4228 12180 5070
rect 12796 4452 12852 4462
rect 12908 4452 12964 6412
rect 13132 5906 13188 6748
rect 13132 5854 13134 5906
rect 13186 5854 13188 5906
rect 13132 5842 13188 5854
rect 13020 5572 13076 5582
rect 13020 5234 13076 5516
rect 13020 5182 13022 5234
rect 13074 5182 13076 5234
rect 13020 5170 13076 5182
rect 13468 5236 13524 7422
rect 13804 7474 13860 8766
rect 13916 8372 13972 8382
rect 14028 8372 14084 9550
rect 13916 8370 14196 8372
rect 13916 8318 13918 8370
rect 13970 8318 14196 8370
rect 13916 8316 14196 8318
rect 13916 8306 13972 8316
rect 13804 7422 13806 7474
rect 13858 7422 13860 7474
rect 13804 7410 13860 7422
rect 14140 7474 14196 8316
rect 14252 8146 14308 10220
rect 14476 9604 14532 12236
rect 14812 12178 14868 12190
rect 14812 12126 14814 12178
rect 14866 12126 14868 12178
rect 14812 11172 14868 12126
rect 14924 11172 14980 11182
rect 14812 11170 14980 11172
rect 14812 11118 14926 11170
rect 14978 11118 14980 11170
rect 14812 11116 14980 11118
rect 15036 11172 15092 12460
rect 15260 13076 15316 13086
rect 15372 13076 15428 13804
rect 15708 13794 15764 13804
rect 16156 14306 16212 14318
rect 16156 14254 16158 14306
rect 16210 14254 16212 14306
rect 16156 13972 16212 14254
rect 15708 13636 15764 13646
rect 15708 13542 15764 13580
rect 16156 13634 16212 13916
rect 16156 13582 16158 13634
rect 16210 13582 16212 13634
rect 15260 13074 15428 13076
rect 15260 13022 15262 13074
rect 15314 13022 15428 13074
rect 15260 13020 15428 13022
rect 15260 11620 15316 13020
rect 15932 12964 15988 12974
rect 15372 12066 15428 12078
rect 15372 12014 15374 12066
rect 15426 12014 15428 12066
rect 15372 11844 15428 12014
rect 15372 11778 15428 11788
rect 15260 11564 15428 11620
rect 15260 11396 15316 11406
rect 15260 11302 15316 11340
rect 15148 11172 15204 11182
rect 15036 11116 15148 11172
rect 14700 10388 14756 10398
rect 14812 10388 14868 11116
rect 14924 11106 14980 11116
rect 14924 10836 14980 10846
rect 14924 10742 14980 10780
rect 15148 10500 15204 11116
rect 15148 10434 15204 10444
rect 14700 10386 14868 10388
rect 14700 10334 14702 10386
rect 14754 10334 14868 10386
rect 14700 10332 14868 10334
rect 14924 10388 14980 10398
rect 14700 10322 14756 10332
rect 14700 10164 14756 10174
rect 14476 9538 14532 9548
rect 14588 9602 14644 9614
rect 14588 9550 14590 9602
rect 14642 9550 14644 9602
rect 14588 9492 14644 9550
rect 14588 9426 14644 9436
rect 14252 8094 14254 8146
rect 14306 8094 14308 8146
rect 14252 8082 14308 8094
rect 14476 9380 14532 9390
rect 14140 7422 14142 7474
rect 14194 7422 14196 7474
rect 14140 7410 14196 7422
rect 14252 7700 14308 7710
rect 13692 6804 13748 6814
rect 13692 6710 13748 6748
rect 13916 6692 13972 6702
rect 13804 6690 13972 6692
rect 13804 6638 13918 6690
rect 13970 6638 13972 6690
rect 13804 6636 13972 6638
rect 13692 5348 13748 5358
rect 13804 5348 13860 6636
rect 13916 6626 13972 6636
rect 14140 6692 14196 6702
rect 14252 6692 14308 7644
rect 14140 6690 14308 6692
rect 14140 6638 14142 6690
rect 14194 6638 14308 6690
rect 14140 6636 14308 6638
rect 14140 6626 14196 6636
rect 14252 6466 14308 6478
rect 14252 6414 14254 6466
rect 14306 6414 14308 6466
rect 14252 6356 14308 6414
rect 14252 6290 14308 6300
rect 14364 6466 14420 6478
rect 14364 6414 14366 6466
rect 14418 6414 14420 6466
rect 14028 5906 14084 5918
rect 14028 5854 14030 5906
rect 14082 5854 14084 5906
rect 13692 5346 13860 5348
rect 13692 5294 13694 5346
rect 13746 5294 13860 5346
rect 13692 5292 13860 5294
rect 13916 5572 13972 5582
rect 13692 5282 13748 5292
rect 13468 5170 13524 5180
rect 13804 4564 13860 4574
rect 13916 4564 13972 5516
rect 14028 5346 14084 5854
rect 14364 5572 14420 6414
rect 14364 5506 14420 5516
rect 14028 5294 14030 5346
rect 14082 5294 14084 5346
rect 14028 5124 14084 5294
rect 14252 5236 14308 5246
rect 14252 5142 14308 5180
rect 14028 5058 14084 5068
rect 13804 4562 13972 4564
rect 13804 4510 13806 4562
rect 13858 4510 13972 4562
rect 13804 4508 13972 4510
rect 14028 4564 14084 4574
rect 13804 4498 13860 4508
rect 12796 4450 12964 4452
rect 12796 4398 12798 4450
rect 12850 4398 12964 4450
rect 12796 4396 12964 4398
rect 12796 4386 12852 4396
rect 12236 4340 12292 4350
rect 12236 4246 12292 4284
rect 12124 4162 12180 4172
rect 13356 4228 13412 4238
rect 13356 4134 13412 4172
rect 12012 4050 12068 4060
rect 13356 3780 13412 3790
rect 11900 3444 11956 3454
rect 11788 3442 11956 3444
rect 11788 3390 11902 3442
rect 11954 3390 11956 3442
rect 11788 3388 11956 3390
rect 11900 3378 11956 3388
rect 12908 3444 12964 3482
rect 12908 3378 12964 3388
rect 11564 3276 11844 3332
rect 11788 868 11844 3276
rect 11788 802 11844 812
rect 13356 800 13412 3724
rect 13580 3780 13636 3790
rect 13580 3554 13636 3724
rect 14028 3666 14084 4508
rect 14028 3614 14030 3666
rect 14082 3614 14084 3666
rect 14028 3602 14084 3614
rect 13580 3502 13582 3554
rect 13634 3502 13636 3554
rect 13580 3490 13636 3502
rect 14476 980 14532 9324
rect 14700 9266 14756 10108
rect 14700 9214 14702 9266
rect 14754 9214 14756 9266
rect 14700 9202 14756 9214
rect 14588 8260 14644 8270
rect 14588 7700 14644 8204
rect 14588 7606 14644 7644
rect 14812 7700 14868 7710
rect 14924 7700 14980 10332
rect 15372 10164 15428 11564
rect 15484 11396 15540 11406
rect 15484 10610 15540 11340
rect 15484 10558 15486 10610
rect 15538 10558 15540 10610
rect 15484 10388 15540 10558
rect 15484 10322 15540 10332
rect 15596 11284 15652 11294
rect 15372 10098 15428 10108
rect 15036 9940 15092 9950
rect 15596 9940 15652 11228
rect 15708 11172 15764 11182
rect 15708 11078 15764 11116
rect 15932 10836 15988 12908
rect 16156 12740 16212 13582
rect 16492 14306 16548 14318
rect 16492 14254 16494 14306
rect 16546 14254 16548 14306
rect 16156 12738 16324 12740
rect 16156 12686 16158 12738
rect 16210 12686 16324 12738
rect 16156 12684 16324 12686
rect 16156 12674 16212 12684
rect 16156 12404 16212 12414
rect 16156 12310 16212 12348
rect 16156 12180 16212 12190
rect 16156 11506 16212 12124
rect 16268 11956 16324 12684
rect 16492 12180 16548 14254
rect 16828 13972 16884 15374
rect 16828 13878 16884 13916
rect 16716 13746 16772 13758
rect 16716 13694 16718 13746
rect 16770 13694 16772 13746
rect 16716 13636 16772 13694
rect 16716 13188 16772 13580
rect 16716 13122 16772 13132
rect 16940 13076 16996 16716
rect 17052 15538 17108 16828
rect 17724 16818 17780 16828
rect 18284 16884 18340 16894
rect 18284 16790 18340 16828
rect 18396 16882 18452 16894
rect 18396 16830 18398 16882
rect 18450 16830 18452 16882
rect 17948 16770 18004 16782
rect 17948 16718 17950 16770
rect 18002 16718 18004 16770
rect 17164 16212 17220 16222
rect 17164 16118 17220 16156
rect 17388 16212 17444 16222
rect 17052 15486 17054 15538
rect 17106 15486 17108 15538
rect 17052 15474 17108 15486
rect 17388 15316 17444 16156
rect 17948 16210 18004 16718
rect 17948 16158 17950 16210
rect 18002 16158 18004 16210
rect 17948 16146 18004 16158
rect 18172 16324 18228 16334
rect 18172 16098 18228 16268
rect 18396 16212 18452 16830
rect 18172 16046 18174 16098
rect 18226 16046 18228 16098
rect 18172 16034 18228 16046
rect 18284 16156 18452 16212
rect 18508 16772 18564 16782
rect 18508 16212 18564 16716
rect 18732 16324 18788 17724
rect 18732 16258 18788 16268
rect 17948 15988 18004 15998
rect 17052 15260 17444 15316
rect 17836 15876 17892 15886
rect 17836 15316 17892 15820
rect 17052 14642 17108 15260
rect 17836 15250 17892 15260
rect 17052 14590 17054 14642
rect 17106 14590 17108 14642
rect 17052 14578 17108 14590
rect 17612 14642 17668 14654
rect 17612 14590 17614 14642
rect 17666 14590 17668 14642
rect 17052 13972 17108 13982
rect 17612 13972 17668 14590
rect 17052 13970 17668 13972
rect 17052 13918 17054 13970
rect 17106 13918 17668 13970
rect 17052 13916 17668 13918
rect 17052 13906 17108 13916
rect 17612 13522 17668 13916
rect 17836 13748 17892 13758
rect 17836 13654 17892 13692
rect 17612 13470 17614 13522
rect 17666 13470 17668 13522
rect 17612 13458 17668 13470
rect 17724 13636 17780 13646
rect 17164 13076 17220 13086
rect 16940 13074 17220 13076
rect 16940 13022 17166 13074
rect 17218 13022 17220 13074
rect 16940 13020 17220 13022
rect 16716 12740 16772 12750
rect 16492 12086 16548 12124
rect 16604 12738 16772 12740
rect 16604 12686 16718 12738
rect 16770 12686 16772 12738
rect 16604 12684 16772 12686
rect 16604 11956 16660 12684
rect 16716 12674 16772 12684
rect 17052 12404 17108 13020
rect 17164 13010 17220 13020
rect 17724 12516 17780 13580
rect 17836 13076 17892 13086
rect 17948 13076 18004 15932
rect 18284 15652 18340 16156
rect 18396 15988 18452 15998
rect 18508 15988 18564 16156
rect 18396 15986 18564 15988
rect 18396 15934 18398 15986
rect 18450 15934 18564 15986
rect 18396 15932 18564 15934
rect 18396 15922 18452 15932
rect 18172 15596 18340 15652
rect 18060 15540 18116 15550
rect 18060 15314 18116 15484
rect 18060 15262 18062 15314
rect 18114 15262 18116 15314
rect 18060 15204 18116 15262
rect 18060 15138 18116 15148
rect 17836 13074 18004 13076
rect 17836 13022 17838 13074
rect 17890 13022 18004 13074
rect 17836 13020 18004 13022
rect 17836 13010 17892 13020
rect 17724 12450 17780 12460
rect 17948 12852 18004 13020
rect 17052 12272 17108 12348
rect 17612 12068 17668 12078
rect 17612 12066 17780 12068
rect 17612 12014 17614 12066
rect 17666 12014 17780 12066
rect 17612 12012 17780 12014
rect 17612 12002 17668 12012
rect 16268 11900 16660 11956
rect 16156 11454 16158 11506
rect 16210 11454 16212 11506
rect 16156 11396 16212 11454
rect 16156 11330 16212 11340
rect 16604 11060 16660 11900
rect 16716 11284 16772 11294
rect 16716 11190 16772 11228
rect 17724 11284 17780 12012
rect 17724 11190 17780 11228
rect 17276 11172 17332 11182
rect 17164 11116 17276 11172
rect 16604 11004 16772 11060
rect 15932 10704 15988 10780
rect 16604 10498 16660 10510
rect 16604 10446 16606 10498
rect 16658 10446 16660 10498
rect 16604 10388 16660 10446
rect 16604 10322 16660 10332
rect 15036 9268 15092 9884
rect 15148 9938 15652 9940
rect 15148 9886 15598 9938
rect 15650 9886 15652 9938
rect 15148 9884 15652 9886
rect 15148 9492 15204 9884
rect 15596 9874 15652 9884
rect 15148 9426 15204 9436
rect 15260 9604 15316 9614
rect 15148 9268 15204 9278
rect 15036 9266 15204 9268
rect 15036 9214 15150 9266
rect 15202 9214 15204 9266
rect 15036 9212 15204 9214
rect 15148 9202 15204 9212
rect 15260 8932 15316 9548
rect 15932 9604 15988 9614
rect 15484 8932 15540 8942
rect 15148 8930 15540 8932
rect 15148 8878 15486 8930
rect 15538 8878 15540 8930
rect 15148 8876 15540 8878
rect 14812 7698 14924 7700
rect 14812 7646 14814 7698
rect 14866 7646 14924 7698
rect 14812 7644 14924 7646
rect 14980 7644 15092 7700
rect 14812 7634 14868 7644
rect 14924 7634 14980 7644
rect 14924 7474 14980 7486
rect 14924 7422 14926 7474
rect 14978 7422 14980 7474
rect 14924 7364 14980 7422
rect 14924 7298 14980 7308
rect 15036 6802 15092 7644
rect 15036 6750 15038 6802
rect 15090 6750 15092 6802
rect 15036 6738 15092 6750
rect 15148 6580 15204 8876
rect 15484 8866 15540 8876
rect 15260 8260 15316 8270
rect 15260 8166 15316 8204
rect 15820 8036 15876 8046
rect 15820 7942 15876 7980
rect 15372 7700 15428 7710
rect 15372 7606 15428 7644
rect 15820 7700 15876 7710
rect 15932 7700 15988 9548
rect 16268 9604 16324 9614
rect 16268 9510 16324 9548
rect 16716 9602 16772 11004
rect 16716 9550 16718 9602
rect 16770 9550 16772 9602
rect 16716 9492 16772 9550
rect 16716 9426 16772 9436
rect 17052 10610 17108 10622
rect 17052 10558 17054 10610
rect 17106 10558 17108 10610
rect 17052 10052 17108 10558
rect 17052 9044 17108 9996
rect 17052 8978 17108 8988
rect 17164 10276 17220 11116
rect 17276 11040 17332 11116
rect 17836 11172 17892 11182
rect 17836 11078 17892 11116
rect 17948 11172 18004 12796
rect 18060 14532 18116 14542
rect 18172 14532 18228 15596
rect 18508 15538 18564 15932
rect 18508 15486 18510 15538
rect 18562 15486 18564 15538
rect 18508 15474 18564 15486
rect 18844 15540 18900 19068
rect 19292 18564 19348 18574
rect 19180 17892 19236 17902
rect 19180 17798 19236 17836
rect 19068 17780 19124 17790
rect 19068 17666 19124 17724
rect 19068 17614 19070 17666
rect 19122 17614 19124 17666
rect 19068 17602 19124 17614
rect 19180 17442 19236 17454
rect 19180 17390 19182 17442
rect 19234 17390 19236 17442
rect 19180 17332 19236 17390
rect 18956 17276 19236 17332
rect 18956 15988 19012 17276
rect 19180 17108 19236 17118
rect 19292 17108 19348 18508
rect 19180 17106 19292 17108
rect 19180 17054 19182 17106
rect 19234 17054 19292 17106
rect 19180 17052 19292 17054
rect 18956 15922 19012 15932
rect 19068 16996 19124 17006
rect 18844 15474 18900 15484
rect 19068 15540 19124 16940
rect 19180 16210 19236 17052
rect 19292 16976 19348 17052
rect 19404 18450 19460 20188
rect 19516 20132 19572 20142
rect 19516 20018 19572 20076
rect 19516 19966 19518 20018
rect 19570 19966 19572 20018
rect 19516 18676 19572 19966
rect 19628 19348 19684 19358
rect 19628 19254 19684 19292
rect 19740 19236 19796 19246
rect 19740 19142 19796 19180
rect 19628 19012 19684 19022
rect 19628 18918 19684 18956
rect 19516 18610 19572 18620
rect 19740 18788 19796 18798
rect 19404 18398 19406 18450
rect 19458 18398 19460 18450
rect 19404 16772 19460 18398
rect 19740 18004 19796 18732
rect 19852 18674 19908 20748
rect 20300 20692 20356 21644
rect 20412 22370 20468 22382
rect 20412 22318 20414 22370
rect 20466 22318 20468 22370
rect 20412 20916 20468 22318
rect 21084 22372 21140 23436
rect 21084 22306 21140 22316
rect 21196 23268 21252 23278
rect 20532 21980 20796 21990
rect 20588 21924 20636 21980
rect 20692 21924 20740 21980
rect 20532 21914 20796 21924
rect 20636 21812 20692 21822
rect 20636 21810 20916 21812
rect 20636 21758 20638 21810
rect 20690 21758 20916 21810
rect 20636 21756 20916 21758
rect 20636 21746 20692 21756
rect 20748 21586 20804 21598
rect 20748 21534 20750 21586
rect 20802 21534 20804 21586
rect 20748 21476 20804 21534
rect 20748 21410 20804 21420
rect 20636 21364 20692 21374
rect 20636 21270 20692 21308
rect 20860 20916 20916 21756
rect 21196 21810 21252 23212
rect 21644 23268 21700 23278
rect 21308 23156 21364 23166
rect 21308 23062 21364 23100
rect 21644 23154 21700 23212
rect 21644 23102 21646 23154
rect 21698 23102 21700 23154
rect 21644 23090 21700 23102
rect 21756 21812 21812 23548
rect 21196 21758 21198 21810
rect 21250 21758 21252 21810
rect 21196 21746 21252 21758
rect 21644 21756 21812 21812
rect 21868 22146 21924 22158
rect 21868 22094 21870 22146
rect 21922 22094 21924 22146
rect 21420 21700 21476 21710
rect 21420 21606 21476 21644
rect 21532 21588 21588 21598
rect 21532 21494 21588 21532
rect 21644 21476 21700 21756
rect 21868 21700 21924 22094
rect 20412 20850 20468 20860
rect 20748 20860 21028 20916
rect 20524 20692 20580 20702
rect 20300 20690 20580 20692
rect 20300 20638 20526 20690
rect 20578 20638 20580 20690
rect 20300 20636 20580 20638
rect 20524 20626 20580 20636
rect 20748 20690 20804 20860
rect 20748 20638 20750 20690
rect 20802 20638 20804 20690
rect 20748 20626 20804 20638
rect 20860 20692 20916 20702
rect 20860 20598 20916 20636
rect 20076 20578 20132 20590
rect 20076 20526 20078 20578
rect 20130 20526 20132 20578
rect 20076 20244 20132 20526
rect 20532 20412 20796 20422
rect 20588 20356 20636 20412
rect 20692 20356 20740 20412
rect 20532 20346 20796 20356
rect 20076 20178 20132 20188
rect 20860 20244 20916 20254
rect 20860 20150 20916 20188
rect 20972 19460 21028 20860
rect 21644 20802 21700 21420
rect 21644 20750 21646 20802
rect 21698 20750 21700 20802
rect 21644 20468 21700 20750
rect 21644 20402 21700 20412
rect 21756 21644 21868 21700
rect 21756 20692 21812 21644
rect 21868 21634 21924 21644
rect 21868 20916 21924 20926
rect 21868 20822 21924 20860
rect 21868 20692 21924 20702
rect 21756 20690 21924 20692
rect 21756 20638 21870 20690
rect 21922 20638 21924 20690
rect 21756 20636 21924 20638
rect 21756 20244 21812 20636
rect 21868 20626 21924 20636
rect 21756 20178 21812 20188
rect 21532 20132 21588 20142
rect 20972 19394 21028 19404
rect 21308 19906 21364 19918
rect 21308 19854 21310 19906
rect 21362 19854 21364 19906
rect 21308 19460 21364 19854
rect 21308 19394 21364 19404
rect 21532 19236 21588 20076
rect 21532 19142 21588 19180
rect 20188 19124 20244 19134
rect 20188 19030 20244 19068
rect 20860 19124 20916 19134
rect 19852 18622 19854 18674
rect 19906 18622 19908 18674
rect 19852 18610 19908 18622
rect 19964 19010 20020 19022
rect 19964 18958 19966 19010
rect 20018 18958 20020 19010
rect 19740 17778 19796 17948
rect 19740 17726 19742 17778
rect 19794 17726 19796 17778
rect 19740 17714 19796 17726
rect 19964 17780 20020 18958
rect 20412 19012 20468 19022
rect 20188 18676 20244 18686
rect 20076 18564 20132 18574
rect 20076 18470 20132 18508
rect 20188 18562 20244 18620
rect 20188 18510 20190 18562
rect 20242 18510 20244 18562
rect 19628 17332 19684 17342
rect 19628 17106 19684 17276
rect 19628 17054 19630 17106
rect 19682 17054 19684 17106
rect 19628 17042 19684 17054
rect 19404 16706 19460 16716
rect 19852 16996 19908 17006
rect 19180 16158 19182 16210
rect 19234 16158 19236 16210
rect 19180 16146 19236 16158
rect 19292 16660 19348 16670
rect 19180 15540 19236 15550
rect 19068 15538 19236 15540
rect 19068 15486 19182 15538
rect 19234 15486 19236 15538
rect 19068 15484 19236 15486
rect 18284 15314 18340 15326
rect 18284 15262 18286 15314
rect 18338 15262 18340 15314
rect 18284 15204 18340 15262
rect 18732 15316 18788 15326
rect 18732 15222 18788 15260
rect 18284 15138 18340 15148
rect 18396 15202 18452 15214
rect 18396 15150 18398 15202
rect 18450 15150 18452 15202
rect 18396 15148 18452 15150
rect 19068 15148 19124 15484
rect 19180 15474 19236 15484
rect 18396 15092 18676 15148
rect 18060 14530 18228 14532
rect 18060 14478 18062 14530
rect 18114 14478 18228 14530
rect 18060 14476 18228 14478
rect 18060 11394 18116 14476
rect 18396 13748 18452 13758
rect 18172 13746 18452 13748
rect 18172 13694 18398 13746
rect 18450 13694 18452 13746
rect 18172 13692 18452 13694
rect 18172 13522 18228 13692
rect 18396 13682 18452 13692
rect 18620 13746 18676 15092
rect 18844 15092 19124 15148
rect 18844 13970 18900 15092
rect 19180 14530 19236 14542
rect 19180 14478 19182 14530
rect 19234 14478 19236 14530
rect 18844 13918 18846 13970
rect 18898 13918 18900 13970
rect 18844 13906 18900 13918
rect 18956 13972 19012 13982
rect 18956 13878 19012 13916
rect 18620 13694 18622 13746
rect 18674 13694 18676 13746
rect 18620 13682 18676 13694
rect 19068 13748 19124 13758
rect 18172 13470 18174 13522
rect 18226 13470 18228 13522
rect 18172 13458 18228 13470
rect 18172 13076 18228 13086
rect 18172 12290 18228 13020
rect 18844 13076 18900 13086
rect 18396 12964 18452 12974
rect 18396 12870 18452 12908
rect 18508 12852 18564 12862
rect 18508 12758 18564 12796
rect 18732 12852 18788 12862
rect 18732 12758 18788 12796
rect 18284 12404 18340 12414
rect 18284 12310 18340 12348
rect 18172 12238 18174 12290
rect 18226 12238 18228 12290
rect 18172 12180 18228 12238
rect 18172 12114 18228 12124
rect 18732 12180 18788 12190
rect 18284 11956 18340 11966
rect 18284 11954 18452 11956
rect 18284 11902 18286 11954
rect 18338 11902 18452 11954
rect 18284 11900 18452 11902
rect 18284 11890 18340 11900
rect 18396 11508 18452 11900
rect 18620 11508 18676 11518
rect 18396 11452 18620 11508
rect 18060 11342 18062 11394
rect 18114 11342 18116 11394
rect 18620 11376 18676 11452
rect 18060 11330 18116 11342
rect 17948 11116 18228 11172
rect 17948 10948 18004 11116
rect 17612 10892 18004 10948
rect 17612 10834 17668 10892
rect 17612 10782 17614 10834
rect 17666 10782 17668 10834
rect 17612 10770 17668 10782
rect 18172 10724 18228 11116
rect 18620 10836 18676 10846
rect 18732 10836 18788 12124
rect 18620 10834 18788 10836
rect 18620 10782 18622 10834
rect 18674 10782 18788 10834
rect 18620 10780 18788 10782
rect 18620 10770 18676 10780
rect 18172 10592 18228 10668
rect 18396 10612 18452 10622
rect 18284 10610 18452 10612
rect 15820 7698 15932 7700
rect 15820 7646 15822 7698
rect 15874 7646 15932 7698
rect 15820 7644 15932 7646
rect 15820 7364 15876 7644
rect 15932 7568 15988 7644
rect 16156 8484 16212 8494
rect 17164 8484 17220 10220
rect 18284 10558 18398 10610
rect 18450 10558 18452 10610
rect 18284 10556 18452 10558
rect 17388 10050 17444 10062
rect 17388 9998 17390 10050
rect 17442 9998 17444 10050
rect 17388 9940 17444 9998
rect 18172 10052 18228 10062
rect 18284 10052 18340 10556
rect 18396 10546 18452 10556
rect 18732 10610 18788 10622
rect 18732 10558 18734 10610
rect 18786 10558 18788 10610
rect 18508 10498 18564 10510
rect 18508 10446 18510 10498
rect 18562 10446 18564 10498
rect 18228 9996 18340 10052
rect 18396 10052 18452 10062
rect 18172 9986 18228 9996
rect 17388 9874 17444 9884
rect 18396 9826 18452 9996
rect 18396 9774 18398 9826
rect 18450 9774 18452 9826
rect 18396 9762 18452 9774
rect 18508 9826 18564 10446
rect 18732 10388 18788 10558
rect 18732 10322 18788 10332
rect 18844 10164 18900 13020
rect 19068 12962 19124 13692
rect 19068 12910 19070 12962
rect 19122 12910 19124 12962
rect 19068 12898 19124 12910
rect 19180 12852 19236 14478
rect 19292 13076 19348 16604
rect 19628 15988 19684 15998
rect 19628 15894 19684 15932
rect 19404 15540 19460 15550
rect 19404 15446 19460 15484
rect 19516 15316 19572 15326
rect 19516 15222 19572 15260
rect 19740 15204 19796 15214
rect 19740 13972 19796 15148
rect 19852 14642 19908 16940
rect 19964 15538 20020 17724
rect 20188 17332 20244 18510
rect 20412 18452 20468 18956
rect 20860 19010 20916 19068
rect 21980 19124 22036 24558
rect 22764 24722 22820 25228
rect 22876 25218 22932 25228
rect 23100 25060 23156 26796
rect 23548 26290 23604 26908
rect 23548 26238 23550 26290
rect 23602 26238 23604 26290
rect 23548 25732 23604 26238
rect 23660 25732 23716 25742
rect 23548 25730 23716 25732
rect 23548 25678 23662 25730
rect 23714 25678 23716 25730
rect 23548 25676 23716 25678
rect 23660 25666 23716 25676
rect 23436 25506 23492 25518
rect 23436 25454 23438 25506
rect 23490 25454 23492 25506
rect 23436 25060 23492 25454
rect 23156 25004 23492 25060
rect 23548 25284 23604 25294
rect 22764 24670 22766 24722
rect 22818 24670 22820 24722
rect 22316 24500 22372 24510
rect 22764 24500 22820 24670
rect 22988 24722 23044 24734
rect 22988 24670 22990 24722
rect 23042 24670 23044 24722
rect 22316 24498 22820 24500
rect 22316 24446 22318 24498
rect 22370 24446 22820 24498
rect 22316 24444 22820 24446
rect 22316 24434 22372 24444
rect 22316 23716 22372 23726
rect 22316 23622 22372 23660
rect 22316 22146 22372 22158
rect 22316 22094 22318 22146
rect 22370 22094 22372 22146
rect 22092 21700 22148 21710
rect 22092 21606 22148 21644
rect 22316 21476 22372 22094
rect 22092 20804 22148 20814
rect 22092 20710 22148 20748
rect 22316 20690 22372 21420
rect 22316 20638 22318 20690
rect 22370 20638 22372 20690
rect 22316 20018 22372 20638
rect 22540 21476 22596 21486
rect 22764 21476 22820 24444
rect 22876 24610 22932 24622
rect 22876 24558 22878 24610
rect 22930 24558 22932 24610
rect 22876 24052 22932 24558
rect 22988 24612 23044 24670
rect 23100 24722 23156 25004
rect 23100 24670 23102 24722
rect 23154 24670 23156 24722
rect 23100 24658 23156 24670
rect 23324 24836 23380 24846
rect 22988 24546 23044 24556
rect 23212 24612 23268 24622
rect 22876 23986 22932 23996
rect 22988 24164 23044 24174
rect 22988 24050 23044 24108
rect 22988 23998 22990 24050
rect 23042 23998 23044 24050
rect 22988 23986 23044 23998
rect 23100 23940 23156 23950
rect 23100 23846 23156 23884
rect 22988 23716 23044 23726
rect 23212 23716 23268 24556
rect 23324 23938 23380 24780
rect 23324 23886 23326 23938
rect 23378 23886 23380 23938
rect 23324 23874 23380 23886
rect 23044 23660 23268 23716
rect 23548 23828 23604 25228
rect 23884 24052 23940 27022
rect 24332 27076 24388 27086
rect 24332 26982 24388 27020
rect 24556 26964 24612 27692
rect 24892 27860 24948 27870
rect 24556 26514 24612 26908
rect 24780 27188 24836 27198
rect 24780 26964 24836 27132
rect 24780 26870 24836 26908
rect 24556 26462 24558 26514
rect 24610 26462 24612 26514
rect 24556 26450 24612 26462
rect 24108 26180 24164 26190
rect 24108 26086 24164 26124
rect 24892 25508 24948 27804
rect 23996 25396 24052 25406
rect 24556 25396 24612 25406
rect 23996 25394 24612 25396
rect 23996 25342 23998 25394
rect 24050 25342 24558 25394
rect 24610 25342 24612 25394
rect 23996 25340 24612 25342
rect 23996 25330 24052 25340
rect 24556 25330 24612 25340
rect 24892 25394 24948 25452
rect 24892 25342 24894 25394
rect 24946 25342 24948 25394
rect 24892 25330 24948 25342
rect 24444 24836 24500 24846
rect 23996 24612 24052 24622
rect 23996 24518 24052 24556
rect 24444 24164 24500 24780
rect 24892 24836 24948 24846
rect 24892 24612 24948 24780
rect 24444 24098 24500 24108
rect 24780 24610 24948 24612
rect 24780 24558 24894 24610
rect 24946 24558 24948 24610
rect 24780 24556 24948 24558
rect 23884 23996 24276 24052
rect 23660 23884 24052 23940
rect 23660 23828 23716 23884
rect 23548 23826 23716 23828
rect 23548 23774 23550 23826
rect 23602 23774 23716 23826
rect 23548 23772 23716 23774
rect 23996 23826 24052 23884
rect 23996 23774 23998 23826
rect 24050 23774 24052 23826
rect 23548 23716 23604 23772
rect 23996 23762 24052 23774
rect 22988 23622 23044 23660
rect 23548 23650 23604 23660
rect 24220 23604 24276 23996
rect 23996 23548 24276 23604
rect 24444 23716 24500 23726
rect 23548 23044 23604 23054
rect 23548 22950 23604 22988
rect 23660 21700 23716 21710
rect 22540 21474 22820 21476
rect 22540 21422 22542 21474
rect 22594 21422 22820 21474
rect 22540 21420 22820 21422
rect 23100 21476 23156 21486
rect 22540 20244 22596 21420
rect 23100 21382 23156 21420
rect 22988 21028 23044 21038
rect 22988 20914 23044 20972
rect 22988 20862 22990 20914
rect 23042 20862 23044 20914
rect 22988 20850 23044 20862
rect 23548 21028 23604 21038
rect 23548 20802 23604 20972
rect 23548 20750 23550 20802
rect 23602 20750 23604 20802
rect 23548 20738 23604 20750
rect 23660 20804 23716 21644
rect 23996 20914 24052 23548
rect 24108 23154 24164 23166
rect 24108 23102 24110 23154
rect 24162 23102 24164 23154
rect 24108 23044 24164 23102
rect 24444 23156 24500 23660
rect 24780 23604 24836 24556
rect 24892 24546 24948 24556
rect 24892 23828 24948 23838
rect 24892 23734 24948 23772
rect 24780 23548 24948 23604
rect 24668 23156 24724 23166
rect 24444 23154 24724 23156
rect 24444 23102 24670 23154
rect 24722 23102 24724 23154
rect 24444 23100 24724 23102
rect 24108 22484 24164 22988
rect 24220 22484 24276 22494
rect 24108 22482 24500 22484
rect 24108 22430 24222 22482
rect 24274 22430 24500 22482
rect 24108 22428 24500 22430
rect 24220 22418 24276 22428
rect 24444 21924 24500 22428
rect 24444 21810 24500 21868
rect 24444 21758 24446 21810
rect 24498 21758 24500 21810
rect 24444 21746 24500 21758
rect 23996 20862 23998 20914
rect 24050 20862 24052 20914
rect 23996 20850 24052 20862
rect 23660 20738 23716 20748
rect 24220 20804 24276 20814
rect 22540 20178 22596 20188
rect 24220 20130 24276 20748
rect 24556 20578 24612 20590
rect 24556 20526 24558 20578
rect 24610 20526 24612 20578
rect 24556 20468 24612 20526
rect 24556 20402 24612 20412
rect 24220 20078 24222 20130
rect 24274 20078 24276 20130
rect 24220 20066 24276 20078
rect 24668 20132 24724 23100
rect 24780 22260 24836 22270
rect 24780 22166 24836 22204
rect 24892 21812 24948 23548
rect 24780 21756 24948 21812
rect 24780 21028 24836 21756
rect 24780 20962 24836 20972
rect 24892 21588 24948 21598
rect 24668 20066 24724 20076
rect 22316 19966 22318 20018
rect 22370 19966 22372 20018
rect 22204 19796 22260 19806
rect 22204 19346 22260 19740
rect 22316 19460 22372 19966
rect 23548 20020 23604 20030
rect 22764 19906 22820 19918
rect 23548 19908 23604 19964
rect 22764 19854 22766 19906
rect 22818 19854 22820 19906
rect 22316 19394 22372 19404
rect 22652 19460 22708 19470
rect 22204 19294 22206 19346
rect 22258 19294 22260 19346
rect 22204 19236 22260 19294
rect 22652 19346 22708 19404
rect 22652 19294 22654 19346
rect 22706 19294 22708 19346
rect 22652 19282 22708 19294
rect 22204 19170 22260 19180
rect 21980 19058 22036 19068
rect 22764 19124 22820 19854
rect 23436 19906 23604 19908
rect 23436 19854 23550 19906
rect 23602 19854 23604 19906
rect 23436 19852 23604 19854
rect 23436 19236 23492 19852
rect 23548 19842 23604 19852
rect 24108 20018 24164 20030
rect 24108 19966 24110 20018
rect 24162 19966 24164 20018
rect 24108 19460 24164 19966
rect 24332 20020 24388 20030
rect 24332 19926 24388 19964
rect 24780 20018 24836 20030
rect 24780 19966 24782 20018
rect 24834 19966 24836 20018
rect 24780 19460 24836 19966
rect 24108 19404 24388 19460
rect 23436 19142 23492 19180
rect 24108 19234 24164 19246
rect 24108 19182 24110 19234
rect 24162 19182 24164 19234
rect 22764 19058 22820 19068
rect 24108 19124 24164 19182
rect 20860 18958 20862 19010
rect 20914 18958 20916 19010
rect 20532 18844 20796 18854
rect 20588 18788 20636 18844
rect 20692 18788 20740 18844
rect 20532 18778 20796 18788
rect 20636 18452 20692 18462
rect 20412 18450 20692 18452
rect 20412 18398 20638 18450
rect 20690 18398 20692 18450
rect 20412 18396 20692 18398
rect 20636 18386 20692 18396
rect 20412 17892 20468 17902
rect 20412 17778 20468 17836
rect 20412 17726 20414 17778
rect 20466 17726 20468 17778
rect 20412 17714 20468 17726
rect 20188 17266 20244 17276
rect 20532 17276 20796 17286
rect 20588 17220 20636 17276
rect 20692 17220 20740 17276
rect 20532 17210 20796 17220
rect 20188 17108 20244 17118
rect 19964 15486 19966 15538
rect 20018 15486 20020 15538
rect 19964 15474 20020 15486
rect 20076 17052 20188 17108
rect 20076 14644 20132 17052
rect 20188 17014 20244 17052
rect 20412 16772 20468 16782
rect 20300 16212 20356 16222
rect 20188 16210 20356 16212
rect 20188 16158 20302 16210
rect 20354 16158 20356 16210
rect 20188 16156 20356 16158
rect 20188 14868 20244 16156
rect 20300 16146 20356 16156
rect 20412 16098 20468 16716
rect 20636 16772 20692 16782
rect 20636 16678 20692 16716
rect 20412 16046 20414 16098
rect 20466 16046 20468 16098
rect 20300 15988 20356 15998
rect 20300 15204 20356 15932
rect 20300 15138 20356 15148
rect 20412 15148 20468 16046
rect 20860 15986 20916 18958
rect 21196 19012 21252 19022
rect 21196 18676 21252 18956
rect 21196 18610 21252 18620
rect 23436 18676 23492 18686
rect 23436 18582 23492 18620
rect 24108 18676 24164 19068
rect 24220 18676 24276 18686
rect 24164 18674 24276 18676
rect 24164 18622 24222 18674
rect 24274 18622 24276 18674
rect 24164 18620 24276 18622
rect 22204 18564 22260 18574
rect 21868 18450 21924 18462
rect 21868 18398 21870 18450
rect 21922 18398 21924 18450
rect 20972 18340 21028 18350
rect 20972 17778 21028 18284
rect 21420 18338 21476 18350
rect 21420 18286 21422 18338
rect 21474 18286 21476 18338
rect 21420 18228 21476 18286
rect 21868 18340 21924 18398
rect 22204 18340 22260 18508
rect 23548 18564 23604 18574
rect 24108 18544 24164 18620
rect 24220 18610 24276 18620
rect 24332 18674 24388 19404
rect 24780 19394 24836 19404
rect 24332 18622 24334 18674
rect 24386 18622 24388 18674
rect 24332 18610 24388 18622
rect 23548 18470 23604 18508
rect 22876 18452 22932 18462
rect 21868 18274 21924 18284
rect 22092 18338 22260 18340
rect 22092 18286 22206 18338
rect 22258 18286 22260 18338
rect 22092 18284 22260 18286
rect 21420 18162 21476 18172
rect 20972 17726 20974 17778
rect 21026 17726 21028 17778
rect 20972 17714 21028 17726
rect 21868 17554 21924 17566
rect 21868 17502 21870 17554
rect 21922 17502 21924 17554
rect 21868 16996 21924 17502
rect 21868 16930 21924 16940
rect 21980 17442 22036 17454
rect 21980 17390 21982 17442
rect 22034 17390 22036 17442
rect 21532 16884 21588 16894
rect 21532 16790 21588 16828
rect 21980 16884 22036 17390
rect 21980 16818 22036 16828
rect 22092 16658 22148 18284
rect 22204 18274 22260 18284
rect 22316 18450 22932 18452
rect 22316 18398 22878 18450
rect 22930 18398 22932 18450
rect 22316 18396 22932 18398
rect 22204 17668 22260 17678
rect 22316 17668 22372 18396
rect 22876 18386 22932 18396
rect 23324 18450 23380 18462
rect 23324 18398 23326 18450
rect 23378 18398 23380 18450
rect 23324 18340 23380 18398
rect 24892 18452 24948 21532
rect 25004 19458 25060 29932
rect 25116 29988 25172 29998
rect 25116 20804 25172 29932
rect 25228 29988 25284 30716
rect 25340 30324 25396 31502
rect 26908 31220 26964 31838
rect 26684 31108 26740 31118
rect 26908 31108 26964 31164
rect 25340 30258 25396 30268
rect 25788 31052 26068 31108
rect 25788 30210 25844 31052
rect 26012 30994 26068 31052
rect 26684 31106 26964 31108
rect 26684 31054 26686 31106
rect 26738 31054 26964 31106
rect 26684 31052 26964 31054
rect 26684 31042 26740 31052
rect 26012 30942 26014 30994
rect 26066 30942 26068 30994
rect 26012 30930 26068 30942
rect 26348 30996 26404 31006
rect 25900 30882 25956 30894
rect 25900 30830 25902 30882
rect 25954 30830 25956 30882
rect 25900 30324 25956 30830
rect 26012 30324 26068 30334
rect 25900 30268 26012 30324
rect 26012 30230 26068 30268
rect 25788 30158 25790 30210
rect 25842 30158 25844 30210
rect 25788 29988 25844 30158
rect 26348 30210 26404 30940
rect 26348 30158 26350 30210
rect 26402 30158 26404 30210
rect 26348 30146 26404 30158
rect 25228 29986 25844 29988
rect 25228 29934 25230 29986
rect 25282 29934 25844 29986
rect 25228 29932 25844 29934
rect 26908 29986 26964 29998
rect 26908 29934 26910 29986
rect 26962 29934 26964 29986
rect 25228 28308 25284 29932
rect 26908 29764 26964 29934
rect 26908 29698 26964 29708
rect 26908 29540 26964 29550
rect 26908 29446 26964 29484
rect 25900 29316 25956 29326
rect 25788 29314 25956 29316
rect 25788 29262 25902 29314
rect 25954 29262 25956 29314
rect 25788 29260 25956 29262
rect 25564 28756 25620 28766
rect 25564 28642 25620 28700
rect 25564 28590 25566 28642
rect 25618 28590 25620 28642
rect 25564 28578 25620 28590
rect 25788 28420 25844 29260
rect 25900 29250 25956 29260
rect 26348 29316 26404 29326
rect 26348 28644 26404 29260
rect 27020 28754 27076 33068
rect 27468 32564 27524 32574
rect 27468 32470 27524 32508
rect 27580 32450 27636 32462
rect 27580 32398 27582 32450
rect 27634 32398 27636 32450
rect 27580 32340 27636 32398
rect 28252 32450 28308 33292
rect 28476 33124 28532 33134
rect 28476 33030 28532 33068
rect 28252 32398 28254 32450
rect 28306 32398 28308 32450
rect 28252 32386 28308 32398
rect 27580 32002 27636 32284
rect 27580 31950 27582 32002
rect 27634 31950 27636 32002
rect 27580 31938 27636 31950
rect 27244 31780 27300 31790
rect 27244 31778 27412 31780
rect 27244 31726 27246 31778
rect 27298 31726 27412 31778
rect 27244 31724 27412 31726
rect 27244 31714 27300 31724
rect 27244 30996 27300 31006
rect 27356 30996 27412 31724
rect 27692 31556 27748 31566
rect 27692 31218 27748 31500
rect 27692 31166 27694 31218
rect 27746 31166 27748 31218
rect 27692 31154 27748 31166
rect 27804 31220 27860 31230
rect 27804 31106 27860 31164
rect 27804 31054 27806 31106
rect 27858 31054 27860 31106
rect 27804 31042 27860 31054
rect 27468 30996 27524 31006
rect 27356 30994 27524 30996
rect 27356 30942 27470 30994
rect 27522 30942 27524 30994
rect 27356 30940 27524 30942
rect 27244 30902 27300 30940
rect 27356 29988 27412 29998
rect 27020 28702 27022 28754
rect 27074 28702 27076 28754
rect 27020 28690 27076 28702
rect 27244 29986 27412 29988
rect 27244 29934 27358 29986
rect 27410 29934 27412 29986
rect 27244 29932 27412 29934
rect 26460 28644 26516 28654
rect 26348 28642 26516 28644
rect 26348 28590 26462 28642
rect 26514 28590 26516 28642
rect 26348 28588 26516 28590
rect 26460 28578 26516 28588
rect 25900 28532 25956 28542
rect 25900 28438 25956 28476
rect 26796 28532 26852 28542
rect 25788 28326 25844 28364
rect 26796 28418 26852 28476
rect 26796 28366 26798 28418
rect 26850 28366 26852 28418
rect 25228 28242 25284 28252
rect 26796 27970 26852 28366
rect 26796 27918 26798 27970
rect 26850 27918 26852 27970
rect 26012 27860 26068 27870
rect 25564 27748 25620 27758
rect 25228 27076 25284 27086
rect 25228 26982 25284 27020
rect 25564 26516 25620 27692
rect 26012 27746 26068 27804
rect 26572 27860 26628 27870
rect 26572 27766 26628 27804
rect 26012 27694 26014 27746
rect 26066 27694 26068 27746
rect 26012 27076 26068 27694
rect 26796 27188 26852 27918
rect 26012 27010 26068 27020
rect 26572 27132 26852 27188
rect 27020 28420 27076 28430
rect 26572 27074 26628 27132
rect 26572 27022 26574 27074
rect 26626 27022 26628 27074
rect 26124 26964 26180 26974
rect 26012 26852 26180 26908
rect 26012 26850 26068 26852
rect 26012 26798 26014 26850
rect 26066 26798 26068 26850
rect 26012 26786 26068 26798
rect 25564 26384 25620 26460
rect 25676 25956 25732 25966
rect 25676 25620 25732 25900
rect 25676 25488 25732 25564
rect 25228 25396 25284 25406
rect 25228 23268 25284 25340
rect 26236 25396 26292 25406
rect 26236 25302 26292 25340
rect 26572 25172 26628 27022
rect 26684 26964 26740 26974
rect 26684 26870 26740 26908
rect 26908 26852 26964 26862
rect 26908 26758 26964 26796
rect 26796 26628 26852 26638
rect 26796 25620 26852 26572
rect 27020 26516 27076 28364
rect 27244 27860 27300 29932
rect 27356 29922 27412 29932
rect 27356 29764 27412 29774
rect 27356 29426 27412 29708
rect 27468 29540 27524 30940
rect 28140 29986 28196 29998
rect 28140 29934 28142 29986
rect 28194 29934 28196 29986
rect 28140 29652 28196 29934
rect 27468 29474 27524 29484
rect 27580 29596 28196 29652
rect 28588 29764 28644 29774
rect 28588 29650 28644 29708
rect 28588 29598 28590 29650
rect 28642 29598 28644 29650
rect 27356 29374 27358 29426
rect 27410 29374 27412 29426
rect 27356 28980 27412 29374
rect 27356 28914 27412 28924
rect 27580 28530 27636 29596
rect 28588 29586 28644 29598
rect 28700 29652 28756 33964
rect 30192 33740 30456 33750
rect 30248 33684 30296 33740
rect 30352 33684 30400 33740
rect 30192 33674 30456 33684
rect 30604 33570 30660 34748
rect 30716 34468 30772 34478
rect 30716 34354 30772 34412
rect 30716 34302 30718 34354
rect 30770 34302 30772 34354
rect 30716 34290 30772 34302
rect 31276 34242 31332 34748
rect 31500 34468 31556 35868
rect 32060 35138 32116 35868
rect 32396 35812 32452 35822
rect 32396 35698 32452 35756
rect 32396 35646 32398 35698
rect 32450 35646 32452 35698
rect 32396 35634 32452 35646
rect 32060 35086 32062 35138
rect 32114 35086 32116 35138
rect 32060 35074 32116 35086
rect 31500 34354 31556 34412
rect 31500 34302 31502 34354
rect 31554 34302 31556 34354
rect 31500 34290 31556 34302
rect 32620 34690 32676 36428
rect 32732 35924 32788 35934
rect 32732 35698 32788 35868
rect 33964 35922 34020 36652
rect 34076 36594 34132 38108
rect 36204 37492 36260 39200
rect 38668 37492 38724 39200
rect 40236 38052 40292 38062
rect 36204 37436 36596 37492
rect 38668 37436 39060 37492
rect 34076 36542 34078 36594
rect 34130 36542 34132 36594
rect 34076 36530 34132 36542
rect 35196 36596 35252 36606
rect 34972 36484 35028 36494
rect 33964 35870 33966 35922
rect 34018 35870 34020 35922
rect 33964 35858 34020 35870
rect 34860 36372 34916 36382
rect 34860 35812 34916 36316
rect 32732 35646 32734 35698
rect 32786 35646 32788 35698
rect 32732 35634 32788 35646
rect 32844 35700 32900 35710
rect 32844 35606 32900 35644
rect 33628 35700 33684 35710
rect 34860 35680 34916 35756
rect 34972 35924 35028 36428
rect 35196 36482 35252 36540
rect 35196 36430 35198 36482
rect 35250 36430 35252 36482
rect 35196 36418 35252 36430
rect 35644 36484 35700 36494
rect 35644 36390 35700 36428
rect 35868 36484 35924 36494
rect 35868 36390 35924 36428
rect 36204 36482 36260 36494
rect 36204 36430 36206 36482
rect 36258 36430 36260 36482
rect 36092 36372 36148 36382
rect 36092 36278 36148 36316
rect 34972 35810 35028 35868
rect 34972 35758 34974 35810
rect 35026 35758 35028 35810
rect 34972 35746 35028 35758
rect 35084 35698 35140 35710
rect 33628 35606 33684 35644
rect 35084 35646 35086 35698
rect 35138 35646 35140 35698
rect 34748 34916 34804 34926
rect 34748 34822 34804 34860
rect 35084 34804 35140 35646
rect 35532 35476 35588 35486
rect 35532 35382 35588 35420
rect 35084 34738 35140 34748
rect 35196 34914 35252 34926
rect 35196 34862 35198 34914
rect 35250 34862 35252 34914
rect 32620 34638 32622 34690
rect 32674 34638 32676 34690
rect 31276 34190 31278 34242
rect 31330 34190 31332 34242
rect 31276 34178 31332 34190
rect 32620 34244 32676 34638
rect 33852 34356 33908 34366
rect 33852 34262 33908 34300
rect 32620 34178 32676 34188
rect 32060 34132 32116 34142
rect 31612 33908 31668 33918
rect 31612 33814 31668 33852
rect 30604 33518 30606 33570
rect 30658 33518 30660 33570
rect 30604 33506 30660 33518
rect 29932 33458 29988 33470
rect 29932 33406 29934 33458
rect 29986 33406 29988 33458
rect 28924 33348 28980 33358
rect 28924 33346 29540 33348
rect 28924 33294 28926 33346
rect 28978 33294 29540 33346
rect 28924 33292 29540 33294
rect 28924 33282 28980 33292
rect 29484 32786 29540 33292
rect 29820 33346 29876 33358
rect 29820 33294 29822 33346
rect 29874 33294 29876 33346
rect 29820 33124 29876 33294
rect 29932 33348 29988 33406
rect 32060 33458 32116 34076
rect 32060 33406 32062 33458
rect 32114 33406 32116 33458
rect 32060 33394 32116 33406
rect 32844 34132 32900 34142
rect 29932 33282 29988 33292
rect 32844 33346 32900 34076
rect 33740 34130 33796 34142
rect 33740 34078 33742 34130
rect 33794 34078 33796 34130
rect 32844 33294 32846 33346
rect 32898 33294 32900 33346
rect 32844 33282 32900 33294
rect 33516 33346 33572 33358
rect 33516 33294 33518 33346
rect 33570 33294 33572 33346
rect 29820 33058 29876 33068
rect 31836 33124 31892 33134
rect 29484 32734 29486 32786
rect 29538 32734 29540 32786
rect 29484 32722 29540 32734
rect 28924 32564 28980 32574
rect 28924 32470 28980 32508
rect 31164 32562 31220 32574
rect 31164 32510 31166 32562
rect 31218 32510 31220 32562
rect 29148 32340 29204 32350
rect 29148 32246 29204 32284
rect 30192 32172 30456 32182
rect 30248 32116 30296 32172
rect 30352 32116 30400 32172
rect 30192 32106 30456 32116
rect 31164 32004 31220 32510
rect 31500 32562 31556 32574
rect 31500 32510 31502 32562
rect 31554 32510 31556 32562
rect 31388 32452 31444 32462
rect 31388 32358 31444 32396
rect 31500 31948 31556 32510
rect 31724 32562 31780 32574
rect 31724 32510 31726 32562
rect 31778 32510 31780 32562
rect 30940 31892 31220 31948
rect 31276 31892 31556 31948
rect 31612 32004 31668 32014
rect 30604 31554 30660 31566
rect 30604 31502 30606 31554
rect 30658 31502 30660 31554
rect 29596 30996 29652 31006
rect 29596 30882 29652 30940
rect 30492 30996 30548 31006
rect 30492 30902 30548 30940
rect 29596 30830 29598 30882
rect 29650 30830 29652 30882
rect 29372 30212 29428 30222
rect 28812 29988 28868 29998
rect 28812 29894 28868 29932
rect 28812 29652 28868 29662
rect 28700 29650 28868 29652
rect 28700 29598 28814 29650
rect 28866 29598 28868 29650
rect 28700 29596 28868 29598
rect 28812 29586 28868 29596
rect 27804 29428 27860 29438
rect 28476 29428 28532 29438
rect 27804 29426 28532 29428
rect 27804 29374 27806 29426
rect 27858 29374 28478 29426
rect 28530 29374 28532 29426
rect 27804 29372 28532 29374
rect 27804 29362 27860 29372
rect 28476 28868 28532 29372
rect 28812 29428 28868 29438
rect 28476 28812 28644 28868
rect 28476 28644 28532 28654
rect 27580 28478 27582 28530
rect 27634 28478 27636 28530
rect 27580 28420 27636 28478
rect 28140 28532 28196 28542
rect 27580 28354 27636 28364
rect 27692 28418 27748 28430
rect 27692 28366 27694 28418
rect 27746 28366 27748 28418
rect 27356 27860 27412 27870
rect 27244 27858 27412 27860
rect 27244 27806 27358 27858
rect 27410 27806 27412 27858
rect 27244 27804 27412 27806
rect 27356 27748 27412 27804
rect 27356 27682 27412 27692
rect 27692 27748 27748 28366
rect 27916 28418 27972 28430
rect 27916 28366 27918 28418
rect 27970 28366 27972 28418
rect 27916 27972 27972 28366
rect 27916 27906 27972 27916
rect 28028 28420 28084 28430
rect 27692 27682 27748 27692
rect 28028 27858 28084 28364
rect 28028 27806 28030 27858
rect 28082 27806 28084 27858
rect 27692 27076 27748 27086
rect 27692 27074 27860 27076
rect 27692 27022 27694 27074
rect 27746 27022 27860 27074
rect 27692 27020 27860 27022
rect 27692 27010 27748 27020
rect 27020 26450 27076 26460
rect 27356 26962 27412 26974
rect 27356 26910 27358 26962
rect 27410 26910 27412 26962
rect 26684 25396 26740 25406
rect 26684 25302 26740 25340
rect 26796 25394 26852 25564
rect 26796 25342 26798 25394
rect 26850 25342 26852 25394
rect 26796 25330 26852 25342
rect 26908 25956 26964 25966
rect 26908 25172 26964 25900
rect 27356 25956 27412 26910
rect 27468 26850 27524 26862
rect 27468 26798 27470 26850
rect 27522 26798 27524 26850
rect 27468 26290 27524 26798
rect 27692 26292 27748 26302
rect 27468 26238 27470 26290
rect 27522 26238 27524 26290
rect 27468 26226 27524 26238
rect 27580 26290 27748 26292
rect 27580 26238 27694 26290
rect 27746 26238 27748 26290
rect 27580 26236 27748 26238
rect 27356 25890 27412 25900
rect 27468 25732 27524 25742
rect 27580 25732 27636 26236
rect 27692 26226 27748 26236
rect 27020 25730 27636 25732
rect 27020 25678 27470 25730
rect 27522 25678 27636 25730
rect 27020 25676 27636 25678
rect 27692 25956 27748 25966
rect 27020 25506 27076 25676
rect 27468 25666 27524 25676
rect 27692 25618 27748 25900
rect 27692 25566 27694 25618
rect 27746 25566 27748 25618
rect 27692 25554 27748 25566
rect 27020 25454 27022 25506
rect 27074 25454 27076 25506
rect 27020 25442 27076 25454
rect 27580 25508 27636 25518
rect 26236 25116 26740 25172
rect 26124 24836 26180 24846
rect 26124 24742 26180 24780
rect 25676 24724 25732 24734
rect 25564 24612 25620 24622
rect 25452 24556 25564 24612
rect 25452 23828 25508 24556
rect 25564 24480 25620 24556
rect 25452 23734 25508 23772
rect 25676 23828 25732 24668
rect 26012 24052 26068 24062
rect 26012 23958 26068 23996
rect 25228 23202 25284 23212
rect 25676 23714 25732 23772
rect 26124 23940 26180 23950
rect 26236 23940 26292 25116
rect 26684 24834 26740 25116
rect 26684 24782 26686 24834
rect 26738 24782 26740 24834
rect 26684 24770 26740 24782
rect 26796 25116 26964 25172
rect 27132 25396 27188 25406
rect 26348 24724 26404 24734
rect 26348 24630 26404 24668
rect 26572 24722 26628 24734
rect 26572 24670 26574 24722
rect 26626 24670 26628 24722
rect 26572 24612 26628 24670
rect 26124 23938 26516 23940
rect 26124 23886 26126 23938
rect 26178 23886 26516 23938
rect 26124 23884 26516 23886
rect 25676 23662 25678 23714
rect 25730 23662 25732 23714
rect 25228 22260 25284 22270
rect 25676 22260 25732 23662
rect 25900 23716 25956 23726
rect 25900 23622 25956 23660
rect 26124 23492 26180 23884
rect 25788 23436 26180 23492
rect 25788 22482 25844 23436
rect 25900 23268 25956 23278
rect 25900 23174 25956 23212
rect 25788 22430 25790 22482
rect 25842 22430 25844 22482
rect 25788 22418 25844 22430
rect 25676 22204 25844 22260
rect 25228 22166 25284 22204
rect 25676 21924 25732 21934
rect 25676 21698 25732 21868
rect 25676 21646 25678 21698
rect 25730 21646 25732 21698
rect 25676 21634 25732 21646
rect 25788 21588 25844 22204
rect 26124 21812 26180 23436
rect 26460 23266 26516 23884
rect 26572 23492 26628 24556
rect 26684 24612 26740 24622
rect 26796 24612 26852 25116
rect 26684 24610 26852 24612
rect 26684 24558 26686 24610
rect 26738 24558 26852 24610
rect 26684 24556 26852 24558
rect 26684 24546 26740 24556
rect 26796 23716 26852 23726
rect 26572 23426 26628 23436
rect 26684 23714 26852 23716
rect 26684 23662 26798 23714
rect 26850 23662 26852 23714
rect 26684 23660 26852 23662
rect 26460 23214 26462 23266
rect 26514 23214 26516 23266
rect 26460 23202 26516 23214
rect 26572 23268 26628 23278
rect 26572 23174 26628 23212
rect 26684 22932 26740 23660
rect 26796 23650 26852 23660
rect 26908 23716 26964 23726
rect 26908 23622 26964 23660
rect 27020 23714 27076 23726
rect 27020 23662 27022 23714
rect 27074 23662 27076 23714
rect 27020 23492 27076 23662
rect 26796 23436 27076 23492
rect 26796 23378 26852 23436
rect 26796 23326 26798 23378
rect 26850 23326 26852 23378
rect 26796 23314 26852 23326
rect 26572 22876 26740 22932
rect 26348 22260 26404 22270
rect 26348 22166 26404 22204
rect 26460 22146 26516 22158
rect 26460 22094 26462 22146
rect 26514 22094 26516 22146
rect 26460 21924 26516 22094
rect 26460 21858 26516 21868
rect 26236 21812 26292 21822
rect 26124 21810 26292 21812
rect 26124 21758 26238 21810
rect 26290 21758 26292 21810
rect 26124 21756 26292 21758
rect 26236 21746 26292 21756
rect 25900 21588 25956 21598
rect 25788 21586 25956 21588
rect 25788 21534 25902 21586
rect 25954 21534 25956 21586
rect 25788 21532 25956 21534
rect 25116 20738 25172 20748
rect 25788 21028 25844 21038
rect 25564 20692 25620 20702
rect 25564 20598 25620 20636
rect 25004 19406 25006 19458
rect 25058 19406 25060 19458
rect 25004 19394 25060 19406
rect 25116 20580 25172 20590
rect 24892 18320 24948 18396
rect 25004 19236 25060 19246
rect 23324 18274 23380 18284
rect 22764 18228 22820 18238
rect 22764 17778 22820 18172
rect 24444 18226 24500 18238
rect 24444 18174 24446 18226
rect 24498 18174 24500 18226
rect 24444 18116 24500 18174
rect 25004 18116 25060 19180
rect 24444 18060 25060 18116
rect 22764 17726 22766 17778
rect 22818 17726 22820 17778
rect 22764 17714 22820 17726
rect 22204 17666 22372 17668
rect 22204 17614 22206 17666
rect 22258 17614 22372 17666
rect 22204 17612 22372 17614
rect 22204 17602 22260 17612
rect 22204 16996 22260 17006
rect 22204 16882 22260 16940
rect 22204 16830 22206 16882
rect 22258 16830 22260 16882
rect 22204 16818 22260 16830
rect 24332 16882 24388 16894
rect 24332 16830 24334 16882
rect 24386 16830 24388 16882
rect 22092 16606 22094 16658
rect 22146 16606 22148 16658
rect 22092 16594 22148 16606
rect 22876 16770 22932 16782
rect 22876 16718 22878 16770
rect 22930 16718 22932 16770
rect 21644 16100 21700 16110
rect 21644 16006 21700 16044
rect 22204 16098 22260 16110
rect 22204 16046 22206 16098
rect 22258 16046 22260 16098
rect 20860 15934 20862 15986
rect 20914 15934 20916 15986
rect 20636 15876 20692 15914
rect 20636 15810 20692 15820
rect 20532 15708 20796 15718
rect 20588 15652 20636 15708
rect 20692 15652 20740 15708
rect 20532 15642 20796 15652
rect 20636 15540 20692 15550
rect 20860 15540 20916 15934
rect 20636 15538 20916 15540
rect 20636 15486 20638 15538
rect 20690 15486 20916 15538
rect 20636 15484 20916 15486
rect 21084 15540 21140 15550
rect 21532 15540 21588 15550
rect 20636 15474 20692 15484
rect 21084 15426 21140 15484
rect 21084 15374 21086 15426
rect 21138 15374 21140 15426
rect 21084 15316 21140 15374
rect 21084 15250 21140 15260
rect 21196 15538 21588 15540
rect 21196 15486 21534 15538
rect 21586 15486 21588 15538
rect 21196 15484 21588 15486
rect 21196 15148 21252 15484
rect 20412 15092 21252 15148
rect 21308 15316 21364 15326
rect 20188 14812 20468 14868
rect 20300 14644 20356 14654
rect 19852 14590 19854 14642
rect 19906 14590 19908 14642
rect 19852 14578 19908 14590
rect 19964 14642 20356 14644
rect 19964 14590 20302 14642
rect 20354 14590 20356 14642
rect 19964 14588 20356 14590
rect 19852 13972 19908 13982
rect 19740 13970 19908 13972
rect 19740 13918 19854 13970
rect 19906 13918 19908 13970
rect 19740 13916 19908 13918
rect 19740 13524 19796 13916
rect 19852 13906 19908 13916
rect 19740 13458 19796 13468
rect 19292 13010 19348 13020
rect 19404 12964 19460 12974
rect 19404 12870 19460 12908
rect 19180 12786 19236 12796
rect 19292 12740 19348 12750
rect 19292 12646 19348 12684
rect 19964 12740 20020 14588
rect 20300 14578 20356 14588
rect 20412 12962 20468 14812
rect 20860 14642 20916 15092
rect 20860 14590 20862 14642
rect 20914 14590 20916 14642
rect 20860 14578 20916 14590
rect 20532 14140 20796 14150
rect 20588 14084 20636 14140
rect 20692 14084 20740 14140
rect 20532 14074 20796 14084
rect 20972 13748 21028 13758
rect 20972 13654 21028 13692
rect 20860 13634 20916 13646
rect 20860 13582 20862 13634
rect 20914 13582 20916 13634
rect 20412 12910 20414 12962
rect 20466 12910 20468 12962
rect 20412 12898 20468 12910
rect 20748 12964 20804 12974
rect 20860 12964 20916 13582
rect 20748 12962 20916 12964
rect 20748 12910 20750 12962
rect 20802 12910 20916 12962
rect 20748 12908 20916 12910
rect 20748 12898 20804 12908
rect 20300 12852 20356 12862
rect 20300 12758 20356 12796
rect 19068 12404 19124 12414
rect 19068 12310 19124 12348
rect 19292 12404 19348 12414
rect 19292 12310 19348 12348
rect 19852 12404 19908 12414
rect 19964 12404 20020 12684
rect 19852 12402 20020 12404
rect 19852 12350 19854 12402
rect 19906 12350 20020 12402
rect 19852 12348 20020 12350
rect 19852 12338 19908 12348
rect 18956 12180 19012 12190
rect 19964 12180 20020 12348
rect 18956 12178 19124 12180
rect 18956 12126 18958 12178
rect 19010 12126 19124 12178
rect 18956 12124 19124 12126
rect 18956 12114 19012 12124
rect 18956 11956 19012 11966
rect 18956 11394 19012 11900
rect 18956 11342 18958 11394
rect 19010 11342 19012 11394
rect 18956 11330 19012 11342
rect 19068 11284 19124 12124
rect 19068 10500 19124 11228
rect 19068 10434 19124 10444
rect 19292 11620 19348 11630
rect 18508 9774 18510 9826
rect 18562 9774 18564 9826
rect 18508 9762 18564 9774
rect 18732 10108 18900 10164
rect 17276 9714 17332 9726
rect 18172 9716 18228 9726
rect 17276 9662 17278 9714
rect 17330 9662 17332 9714
rect 17276 9604 17332 9662
rect 17500 9714 18228 9716
rect 17500 9662 18174 9714
rect 18226 9662 18228 9714
rect 17500 9660 18228 9662
rect 17276 9538 17332 9548
rect 17388 9602 17444 9614
rect 17388 9550 17390 9602
rect 17442 9550 17444 9602
rect 17388 9492 17444 9550
rect 17388 9426 17444 9436
rect 17164 8428 17332 8484
rect 15820 7298 15876 7308
rect 15596 6692 15652 6702
rect 15596 6598 15652 6636
rect 16044 6692 16100 6702
rect 15092 6524 15204 6580
rect 14812 6468 14868 6478
rect 15092 6468 15148 6524
rect 14868 6412 15148 6468
rect 14700 5796 14756 5806
rect 14700 5702 14756 5740
rect 14812 5572 14868 6412
rect 15484 6132 15540 6142
rect 15484 6130 15988 6132
rect 15484 6078 15486 6130
rect 15538 6078 15988 6130
rect 15484 6076 15988 6078
rect 15484 6066 15540 6076
rect 15820 5906 15876 5918
rect 15820 5854 15822 5906
rect 15874 5854 15876 5906
rect 14700 5516 14868 5572
rect 14924 5572 14980 5582
rect 14700 2212 14756 5516
rect 14924 5236 14980 5516
rect 14812 5234 14980 5236
rect 14812 5182 14926 5234
rect 14978 5182 14980 5234
rect 14812 5180 14980 5182
rect 14812 4450 14868 5180
rect 14924 5170 14980 5180
rect 15036 5124 15092 5134
rect 15036 4900 15092 5068
rect 15148 5124 15204 5134
rect 15820 5124 15876 5854
rect 15932 5908 15988 6076
rect 16044 6130 16100 6636
rect 16044 6078 16046 6130
rect 16098 6078 16100 6130
rect 16044 6066 16100 6078
rect 16156 6018 16212 8428
rect 16604 8260 16660 8270
rect 16604 8166 16660 8204
rect 17164 8260 17220 8270
rect 16604 7700 16660 7710
rect 16268 7362 16324 7374
rect 16268 7310 16270 7362
rect 16322 7310 16324 7362
rect 16268 6692 16324 7310
rect 16604 6692 16660 7644
rect 16828 7364 16884 7374
rect 16828 7362 16996 7364
rect 16828 7310 16830 7362
rect 16882 7310 16996 7362
rect 16828 7308 16996 7310
rect 16828 7298 16884 7308
rect 16324 6636 16436 6692
rect 16268 6626 16324 6636
rect 16156 5966 16158 6018
rect 16210 5966 16212 6018
rect 16156 5908 16212 5966
rect 15932 5852 16212 5908
rect 16268 6466 16324 6478
rect 16268 6414 16270 6466
rect 16322 6414 16324 6466
rect 16268 5236 16324 6414
rect 16268 5170 16324 5180
rect 15148 5122 15652 5124
rect 15148 5070 15150 5122
rect 15202 5070 15652 5122
rect 15148 5068 15652 5070
rect 15148 5058 15204 5068
rect 15036 4844 15316 4900
rect 14812 4398 14814 4450
rect 14866 4398 14868 4450
rect 14812 4386 14868 4398
rect 14924 4338 14980 4350
rect 14924 4286 14926 4338
rect 14978 4286 14980 4338
rect 14924 4228 14980 4286
rect 14924 3556 14980 4172
rect 14924 3490 14980 3500
rect 15036 3780 15092 3790
rect 15036 3444 15092 3724
rect 15260 3554 15316 4844
rect 15484 4898 15540 4910
rect 15484 4846 15486 4898
rect 15538 4846 15540 4898
rect 15260 3502 15262 3554
rect 15314 3502 15316 3554
rect 15260 3490 15316 3502
rect 15372 4116 15428 4126
rect 15036 3378 15092 3388
rect 15148 3332 15204 3342
rect 15372 3332 15428 4060
rect 15484 3666 15540 4846
rect 15596 4900 15652 5068
rect 15820 5058 15876 5068
rect 16380 5124 16436 6636
rect 16604 6690 16884 6692
rect 16604 6638 16606 6690
rect 16658 6638 16884 6690
rect 16604 6636 16884 6638
rect 16604 6626 16660 6636
rect 16492 6466 16548 6478
rect 16492 6414 16494 6466
rect 16546 6414 16548 6466
rect 16492 5908 16548 6414
rect 16828 6130 16884 6636
rect 16828 6078 16830 6130
rect 16882 6078 16884 6130
rect 16828 6066 16884 6078
rect 16492 5842 16548 5852
rect 16940 5572 16996 7308
rect 16940 5506 16996 5516
rect 16380 5012 16436 5068
rect 16716 5236 16772 5246
rect 16492 5012 16548 5022
rect 16380 5010 16548 5012
rect 16380 4958 16494 5010
rect 16546 4958 16548 5010
rect 16380 4956 16548 4958
rect 16268 4900 16324 4910
rect 15596 4898 16324 4900
rect 15596 4846 16270 4898
rect 16322 4846 16324 4898
rect 15596 4844 16324 4846
rect 16268 4450 16324 4844
rect 16380 4564 16436 4574
rect 16380 4470 16436 4508
rect 16268 4398 16270 4450
rect 16322 4398 16324 4450
rect 16268 4386 16324 4398
rect 15484 3614 15486 3666
rect 15538 3614 15540 3666
rect 15484 3602 15540 3614
rect 15708 3556 15764 3566
rect 15708 3462 15764 3500
rect 15148 3330 15428 3332
rect 15148 3278 15150 3330
rect 15202 3278 15428 3330
rect 15148 3276 15428 3278
rect 16268 3332 16324 3342
rect 15148 3266 15204 3276
rect 16268 3238 16324 3276
rect 14700 2146 14756 2156
rect 16492 1316 16548 4956
rect 16604 5012 16660 5022
rect 16604 4918 16660 4956
rect 16492 1250 16548 1260
rect 16604 3556 16660 3566
rect 16716 3556 16772 5180
rect 17052 5124 17108 5134
rect 17052 5030 17108 5068
rect 17164 5012 17220 8204
rect 17276 8036 17332 8428
rect 17500 8260 17556 9660
rect 18172 9650 18228 9660
rect 18284 9602 18340 9614
rect 18284 9550 18286 9602
rect 18338 9550 18340 9602
rect 17948 9380 18004 9390
rect 17500 8258 17780 8260
rect 17500 8206 17502 8258
rect 17554 8206 17780 8258
rect 17500 8204 17780 8206
rect 17500 8194 17556 8204
rect 17276 8034 17668 8036
rect 17276 7982 17278 8034
rect 17330 7982 17668 8034
rect 17276 7980 17668 7982
rect 17276 7970 17332 7980
rect 17612 7698 17668 7980
rect 17612 7646 17614 7698
rect 17666 7646 17668 7698
rect 17612 7634 17668 7646
rect 17724 6690 17780 8204
rect 17724 6638 17726 6690
rect 17778 6638 17780 6690
rect 17724 6626 17780 6638
rect 17612 5908 17668 5918
rect 17612 5794 17668 5852
rect 17612 5742 17614 5794
rect 17666 5742 17668 5794
rect 17500 5124 17556 5134
rect 17612 5124 17668 5742
rect 17948 5684 18004 9324
rect 18172 9268 18228 9278
rect 18060 9044 18116 9054
rect 18060 8950 18116 8988
rect 18172 7140 18228 9212
rect 18284 9156 18340 9550
rect 18284 8258 18340 9100
rect 18284 8206 18286 8258
rect 18338 8206 18340 8258
rect 18284 8194 18340 8206
rect 18396 9492 18452 9502
rect 18396 7252 18452 9436
rect 18620 9042 18676 9054
rect 18620 8990 18622 9042
rect 18674 8990 18676 9042
rect 18620 8932 18676 8990
rect 18620 8260 18676 8876
rect 18620 8194 18676 8204
rect 18508 8036 18564 8046
rect 18508 7474 18564 7980
rect 18508 7422 18510 7474
rect 18562 7422 18564 7474
rect 18508 7410 18564 7422
rect 18396 7196 18564 7252
rect 18172 7084 18452 7140
rect 18060 6692 18116 6702
rect 18060 6690 18340 6692
rect 18060 6638 18062 6690
rect 18114 6638 18340 6690
rect 18060 6636 18340 6638
rect 18060 6626 18116 6636
rect 18284 5908 18340 6636
rect 18284 5814 18340 5852
rect 17948 5628 18340 5684
rect 17724 5124 17780 5134
rect 17612 5068 17724 5124
rect 17500 5030 17556 5068
rect 17724 5058 17780 5068
rect 17052 4564 17108 4574
rect 17164 4564 17220 4956
rect 17052 4562 17220 4564
rect 17052 4510 17054 4562
rect 17106 4510 17220 4562
rect 17052 4508 17220 4510
rect 17948 4898 18004 4910
rect 17948 4846 17950 4898
rect 18002 4846 18004 4898
rect 17052 4498 17108 4508
rect 17948 4340 18004 4846
rect 17612 4338 18004 4340
rect 17612 4286 17950 4338
rect 18002 4286 18004 4338
rect 17612 4284 18004 4286
rect 16604 3554 16772 3556
rect 16604 3502 16606 3554
rect 16658 3502 16772 3554
rect 16604 3500 16772 3502
rect 17500 3556 17556 3566
rect 14476 914 14532 924
rect 15484 924 15764 980
rect 15484 800 15540 924
rect 2688 0 2800 800
rect 4816 0 4928 800
rect 6944 0 7056 800
rect 9072 0 9184 800
rect 11200 0 11312 800
rect 13328 0 13440 800
rect 15456 0 15568 800
rect 15708 756 15764 924
rect 16604 868 16660 3500
rect 17500 1652 17556 3500
rect 17500 1586 17556 1596
rect 16268 812 16660 868
rect 16268 756 16324 812
rect 17612 800 17668 4284
rect 17948 4274 18004 4284
rect 18284 4452 18340 5628
rect 18284 4226 18340 4396
rect 18284 4174 18286 4226
rect 18338 4174 18340 4226
rect 18284 4162 18340 4174
rect 18396 3668 18452 7084
rect 18508 6020 18564 7196
rect 18508 5926 18564 5964
rect 18620 5906 18676 5918
rect 18620 5854 18622 5906
rect 18674 5854 18676 5906
rect 18620 5124 18676 5854
rect 18732 5796 18788 10108
rect 18844 9940 18900 9950
rect 18844 9846 18900 9884
rect 19292 9380 19348 11564
rect 19628 10724 19684 10734
rect 19516 10610 19572 10622
rect 19516 10558 19518 10610
rect 19570 10558 19572 10610
rect 19404 10388 19460 10398
rect 19404 9714 19460 10332
rect 19516 10276 19572 10558
rect 19516 10210 19572 10220
rect 19516 10052 19572 10062
rect 19516 9958 19572 9996
rect 19404 9662 19406 9714
rect 19458 9662 19460 9714
rect 19404 9492 19460 9662
rect 19516 9716 19572 9726
rect 19628 9716 19684 10668
rect 19964 10610 20020 12124
rect 20076 12738 20132 12750
rect 20076 12686 20078 12738
rect 20130 12686 20132 12738
rect 20076 11956 20132 12686
rect 20188 12740 20244 12750
rect 20188 12646 20244 12684
rect 20532 12572 20796 12582
rect 20588 12516 20636 12572
rect 20692 12516 20740 12572
rect 20532 12506 20796 12516
rect 20860 12404 20916 12908
rect 20860 12338 20916 12348
rect 21084 12404 21140 12414
rect 20524 12290 20580 12302
rect 20524 12238 20526 12290
rect 20578 12238 20580 12290
rect 20524 12180 20580 12238
rect 20076 11890 20132 11900
rect 20412 12124 20524 12180
rect 19964 10558 19966 10610
rect 20018 10558 20020 10610
rect 19964 10546 20020 10558
rect 20188 11394 20244 11406
rect 20188 11342 20190 11394
rect 20242 11342 20244 11394
rect 20188 10052 20244 11342
rect 20412 10836 20468 12124
rect 20524 12114 20580 12124
rect 20636 12180 20692 12190
rect 20860 12180 20916 12190
rect 20636 12178 20804 12180
rect 20636 12126 20638 12178
rect 20690 12126 20804 12178
rect 20636 12124 20804 12126
rect 20636 12114 20692 12124
rect 20524 11956 20580 11966
rect 20524 11862 20580 11900
rect 20748 11956 20804 12124
rect 20748 11890 20804 11900
rect 20860 11506 20916 12124
rect 21084 11956 21140 12348
rect 21308 12292 21364 15260
rect 21420 15202 21476 15214
rect 21420 15150 21422 15202
rect 21474 15150 21476 15202
rect 21420 13860 21476 15150
rect 21532 14644 21588 15484
rect 21644 15540 21700 15550
rect 21644 15446 21700 15484
rect 21868 15540 21924 15550
rect 21868 15148 21924 15484
rect 22204 15204 22260 16046
rect 21868 15092 22036 15148
rect 22204 15138 22260 15148
rect 22316 16100 22372 16110
rect 21644 14644 21700 14654
rect 21532 14642 21700 14644
rect 21532 14590 21646 14642
rect 21698 14590 21700 14642
rect 21532 14588 21700 14590
rect 21644 14578 21700 14588
rect 21980 14306 22036 15092
rect 21980 14254 21982 14306
rect 22034 14254 22036 14306
rect 21420 13804 21924 13860
rect 21644 12852 21700 12862
rect 21644 12758 21700 12796
rect 21308 12236 21476 12292
rect 21084 11890 21140 11900
rect 21308 12068 21364 12078
rect 20860 11454 20862 11506
rect 20914 11454 20916 11506
rect 20860 11442 20916 11454
rect 20532 11004 20796 11014
rect 20588 10948 20636 11004
rect 20692 10948 20740 11004
rect 20532 10938 20796 10948
rect 20636 10836 20692 10846
rect 20412 10834 20692 10836
rect 20412 10782 20638 10834
rect 20690 10782 20692 10834
rect 20412 10780 20692 10782
rect 20188 9986 20244 9996
rect 20300 10276 20356 10286
rect 19516 9714 20132 9716
rect 19516 9662 19518 9714
rect 19570 9662 20132 9714
rect 19516 9660 20132 9662
rect 19516 9650 19572 9660
rect 19404 9436 19572 9492
rect 19292 9324 19460 9380
rect 19292 9156 19348 9166
rect 19292 9062 19348 9100
rect 19180 9044 19236 9054
rect 18956 9042 19236 9044
rect 18956 8990 19182 9042
rect 19234 8990 19236 9042
rect 18956 8988 19236 8990
rect 18844 8260 18900 8270
rect 18956 8260 19012 8988
rect 19180 8978 19236 8988
rect 19404 8820 19460 9324
rect 19516 9268 19572 9436
rect 19516 9202 19572 9212
rect 20076 9266 20132 9660
rect 20188 9604 20244 9614
rect 20300 9604 20356 10220
rect 20636 9940 20692 10780
rect 21308 10834 21364 12012
rect 21308 10782 21310 10834
rect 21362 10782 21364 10834
rect 21308 10770 21364 10782
rect 21196 10610 21252 10622
rect 21196 10558 21198 10610
rect 21250 10558 21252 10610
rect 21196 10052 21252 10558
rect 20748 9940 20804 9950
rect 20636 9938 20804 9940
rect 20636 9886 20750 9938
rect 20802 9886 20804 9938
rect 20636 9884 20804 9886
rect 20748 9874 20804 9884
rect 20188 9602 20356 9604
rect 20188 9550 20190 9602
rect 20242 9550 20356 9602
rect 20188 9548 20356 9550
rect 20188 9538 20244 9548
rect 20076 9214 20078 9266
rect 20130 9214 20132 9266
rect 20076 9202 20132 9214
rect 18844 8258 19012 8260
rect 18844 8206 18846 8258
rect 18898 8206 19012 8258
rect 18844 8204 19012 8206
rect 18844 8194 18900 8204
rect 18956 6914 19012 8204
rect 19180 8764 19460 8820
rect 19516 9042 19572 9054
rect 19516 8990 19518 9042
rect 19570 8990 19572 9042
rect 19068 8148 19124 8158
rect 19068 7474 19124 8092
rect 19180 7586 19236 8764
rect 19516 8258 19572 8990
rect 20076 8372 20132 8382
rect 20076 8278 20132 8316
rect 19516 8206 19518 8258
rect 19570 8206 19572 8258
rect 19516 8194 19572 8206
rect 20188 8148 20244 8158
rect 20188 8054 20244 8092
rect 19964 8036 20020 8046
rect 19964 7942 20020 7980
rect 20300 7588 20356 9548
rect 20532 9436 20796 9446
rect 20588 9380 20636 9436
rect 20692 9380 20740 9436
rect 20532 9370 20796 9380
rect 20524 9268 20580 9278
rect 20524 8930 20580 9212
rect 20524 8878 20526 8930
rect 20578 8878 20580 8930
rect 20524 8596 20580 8878
rect 20524 8530 20580 8540
rect 20972 8932 21028 8942
rect 20532 7868 20796 7878
rect 20588 7812 20636 7868
rect 20692 7812 20740 7868
rect 20532 7802 20796 7812
rect 19180 7534 19182 7586
rect 19234 7534 19236 7586
rect 19180 7522 19236 7534
rect 20188 7532 20356 7588
rect 19068 7422 19070 7474
rect 19122 7422 19124 7474
rect 19068 7410 19124 7422
rect 18956 6862 18958 6914
rect 19010 6862 19012 6914
rect 18956 6850 19012 6862
rect 19068 6692 19124 6702
rect 19964 6692 20020 6702
rect 19068 6690 20020 6692
rect 19068 6638 19070 6690
rect 19122 6638 19966 6690
rect 20018 6638 20020 6690
rect 19068 6636 20020 6638
rect 19068 6626 19124 6636
rect 19516 6020 19572 6030
rect 18732 5740 19012 5796
rect 18844 5572 18900 5582
rect 18844 5348 18900 5516
rect 18508 5068 18676 5124
rect 18732 5124 18788 5134
rect 18508 5012 18564 5068
rect 18508 4918 18564 4956
rect 18620 4900 18676 4910
rect 18732 4900 18788 5068
rect 18844 5122 18900 5292
rect 18844 5070 18846 5122
rect 18898 5070 18900 5122
rect 18844 5058 18900 5070
rect 18620 4898 18788 4900
rect 18620 4846 18622 4898
rect 18674 4846 18788 4898
rect 18620 4844 18788 4846
rect 18620 4834 18676 4844
rect 18956 4788 19012 5740
rect 18956 4452 19012 4732
rect 18620 4396 19012 4452
rect 19068 5794 19124 5806
rect 19068 5742 19070 5794
rect 19122 5742 19124 5794
rect 19068 5012 19124 5742
rect 19516 5794 19572 5964
rect 19516 5742 19518 5794
rect 19570 5742 19572 5794
rect 19180 5124 19236 5134
rect 19180 5030 19236 5068
rect 18396 3602 18452 3612
rect 18508 3668 18564 3678
rect 18620 3668 18676 4396
rect 18956 4228 19012 4238
rect 19068 4228 19124 4956
rect 18956 4226 19124 4228
rect 18956 4174 18958 4226
rect 19010 4174 19124 4226
rect 18956 4172 19124 4174
rect 18956 4162 19012 4172
rect 18508 3666 18676 3668
rect 18508 3614 18510 3666
rect 18562 3614 18676 3666
rect 18508 3612 18676 3614
rect 18508 3602 18564 3612
rect 17948 3556 18004 3566
rect 17948 3462 18004 3500
rect 18844 3556 18900 3566
rect 18844 3462 18900 3500
rect 19068 2772 19124 4172
rect 19516 3892 19572 5742
rect 19740 5012 19796 6636
rect 19964 6626 20020 6636
rect 19964 5794 20020 5806
rect 19964 5742 19966 5794
rect 20018 5742 20020 5794
rect 19964 5236 20020 5742
rect 19964 5170 20020 5180
rect 19740 4946 19796 4956
rect 19852 4898 19908 4910
rect 19852 4846 19854 4898
rect 19906 4846 19908 4898
rect 19740 4564 19796 4574
rect 19740 4004 19796 4508
rect 19852 4116 19908 4846
rect 19964 4900 20020 4910
rect 19964 4806 20020 4844
rect 20076 4898 20132 4910
rect 20076 4846 20078 4898
rect 20130 4846 20132 4898
rect 20076 4564 20132 4846
rect 20076 4498 20132 4508
rect 20076 4116 20132 4126
rect 19852 4114 20132 4116
rect 19852 4062 20078 4114
rect 20130 4062 20132 4114
rect 19852 4060 20132 4062
rect 19740 3948 19908 4004
rect 19516 3826 19572 3836
rect 19068 2706 19124 2716
rect 19740 3556 19796 3566
rect 19740 800 19796 3500
rect 19852 3554 19908 3948
rect 20076 3666 20132 4060
rect 20188 4004 20244 7532
rect 20412 7364 20468 7374
rect 20412 4564 20468 7308
rect 20972 6356 21028 8876
rect 21196 8484 21252 9996
rect 21420 8596 21476 12236
rect 21532 12068 21588 12078
rect 21532 11974 21588 12012
rect 21644 11508 21700 11518
rect 21644 11414 21700 11452
rect 21868 11506 21924 13804
rect 21980 12404 22036 14254
rect 22092 12852 22148 12862
rect 22092 12758 22148 12796
rect 21980 12338 22036 12348
rect 22204 12404 22260 12414
rect 22204 12290 22260 12348
rect 22204 12238 22206 12290
rect 22258 12238 22260 12290
rect 22204 12226 22260 12238
rect 22316 12290 22372 16044
rect 22652 16100 22708 16110
rect 22652 16006 22708 16044
rect 22876 15540 22932 16718
rect 23772 16770 23828 16782
rect 23772 16718 23774 16770
rect 23826 16718 23828 16770
rect 23436 16212 23492 16222
rect 22876 15474 22932 15484
rect 23324 16100 23380 16110
rect 23324 15874 23380 16044
rect 23324 15822 23326 15874
rect 23378 15822 23380 15874
rect 23324 15428 23380 15822
rect 23436 15652 23492 16156
rect 23772 16100 23828 16718
rect 23772 16034 23828 16044
rect 24220 16100 24276 16110
rect 24220 16006 24276 16044
rect 24332 15876 24388 16830
rect 24668 16882 24724 16894
rect 24668 16830 24670 16882
rect 24722 16830 24724 16882
rect 24668 16100 24724 16830
rect 24780 16884 24836 16894
rect 24780 16790 24836 16828
rect 24892 16882 24948 16894
rect 24892 16830 24894 16882
rect 24946 16830 24948 16882
rect 24892 16324 24948 16830
rect 24668 16034 24724 16044
rect 24780 16268 24948 16324
rect 24780 16098 24836 16268
rect 24780 16046 24782 16098
rect 24834 16046 24836 16098
rect 23436 15586 23492 15596
rect 24220 15820 24388 15876
rect 23324 15362 23380 15372
rect 22876 15316 22932 15326
rect 22428 15204 22484 15242
rect 22876 15222 22932 15260
rect 23996 15314 24052 15326
rect 23996 15262 23998 15314
rect 24050 15262 24052 15314
rect 22428 14644 22484 15148
rect 23884 15202 23940 15214
rect 23884 15150 23886 15202
rect 23938 15150 23940 15202
rect 22540 14644 22596 14654
rect 22428 14642 22596 14644
rect 22428 14590 22542 14642
rect 22594 14590 22596 14642
rect 22428 14588 22596 14590
rect 22540 14578 22596 14588
rect 23884 14418 23940 15150
rect 23884 14366 23886 14418
rect 23938 14366 23940 14418
rect 23100 13860 23156 13870
rect 23100 13766 23156 13804
rect 23884 13860 23940 14366
rect 23996 14306 24052 15262
rect 24220 14530 24276 15820
rect 24556 15428 24612 15438
rect 24780 15428 24836 16046
rect 24892 16100 24948 16110
rect 25004 16100 25060 18060
rect 24892 16098 25060 16100
rect 24892 16046 24894 16098
rect 24946 16046 25060 16098
rect 24892 16044 25060 16046
rect 24892 16034 24948 16044
rect 24556 15426 24836 15428
rect 24556 15374 24558 15426
rect 24610 15374 24836 15426
rect 24556 15372 24836 15374
rect 24556 15362 24612 15372
rect 24668 14868 24724 14878
rect 24668 14642 24724 14812
rect 24668 14590 24670 14642
rect 24722 14590 24724 14642
rect 24668 14578 24724 14590
rect 24220 14478 24222 14530
rect 24274 14478 24276 14530
rect 24220 14466 24276 14478
rect 23996 14254 23998 14306
rect 24050 14254 24052 14306
rect 23996 13972 24052 14254
rect 23996 13906 24052 13916
rect 23884 13794 23940 13804
rect 24780 13858 24836 13870
rect 24780 13806 24782 13858
rect 24834 13806 24836 13858
rect 22540 13746 22596 13758
rect 22540 13694 22542 13746
rect 22594 13694 22596 13746
rect 22540 12404 22596 13694
rect 24668 13746 24724 13758
rect 24668 13694 24670 13746
rect 24722 13694 24724 13746
rect 24556 13300 24612 13310
rect 22316 12238 22318 12290
rect 22370 12238 22372 12290
rect 22316 12068 22372 12238
rect 21868 11454 21870 11506
rect 21922 11454 21924 11506
rect 21868 11442 21924 11454
rect 21980 12012 22372 12068
rect 22428 12402 22596 12404
rect 22428 12350 22542 12402
rect 22594 12350 22596 12402
rect 22428 12348 22596 12350
rect 21980 11732 22036 12012
rect 22428 11844 22484 12348
rect 22540 12338 22596 12348
rect 22988 12964 23044 12974
rect 21532 10724 21588 10734
rect 21532 10630 21588 10668
rect 21644 10052 21700 10062
rect 21644 9938 21700 9996
rect 21644 9886 21646 9938
rect 21698 9886 21700 9938
rect 21644 9874 21700 9886
rect 21644 9268 21700 9278
rect 21644 9174 21700 9212
rect 21980 9044 22036 11676
rect 22092 11788 22484 11844
rect 22876 12066 22932 12078
rect 22876 12014 22878 12066
rect 22930 12014 22932 12066
rect 22092 11394 22148 11788
rect 22876 11732 22932 12014
rect 22876 11666 22932 11676
rect 22092 11342 22094 11394
rect 22146 11342 22148 11394
rect 22092 11330 22148 11342
rect 22204 11396 22260 11406
rect 22204 11302 22260 11340
rect 22316 11170 22372 11182
rect 22316 11118 22318 11170
rect 22370 11118 22372 11170
rect 22316 10724 22372 11118
rect 22316 10610 22372 10668
rect 22316 10558 22318 10610
rect 22370 10558 22372 10610
rect 22316 10546 22372 10558
rect 22092 10498 22148 10510
rect 22092 10446 22094 10498
rect 22146 10446 22148 10498
rect 22092 9940 22148 10446
rect 22092 9874 22148 9884
rect 22316 9940 22372 9950
rect 22092 9044 22148 9054
rect 21980 9042 22148 9044
rect 21980 8990 22094 9042
rect 22146 8990 22148 9042
rect 21980 8988 22148 8990
rect 22092 8978 22148 8988
rect 22316 9044 22372 9884
rect 22988 9940 23044 12908
rect 23324 12404 23380 12414
rect 23324 12310 23380 12348
rect 24332 11508 24388 11518
rect 24332 10722 24388 11452
rect 24332 10670 24334 10722
rect 24386 10670 24388 10722
rect 24332 10658 24388 10670
rect 22876 9828 22932 9838
rect 22988 9828 23044 9884
rect 22876 9826 23044 9828
rect 22876 9774 22878 9826
rect 22930 9774 23044 9826
rect 22876 9772 23044 9774
rect 23548 10610 23604 10622
rect 23548 10558 23550 10610
rect 23602 10558 23604 10610
rect 22876 9762 22932 9772
rect 22652 9604 22708 9614
rect 22652 9268 22708 9548
rect 22988 9604 23044 9614
rect 22988 9510 23044 9548
rect 23212 9604 23268 9614
rect 23548 9604 23604 10558
rect 23212 9602 23604 9604
rect 23212 9550 23214 9602
rect 23266 9550 23604 9602
rect 23212 9548 23604 9550
rect 23660 9714 23716 9726
rect 23660 9662 23662 9714
rect 23714 9662 23716 9714
rect 23212 9538 23268 9548
rect 22652 9136 22708 9212
rect 22316 8978 22372 8988
rect 21420 8530 21476 8540
rect 21196 8418 21252 8428
rect 22652 8260 22708 8270
rect 21644 8036 21700 8046
rect 21644 7588 21700 7980
rect 22204 8034 22260 8046
rect 22204 7982 22206 8034
rect 22258 7982 22260 8034
rect 22204 7700 22260 7982
rect 22428 8036 22484 8046
rect 22428 7942 22484 7980
rect 22540 8034 22596 8046
rect 22540 7982 22542 8034
rect 22594 7982 22596 8034
rect 22540 7924 22596 7982
rect 22540 7858 22596 7868
rect 22204 7634 22260 7644
rect 21644 7522 21700 7532
rect 22092 7588 22148 7598
rect 20532 6300 20796 6310
rect 20588 6244 20636 6300
rect 20692 6244 20740 6300
rect 20972 6290 21028 6300
rect 21980 6690 22036 6702
rect 21980 6638 21982 6690
rect 22034 6638 22036 6690
rect 20532 6234 20796 6244
rect 21756 6018 21812 6030
rect 21756 5966 21758 6018
rect 21810 5966 21812 6018
rect 20524 5124 20580 5134
rect 20524 5122 21140 5124
rect 20524 5070 20526 5122
rect 20578 5070 21140 5122
rect 20524 5068 21140 5070
rect 20524 5058 20580 5068
rect 20972 4898 21028 4910
rect 20972 4846 20974 4898
rect 21026 4846 21028 4898
rect 20532 4732 20796 4742
rect 20588 4676 20636 4732
rect 20692 4676 20740 4732
rect 20532 4666 20796 4676
rect 20412 4508 20580 4564
rect 20300 4340 20356 4350
rect 20300 4226 20356 4284
rect 20300 4174 20302 4226
rect 20354 4174 20356 4226
rect 20300 4162 20356 4174
rect 20412 4338 20468 4350
rect 20412 4286 20414 4338
rect 20466 4286 20468 4338
rect 20412 4228 20468 4286
rect 20412 4162 20468 4172
rect 20188 3938 20244 3948
rect 20076 3614 20078 3666
rect 20130 3614 20132 3666
rect 20076 3602 20132 3614
rect 20524 3666 20580 4508
rect 20524 3614 20526 3666
rect 20578 3614 20580 3666
rect 20524 3602 20580 3614
rect 19852 3502 19854 3554
rect 19906 3502 19908 3554
rect 19852 3490 19908 3502
rect 20972 3556 21028 4846
rect 21084 4562 21140 5068
rect 21084 4510 21086 4562
rect 21138 4510 21140 4562
rect 21084 4498 21140 4510
rect 21308 4450 21364 4462
rect 21308 4398 21310 4450
rect 21362 4398 21364 4450
rect 21308 4228 21364 4398
rect 21308 4162 21364 4172
rect 21420 4340 21476 4350
rect 20972 3490 21028 3500
rect 21420 3220 21476 4284
rect 21756 4116 21812 5966
rect 21980 5906 22036 6638
rect 22092 6130 22148 7532
rect 22316 7364 22372 7374
rect 22316 7270 22372 7308
rect 22652 7250 22708 8204
rect 22764 7588 22820 7598
rect 22764 7474 22820 7532
rect 22764 7422 22766 7474
rect 22818 7422 22820 7474
rect 22764 7410 22820 7422
rect 22652 7198 22654 7250
rect 22706 7198 22708 7250
rect 22652 7186 22708 7198
rect 22092 6078 22094 6130
rect 22146 6078 22148 6130
rect 22092 6066 22148 6078
rect 22204 6802 22260 6814
rect 22204 6750 22206 6802
rect 22258 6750 22260 6802
rect 21980 5854 21982 5906
rect 22034 5854 22036 5906
rect 21980 5796 22036 5854
rect 21980 5730 22036 5740
rect 22204 5906 22260 6750
rect 22652 6692 22708 6702
rect 22652 6598 22708 6636
rect 23212 6468 23268 6478
rect 23100 6466 23268 6468
rect 23100 6414 23214 6466
rect 23266 6414 23268 6466
rect 23100 6412 23268 6414
rect 22204 5854 22206 5906
rect 22258 5854 22260 5906
rect 22204 5346 22260 5854
rect 22876 5908 22932 5918
rect 22876 5814 22932 5852
rect 22204 5294 22206 5346
rect 22258 5294 22260 5346
rect 22204 5282 22260 5294
rect 22540 5796 22596 5806
rect 21980 5236 22036 5246
rect 21980 4450 22036 5180
rect 22540 5124 22596 5740
rect 22092 5122 22596 5124
rect 22092 5070 22542 5122
rect 22594 5070 22596 5122
rect 22092 5068 22596 5070
rect 22092 4562 22148 5068
rect 22540 5058 22596 5068
rect 22092 4510 22094 4562
rect 22146 4510 22148 4562
rect 22092 4498 22148 4510
rect 21980 4398 21982 4450
rect 22034 4398 22036 4450
rect 21980 4386 22036 4398
rect 23100 4452 23156 6412
rect 23212 6402 23268 6412
rect 23212 6244 23268 6254
rect 23212 5906 23268 6188
rect 23324 6130 23380 9548
rect 23548 9380 23604 9390
rect 23548 9042 23604 9324
rect 23548 8990 23550 9042
rect 23602 8990 23604 9042
rect 23548 8484 23604 8990
rect 23660 8932 23716 9662
rect 23772 9602 23828 9614
rect 23772 9550 23774 9602
rect 23826 9550 23828 9602
rect 23772 9380 23828 9550
rect 23772 9314 23828 9324
rect 23996 9602 24052 9614
rect 23996 9550 23998 9602
rect 24050 9550 24052 9602
rect 23996 9268 24052 9550
rect 23996 9202 24052 9212
rect 24444 9604 24500 9614
rect 24332 9156 24388 9166
rect 24332 9062 24388 9100
rect 23772 8932 23828 8942
rect 23660 8930 23828 8932
rect 23660 8878 23774 8930
rect 23826 8878 23828 8930
rect 23660 8876 23828 8878
rect 23548 8418 23604 8428
rect 23436 8370 23492 8382
rect 23436 8318 23438 8370
rect 23490 8318 23492 8370
rect 23436 8260 23492 8318
rect 23436 8194 23492 8204
rect 23548 8258 23604 8270
rect 23548 8206 23550 8258
rect 23602 8206 23604 8258
rect 23548 8036 23604 8206
rect 23548 7970 23604 7980
rect 23660 7700 23716 7710
rect 23660 7606 23716 7644
rect 23772 7476 23828 8876
rect 24220 8372 24276 8382
rect 24220 8278 24276 8316
rect 23884 7588 23940 7598
rect 23884 7494 23940 7532
rect 23548 7420 23828 7476
rect 23996 7474 24052 7486
rect 23996 7422 23998 7474
rect 24050 7422 24052 7474
rect 23548 6692 23604 7420
rect 23996 7364 24052 7422
rect 23996 7298 24052 7308
rect 24220 7364 24276 7374
rect 23996 6692 24052 6702
rect 23548 6626 23604 6636
rect 23660 6690 24052 6692
rect 23660 6638 23998 6690
rect 24050 6638 24052 6690
rect 23660 6636 24052 6638
rect 23660 6244 23716 6636
rect 23996 6626 24052 6636
rect 24108 6580 24164 6590
rect 24108 6486 24164 6524
rect 23772 6466 23828 6478
rect 23772 6414 23774 6466
rect 23826 6414 23828 6466
rect 23772 6356 23828 6414
rect 23884 6466 23940 6478
rect 23884 6414 23886 6466
rect 23938 6414 23940 6466
rect 23884 6356 23940 6414
rect 23884 6300 24164 6356
rect 23772 6290 23828 6300
rect 23660 6178 23716 6188
rect 23324 6078 23326 6130
rect 23378 6078 23380 6130
rect 23324 6066 23380 6078
rect 23212 5854 23214 5906
rect 23266 5854 23268 5906
rect 23212 5842 23268 5854
rect 23548 5908 23604 5918
rect 23548 5906 23940 5908
rect 23548 5854 23550 5906
rect 23602 5854 23940 5906
rect 23548 5852 23940 5854
rect 23548 5842 23604 5852
rect 23436 5796 23492 5806
rect 23436 5702 23492 5740
rect 23884 5122 23940 5852
rect 23884 5070 23886 5122
rect 23938 5070 23940 5122
rect 23436 5012 23492 5022
rect 23436 4562 23492 4956
rect 23436 4510 23438 4562
rect 23490 4510 23492 4562
rect 23436 4498 23492 4510
rect 23772 4564 23828 4574
rect 23884 4564 23940 5070
rect 23772 4562 23940 4564
rect 23772 4510 23774 4562
rect 23826 4510 23940 4562
rect 23772 4508 23940 4510
rect 23996 4788 24052 4798
rect 24108 4788 24164 6300
rect 24052 4732 24164 4788
rect 23772 4498 23828 4508
rect 23100 4386 23156 4396
rect 23996 4450 24052 4732
rect 23996 4398 23998 4450
rect 24050 4398 24052 4450
rect 22876 4226 22932 4238
rect 22876 4174 22878 4226
rect 22930 4174 22932 4226
rect 22092 4116 22148 4126
rect 21756 4114 22148 4116
rect 21756 4062 22094 4114
rect 22146 4062 22148 4114
rect 21756 4060 22148 4062
rect 22092 4050 22148 4060
rect 21644 4004 21700 4014
rect 21644 3666 21700 3948
rect 22876 3892 22932 4174
rect 23996 4004 24052 4398
rect 24108 4452 24164 4462
rect 24108 4116 24164 4396
rect 24108 4050 24164 4060
rect 23996 3938 24052 3948
rect 22876 3826 22932 3836
rect 21644 3614 21646 3666
rect 21698 3614 21700 3666
rect 21644 3602 21700 3614
rect 22652 3668 22708 3678
rect 22652 3574 22708 3612
rect 24108 3666 24164 3678
rect 24108 3614 24110 3666
rect 24162 3614 24164 3666
rect 20532 3164 20796 3174
rect 20588 3108 20636 3164
rect 20692 3108 20740 3164
rect 21420 3154 21476 3164
rect 21868 3556 21924 3566
rect 20532 3098 20796 3108
rect 21868 800 21924 3500
rect 22092 3556 22148 3566
rect 22092 3462 22148 3500
rect 23548 3444 23604 3482
rect 23548 3378 23604 3388
rect 24108 3388 24164 3614
rect 24220 3388 24276 7308
rect 24332 6692 24388 6702
rect 24444 6692 24500 9548
rect 24388 6636 24500 6692
rect 24332 6598 24388 6636
rect 24444 6356 24500 6366
rect 24444 5908 24500 6300
rect 24444 5814 24500 5852
rect 24556 5348 24612 13244
rect 24668 12180 24724 13694
rect 24780 12964 24836 13806
rect 25004 13748 25060 13758
rect 25004 13654 25060 13692
rect 25004 12964 25060 12974
rect 24780 12962 25060 12964
rect 24780 12910 25006 12962
rect 25058 12910 25060 12962
rect 24780 12908 25060 12910
rect 25004 12740 25060 12908
rect 25004 12674 25060 12684
rect 24668 12114 24724 12124
rect 24892 12066 24948 12078
rect 24892 12014 24894 12066
rect 24946 12014 24948 12066
rect 24892 11844 24948 12014
rect 24892 11778 24948 11788
rect 25004 11508 25060 11518
rect 25004 11414 25060 11452
rect 24892 11396 24948 11406
rect 24892 11302 24948 11340
rect 25116 10164 25172 20524
rect 25788 20244 25844 20972
rect 25900 20914 25956 21532
rect 26124 21588 26180 21598
rect 26124 21494 26180 21532
rect 26572 21588 26628 22876
rect 26684 22708 26740 22718
rect 26684 22370 26740 22652
rect 26684 22318 26686 22370
rect 26738 22318 26740 22370
rect 26684 22306 26740 22318
rect 25900 20862 25902 20914
rect 25954 20862 25956 20914
rect 25900 20850 25956 20862
rect 26012 21474 26068 21486
rect 26012 21422 26014 21474
rect 26066 21422 26068 21474
rect 26012 20916 26068 21422
rect 26572 21026 26628 21532
rect 26572 20974 26574 21026
rect 26626 20974 26628 21026
rect 26572 20962 26628 20974
rect 26796 22260 26852 22270
rect 26796 21474 26852 22204
rect 27132 22148 27188 25340
rect 27580 24946 27636 25452
rect 27580 24894 27582 24946
rect 27634 24894 27636 24946
rect 27580 24882 27636 24894
rect 27692 24948 27748 24958
rect 27804 24948 27860 27020
rect 28028 26964 28084 27806
rect 28140 27970 28196 28476
rect 28140 27918 28142 27970
rect 28194 27918 28196 27970
rect 28140 27188 28196 27918
rect 28364 27300 28420 27310
rect 28364 27206 28420 27244
rect 28252 27188 28308 27198
rect 28140 27186 28308 27188
rect 28140 27134 28254 27186
rect 28306 27134 28308 27186
rect 28140 27132 28308 27134
rect 28252 27122 28308 27132
rect 28252 26964 28308 26974
rect 28028 26908 28252 26964
rect 27916 26852 27972 26862
rect 27916 25508 27972 26796
rect 28028 25620 28084 25630
rect 28028 25526 28084 25564
rect 27916 25376 27972 25452
rect 27692 24946 27860 24948
rect 27692 24894 27694 24946
rect 27746 24894 27860 24946
rect 27692 24892 27860 24894
rect 28140 25282 28196 25294
rect 28140 25230 28142 25282
rect 28194 25230 28196 25282
rect 27692 24882 27748 24892
rect 27804 24500 27860 24510
rect 28140 24500 28196 25230
rect 27804 24498 28196 24500
rect 27804 24446 27806 24498
rect 27858 24446 28196 24498
rect 27804 24444 28196 24446
rect 28252 24610 28308 26908
rect 28364 26404 28420 26414
rect 28476 26404 28532 28588
rect 28588 28308 28644 28812
rect 28812 28866 28868 29372
rect 29372 29316 29428 30156
rect 28812 28814 28814 28866
rect 28866 28814 28868 28866
rect 28812 28802 28868 28814
rect 29260 29314 29428 29316
rect 29260 29262 29374 29314
rect 29426 29262 29428 29314
rect 29260 29260 29428 29262
rect 28700 28532 28756 28542
rect 28700 28438 28756 28476
rect 28588 28252 28756 28308
rect 28700 28082 28756 28252
rect 28700 28030 28702 28082
rect 28754 28030 28756 28082
rect 28700 28018 28756 28030
rect 28588 27972 28644 27982
rect 28588 27878 28644 27916
rect 28924 27858 28980 27870
rect 28924 27806 28926 27858
rect 28978 27806 28980 27858
rect 28364 26402 28532 26404
rect 28364 26350 28366 26402
rect 28418 26350 28532 26402
rect 28364 26348 28532 26350
rect 28700 27748 28756 27758
rect 28364 26338 28420 26348
rect 28252 24558 28254 24610
rect 28306 24558 28308 24610
rect 27244 24052 27300 24062
rect 27244 23958 27300 23996
rect 27468 23938 27524 23950
rect 27468 23886 27470 23938
rect 27522 23886 27524 23938
rect 27356 23492 27412 23502
rect 27356 22932 27412 23436
rect 27468 23044 27524 23886
rect 27804 23268 27860 24444
rect 28252 24052 28308 24558
rect 27916 23828 27972 23838
rect 27916 23734 27972 23772
rect 28252 23828 28308 23996
rect 28252 23762 28308 23772
rect 28252 23268 28308 23278
rect 27804 23266 28308 23268
rect 27804 23214 28254 23266
rect 28306 23214 28308 23266
rect 27804 23212 28308 23214
rect 27804 23044 27860 23054
rect 27468 23042 27860 23044
rect 27468 22990 27806 23042
rect 27858 22990 27860 23042
rect 27468 22988 27860 22990
rect 27356 22876 27636 22932
rect 27132 22082 27188 22092
rect 27356 22146 27412 22158
rect 27356 22094 27358 22146
rect 27410 22094 27412 22146
rect 26796 21422 26798 21474
rect 26850 21422 26852 21474
rect 26012 20850 26068 20860
rect 26460 20692 26516 20702
rect 25788 20132 25844 20188
rect 26124 20468 26180 20478
rect 25900 20132 25956 20142
rect 25788 20130 25956 20132
rect 25788 20078 25902 20130
rect 25954 20078 25956 20130
rect 25788 20076 25956 20078
rect 25900 20066 25956 20076
rect 25900 19572 25956 19582
rect 25676 18564 25732 18574
rect 25676 18470 25732 18508
rect 25900 18452 25956 19516
rect 25900 18386 25956 18396
rect 26012 18900 26068 18910
rect 25228 17668 25284 17678
rect 25228 13300 25284 17612
rect 25788 17444 25844 17454
rect 25900 17444 25956 17454
rect 25788 17442 25900 17444
rect 25788 17390 25790 17442
rect 25842 17390 25900 17442
rect 25788 17388 25900 17390
rect 25788 17378 25844 17388
rect 25788 16884 25844 16894
rect 25788 16770 25844 16828
rect 25788 16718 25790 16770
rect 25842 16718 25844 16770
rect 25788 16706 25844 16718
rect 25900 16882 25956 17388
rect 25900 16830 25902 16882
rect 25954 16830 25956 16882
rect 25452 15876 25508 15886
rect 25900 15876 25956 16830
rect 25340 15874 25956 15876
rect 25340 15822 25454 15874
rect 25506 15822 25956 15874
rect 25340 15820 25956 15822
rect 25340 13412 25396 15820
rect 25452 15810 25508 15820
rect 26012 15148 26068 18844
rect 26124 18340 26180 20412
rect 26460 20356 26516 20636
rect 26572 20580 26628 20590
rect 26572 20486 26628 20524
rect 26460 20290 26516 20300
rect 26348 19906 26404 19918
rect 26348 19854 26350 19906
rect 26402 19854 26404 19906
rect 26348 19572 26404 19854
rect 26348 19506 26404 19516
rect 26236 19460 26292 19470
rect 26236 19366 26292 19404
rect 26348 19236 26404 19246
rect 26348 19142 26404 19180
rect 26236 19124 26292 19134
rect 26796 19124 26852 21422
rect 27356 21476 27412 22094
rect 27580 22146 27636 22876
rect 27580 22094 27582 22146
rect 27634 22094 27636 22146
rect 27580 22036 27636 22094
rect 27692 22258 27748 22270
rect 27692 22206 27694 22258
rect 27746 22206 27748 22258
rect 27692 22148 27748 22206
rect 27692 22082 27748 22092
rect 27580 21970 27636 21980
rect 27580 21588 27636 21598
rect 27580 21494 27636 21532
rect 27468 21476 27524 21486
rect 27356 21474 27524 21476
rect 27356 21422 27470 21474
rect 27522 21422 27524 21474
rect 27356 21420 27524 21422
rect 27244 21028 27300 21038
rect 27356 21028 27412 21420
rect 27468 21410 27524 21420
rect 27804 21364 27860 22988
rect 27244 21026 27412 21028
rect 27244 20974 27246 21026
rect 27298 20974 27412 21026
rect 27244 20972 27412 20974
rect 27580 21308 27860 21364
rect 27916 22708 27972 22718
rect 27244 20962 27300 20972
rect 27468 20916 27524 20926
rect 27468 20822 27524 20860
rect 27580 20692 27636 21308
rect 27916 21252 27972 22652
rect 28140 22148 28196 22158
rect 28140 22054 28196 22092
rect 27692 21196 27972 21252
rect 27692 20802 27748 21196
rect 27692 20750 27694 20802
rect 27746 20750 27748 20802
rect 27692 20738 27748 20750
rect 28252 20804 28308 23212
rect 28588 22146 28644 22158
rect 28588 22094 28590 22146
rect 28642 22094 28644 22146
rect 28588 22036 28644 22094
rect 28588 21970 28644 21980
rect 28476 20804 28532 20814
rect 28700 20804 28756 27692
rect 28812 26964 28868 26974
rect 28812 26870 28868 26908
rect 28924 26852 28980 27806
rect 29036 27858 29092 27870
rect 29036 27806 29038 27858
rect 29090 27806 29092 27858
rect 29036 27300 29092 27806
rect 29036 27234 29092 27244
rect 28924 26786 28980 26796
rect 29148 23154 29204 23166
rect 29148 23102 29150 23154
rect 29202 23102 29204 23154
rect 29148 22708 29204 23102
rect 29148 22642 29204 22652
rect 28252 20802 28532 20804
rect 28252 20750 28478 20802
rect 28530 20750 28532 20802
rect 28252 20748 28532 20750
rect 28476 20738 28532 20748
rect 28588 20748 28756 20804
rect 29148 21586 29204 21598
rect 29148 21534 29150 21586
rect 29202 21534 29204 21586
rect 27356 20636 27636 20692
rect 27244 20244 27300 20254
rect 27356 20244 27412 20636
rect 27804 20580 27860 20590
rect 27804 20486 27860 20524
rect 27916 20578 27972 20590
rect 27916 20526 27918 20578
rect 27970 20526 27972 20578
rect 27244 20242 27412 20244
rect 27244 20190 27246 20242
rect 27298 20190 27412 20242
rect 27244 20188 27412 20190
rect 27468 20468 27524 20478
rect 27468 20244 27524 20412
rect 27244 20178 27300 20188
rect 27468 20178 27524 20188
rect 27804 20244 27860 20254
rect 27580 20020 27636 20030
rect 27580 20018 27748 20020
rect 27580 19966 27582 20018
rect 27634 19966 27748 20018
rect 27580 19964 27748 19966
rect 27580 19954 27636 19964
rect 26908 19908 26964 19918
rect 26908 19814 26964 19852
rect 27692 19908 27748 19964
rect 26908 19124 26964 19134
rect 26796 19068 26908 19124
rect 26236 19030 26292 19068
rect 26908 19030 26964 19068
rect 27468 19124 27524 19134
rect 26684 18452 26740 18462
rect 26684 18358 26740 18396
rect 27132 18452 27188 18462
rect 27132 18358 27188 18396
rect 26236 18340 26292 18350
rect 26124 18338 26292 18340
rect 26124 18286 26238 18338
rect 26290 18286 26292 18338
rect 26124 18284 26292 18286
rect 26236 18228 26292 18284
rect 26236 18172 26628 18228
rect 26348 17556 26404 17566
rect 26348 17462 26404 17500
rect 26236 17442 26292 17454
rect 26236 17390 26238 17442
rect 26290 17390 26292 17442
rect 26124 16884 26180 16894
rect 26124 16098 26180 16828
rect 26236 16210 26292 17390
rect 26460 17444 26516 17454
rect 26460 17350 26516 17388
rect 26572 17332 26628 18172
rect 26572 17266 26628 17276
rect 26796 17666 26852 17678
rect 26796 17614 26798 17666
rect 26850 17614 26852 17666
rect 26236 16158 26238 16210
rect 26290 16158 26292 16210
rect 26236 16146 26292 16158
rect 26124 16046 26126 16098
rect 26178 16046 26180 16098
rect 26124 15988 26180 16046
rect 26124 15922 26180 15932
rect 26460 16100 26516 16110
rect 26796 16100 26852 17614
rect 27468 17444 27524 19068
rect 27580 19010 27636 19022
rect 27580 18958 27582 19010
rect 27634 18958 27636 19010
rect 27580 18452 27636 18958
rect 27580 18386 27636 18396
rect 27692 18450 27748 19852
rect 27804 19234 27860 20188
rect 27916 19796 27972 20526
rect 28364 20356 28420 20366
rect 28252 20132 28308 20142
rect 27916 19730 27972 19740
rect 28140 20130 28308 20132
rect 28140 20078 28254 20130
rect 28306 20078 28308 20130
rect 28140 20076 28308 20078
rect 27804 19182 27806 19234
rect 27858 19182 27860 19234
rect 27804 19170 27860 19182
rect 28140 18676 28196 20076
rect 28252 20066 28308 20076
rect 28364 20018 28420 20300
rect 28588 20188 28644 20748
rect 28812 20690 28868 20702
rect 28812 20638 28814 20690
rect 28866 20638 28868 20690
rect 28364 19966 28366 20018
rect 28418 19966 28420 20018
rect 28252 19796 28308 19806
rect 28252 19702 28308 19740
rect 28252 19010 28308 19022
rect 28252 18958 28254 19010
rect 28306 18958 28308 19010
rect 28252 18900 28308 18958
rect 28252 18834 28308 18844
rect 27916 18620 28196 18676
rect 27692 18398 27694 18450
rect 27746 18398 27748 18450
rect 27692 17444 27748 18398
rect 27804 18564 27860 18574
rect 27916 18564 27972 18620
rect 27804 18562 27972 18564
rect 27804 18510 27806 18562
rect 27858 18510 27972 18562
rect 27804 18508 27972 18510
rect 27804 18452 27860 18508
rect 27804 18386 27860 18396
rect 28028 18452 28084 18462
rect 28028 18358 28084 18396
rect 28364 18340 28420 19966
rect 28364 18274 28420 18284
rect 28476 20132 28644 20188
rect 28700 20578 28756 20590
rect 28700 20526 28702 20578
rect 28754 20526 28756 20578
rect 28140 17444 28196 17454
rect 27692 17442 28196 17444
rect 27692 17390 28142 17442
rect 28194 17390 28196 17442
rect 27692 17388 28196 17390
rect 27244 16882 27300 16894
rect 27244 16830 27246 16882
rect 27298 16830 27300 16882
rect 26908 16100 26964 16110
rect 26796 16098 26964 16100
rect 26796 16046 26910 16098
rect 26962 16046 26964 16098
rect 26796 16044 26964 16046
rect 26460 15986 26516 16044
rect 26908 16034 26964 16044
rect 27244 16100 27300 16830
rect 27468 16436 27524 17388
rect 28028 16996 28084 17388
rect 28140 17378 28196 17388
rect 28476 17220 28532 20132
rect 28700 19348 28756 20526
rect 28812 20356 28868 20638
rect 28812 20290 28868 20300
rect 29036 20692 29092 20702
rect 29036 20188 29092 20636
rect 28700 18900 28756 19292
rect 28812 20132 29092 20188
rect 29148 20244 29204 21534
rect 29148 20178 29204 20188
rect 28812 19346 28868 20132
rect 29036 19908 29092 19918
rect 29036 19814 29092 19852
rect 28812 19294 28814 19346
rect 28866 19294 28868 19346
rect 28812 19282 28868 19294
rect 28700 18834 28756 18844
rect 28028 16930 28084 16940
rect 28140 17164 28532 17220
rect 28588 18340 28644 18350
rect 28028 16772 28084 16782
rect 28028 16678 28084 16716
rect 27468 16380 27860 16436
rect 27244 16006 27300 16044
rect 26460 15934 26462 15986
rect 26514 15934 26516 15986
rect 26460 15148 26516 15934
rect 27132 15988 27188 15998
rect 27132 15894 27188 15932
rect 25788 15092 26068 15148
rect 26124 15092 26516 15148
rect 27468 15202 27524 15214
rect 27468 15150 27470 15202
rect 27522 15150 27524 15202
rect 25452 14868 25508 14878
rect 25452 14530 25508 14812
rect 25452 14478 25454 14530
rect 25506 14478 25508 14530
rect 25452 13860 25508 14478
rect 25452 13794 25508 13804
rect 25564 13748 25620 13758
rect 25564 13654 25620 13692
rect 25452 13412 25508 13422
rect 25340 13356 25452 13412
rect 25452 13346 25508 13356
rect 25228 13244 25396 13300
rect 25228 13074 25284 13086
rect 25228 13022 25230 13074
rect 25282 13022 25284 13074
rect 25228 12180 25284 13022
rect 25228 12114 25284 12124
rect 25116 10098 25172 10108
rect 25004 9828 25060 9838
rect 25004 9266 25060 9772
rect 25004 9214 25006 9266
rect 25058 9214 25060 9266
rect 25004 9202 25060 9214
rect 24668 8036 24724 8046
rect 25116 8036 25172 8046
rect 24668 7942 24724 7980
rect 25004 8034 25172 8036
rect 25004 7982 25118 8034
rect 25170 7982 25172 8034
rect 25004 7980 25172 7982
rect 24780 7362 24836 7374
rect 24780 7310 24782 7362
rect 24834 7310 24836 7362
rect 24780 6580 24836 7310
rect 24780 6514 24836 6524
rect 24892 6466 24948 6478
rect 24892 6414 24894 6466
rect 24946 6414 24948 6466
rect 24892 6356 24948 6414
rect 24444 5292 24612 5348
rect 24668 6300 24948 6356
rect 24444 3668 24500 5292
rect 24556 5122 24612 5134
rect 24556 5070 24558 5122
rect 24610 5070 24612 5122
rect 24556 4562 24612 5070
rect 24556 4510 24558 4562
rect 24610 4510 24612 4562
rect 24556 4340 24612 4510
rect 24668 5012 24724 6300
rect 24892 5796 24948 5806
rect 24668 4564 24724 4956
rect 24780 5794 24948 5796
rect 24780 5742 24894 5794
rect 24946 5742 24948 5794
rect 24780 5740 24948 5742
rect 24780 4788 24836 5740
rect 24892 5730 24948 5740
rect 24780 4722 24836 4732
rect 24892 5012 24948 5022
rect 24668 4498 24724 4508
rect 24556 4274 24612 4284
rect 24780 4450 24836 4462
rect 24780 4398 24782 4450
rect 24834 4398 24836 4450
rect 24444 3602 24500 3612
rect 24780 3892 24836 4398
rect 24892 4450 24948 4956
rect 24892 4398 24894 4450
rect 24946 4398 24948 4450
rect 24892 4386 24948 4398
rect 24556 3556 24612 3566
rect 24556 3388 24612 3500
rect 24108 3332 24276 3388
rect 24444 3332 24612 3388
rect 24108 2884 24164 3332
rect 24108 2818 24164 2828
rect 24444 980 24500 3332
rect 24780 2884 24836 3836
rect 25004 3556 25060 7980
rect 25116 7970 25172 7980
rect 25340 7364 25396 13244
rect 25788 12292 25844 15092
rect 26124 14642 26180 15092
rect 26124 14590 26126 14642
rect 26178 14590 26180 14642
rect 26124 14578 26180 14590
rect 26012 14530 26068 14542
rect 26012 14478 26014 14530
rect 26066 14478 26068 14530
rect 26012 14084 26068 14478
rect 26796 14420 26852 14430
rect 25900 14028 26292 14084
rect 25900 12962 25956 14028
rect 26236 13970 26292 14028
rect 26236 13918 26238 13970
rect 26290 13918 26292 13970
rect 26236 13906 26292 13918
rect 26012 13860 26068 13870
rect 26012 13766 26068 13804
rect 26684 13860 26740 13870
rect 26684 13766 26740 13804
rect 26124 13636 26180 13646
rect 26124 13542 26180 13580
rect 26796 13188 26852 14364
rect 27468 14308 27524 15150
rect 27692 14420 27748 14430
rect 27692 14326 27748 14364
rect 27468 13748 27524 14252
rect 27468 13654 27524 13692
rect 25900 12910 25902 12962
rect 25954 12910 25956 12962
rect 25900 12898 25956 12910
rect 26684 13132 26852 13188
rect 25564 12236 25844 12292
rect 26684 12290 26740 13132
rect 26684 12238 26686 12290
rect 26738 12238 26740 12290
rect 25452 9828 25508 9838
rect 25452 9734 25508 9772
rect 25564 7588 25620 12236
rect 26684 12226 26740 12238
rect 27356 12740 27412 12750
rect 26012 12178 26068 12190
rect 26012 12126 26014 12178
rect 26066 12126 26068 12178
rect 25788 12066 25844 12078
rect 25788 12014 25790 12066
rect 25842 12014 25844 12066
rect 25676 11508 25732 11518
rect 25676 10722 25732 11452
rect 25788 11396 25844 12014
rect 26012 11844 26068 12126
rect 26796 12180 26852 12190
rect 26012 11778 26068 11788
rect 26684 11844 26740 11854
rect 26236 11396 26292 11406
rect 26684 11396 26740 11788
rect 26796 11506 26852 12124
rect 27356 11956 27412 12684
rect 27580 11956 27636 11966
rect 27356 11954 27636 11956
rect 27356 11902 27582 11954
rect 27634 11902 27636 11954
rect 27356 11900 27636 11902
rect 27580 11620 27636 11900
rect 27580 11554 27636 11564
rect 26796 11454 26798 11506
rect 26850 11454 26852 11506
rect 26796 11442 26852 11454
rect 25788 11302 25844 11340
rect 26012 11394 26292 11396
rect 26012 11342 26238 11394
rect 26290 11342 26292 11394
rect 26012 11340 26292 11342
rect 25788 11172 25844 11182
rect 25788 10834 25844 11116
rect 25788 10782 25790 10834
rect 25842 10782 25844 10834
rect 25788 10770 25844 10782
rect 26012 10834 26068 11340
rect 26236 11330 26292 11340
rect 26460 11394 26740 11396
rect 26460 11342 26686 11394
rect 26738 11342 26740 11394
rect 26460 11340 26740 11342
rect 26012 10782 26014 10834
rect 26066 10782 26068 10834
rect 26012 10770 26068 10782
rect 26460 10834 26516 11340
rect 26684 11330 26740 11340
rect 26908 11396 26964 11406
rect 26908 11302 26964 11340
rect 26460 10782 26462 10834
rect 26514 10782 26516 10834
rect 26460 10770 26516 10782
rect 27804 10724 27860 16380
rect 28140 15538 28196 17164
rect 28588 16660 28644 18284
rect 28812 17668 28868 17678
rect 28812 17574 28868 17612
rect 29148 17668 29204 17678
rect 29148 17108 29204 17612
rect 29148 16976 29204 17052
rect 29260 16772 29316 29260
rect 29372 29250 29428 29260
rect 29596 23380 29652 30830
rect 30604 30772 30660 31502
rect 30192 30604 30456 30614
rect 30248 30548 30296 30604
rect 30352 30548 30400 30604
rect 30192 30538 30456 30548
rect 30268 30324 30324 30334
rect 30044 30212 30100 30222
rect 30044 30118 30100 30156
rect 30268 30210 30324 30268
rect 30268 30158 30270 30210
rect 30322 30158 30324 30210
rect 30268 29988 30324 30158
rect 30604 30212 30660 30716
rect 30940 30322 30996 31892
rect 31276 31780 31332 31892
rect 31612 31890 31668 31948
rect 31612 31838 31614 31890
rect 31666 31838 31668 31890
rect 31612 31826 31668 31838
rect 31164 31778 31332 31780
rect 31164 31726 31278 31778
rect 31330 31726 31332 31778
rect 31164 31724 31332 31726
rect 31164 31106 31220 31724
rect 31276 31714 31332 31724
rect 31724 31218 31780 32510
rect 31724 31166 31726 31218
rect 31778 31166 31780 31218
rect 31724 31154 31780 31166
rect 31164 31054 31166 31106
rect 31218 31054 31220 31106
rect 31164 31042 31220 31054
rect 30940 30270 30942 30322
rect 30994 30270 30996 30322
rect 30940 30258 30996 30270
rect 31052 30994 31108 31006
rect 31052 30942 31054 30994
rect 31106 30942 31108 30994
rect 31052 30324 31108 30942
rect 31612 30996 31668 31006
rect 31052 30268 31556 30324
rect 30604 30146 30660 30156
rect 30268 29922 30324 29932
rect 31052 29876 31108 30268
rect 31500 30210 31556 30268
rect 31500 30158 31502 30210
rect 31554 30158 31556 30210
rect 31500 30146 31556 30158
rect 31612 30100 31668 30940
rect 31836 30210 31892 33068
rect 33516 32676 33572 33294
rect 33628 32676 33684 32686
rect 33516 32674 33684 32676
rect 33516 32622 33630 32674
rect 33682 32622 33684 32674
rect 33516 32620 33684 32622
rect 33404 32564 33460 32574
rect 32172 32004 32228 32014
rect 32172 31778 32228 31948
rect 33404 32004 33460 32508
rect 33404 31890 33460 31948
rect 33404 31838 33406 31890
rect 33458 31838 33460 31890
rect 33404 31826 33460 31838
rect 32172 31726 32174 31778
rect 32226 31726 32228 31778
rect 32172 31714 32228 31726
rect 33180 31778 33236 31790
rect 33180 31726 33182 31778
rect 33234 31726 33236 31778
rect 33180 31556 33236 31726
rect 33180 31490 33236 31500
rect 33516 31556 33572 32620
rect 33628 32610 33684 32620
rect 33740 31890 33796 34078
rect 33964 34132 34020 34142
rect 33964 34038 34020 34076
rect 34300 34130 34356 34142
rect 34300 34078 34302 34130
rect 34354 34078 34356 34130
rect 34188 33348 34244 33358
rect 33852 33346 34244 33348
rect 33852 33294 34190 33346
rect 34242 33294 34244 33346
rect 33852 33292 34244 33294
rect 33852 32564 33908 33292
rect 34188 33282 34244 33292
rect 34188 32788 34244 32798
rect 34300 32788 34356 34078
rect 35196 34018 35252 34862
rect 35420 34916 35476 34926
rect 35420 34130 35476 34860
rect 35644 34916 35700 34926
rect 35644 34822 35700 34860
rect 36204 34802 36260 36430
rect 36540 35810 36596 37436
rect 37212 36594 37268 36606
rect 37212 36542 37214 36594
rect 37266 36542 37268 36594
rect 36540 35758 36542 35810
rect 36594 35758 36596 35810
rect 36540 35746 36596 35758
rect 36988 36260 37044 36270
rect 36988 35252 37044 36204
rect 36988 35186 37044 35196
rect 36540 34916 36596 34926
rect 36540 34822 36596 34860
rect 36204 34750 36206 34802
rect 36258 34750 36260 34802
rect 36204 34692 36260 34750
rect 36652 34804 36708 34814
rect 36652 34710 36708 34748
rect 36764 34802 36820 34814
rect 36764 34750 36766 34802
rect 36818 34750 36820 34802
rect 36204 34626 36260 34636
rect 35756 34244 35812 34254
rect 35756 34150 35812 34188
rect 35420 34078 35422 34130
rect 35474 34078 35476 34130
rect 35420 34066 35476 34078
rect 35196 33966 35198 34018
rect 35250 33966 35252 34018
rect 34972 33460 35028 33470
rect 35196 33460 35252 33966
rect 36764 33908 36820 34750
rect 36764 33842 36820 33852
rect 37212 33908 37268 36542
rect 37436 36482 37492 36494
rect 37436 36430 37438 36482
rect 37490 36430 37492 36482
rect 37436 34916 37492 36430
rect 38668 36484 38724 36494
rect 38668 36390 38724 36428
rect 39004 35810 39060 37436
rect 39004 35758 39006 35810
rect 39058 35758 39060 35810
rect 39004 35746 39060 35758
rect 39452 36370 39508 36382
rect 39452 36318 39454 36370
rect 39506 36318 39508 36370
rect 37660 35698 37716 35710
rect 37660 35646 37662 35698
rect 37714 35646 37716 35698
rect 37660 35588 37716 35646
rect 37660 35522 37716 35532
rect 38108 35588 38164 35598
rect 38108 35494 38164 35532
rect 37436 34354 37492 34860
rect 37548 34804 37604 34814
rect 37548 34710 37604 34748
rect 37660 34692 37716 34702
rect 37660 34598 37716 34636
rect 37772 34690 37828 34702
rect 37772 34638 37774 34690
rect 37826 34638 37828 34690
rect 37436 34302 37438 34354
rect 37490 34302 37492 34354
rect 37436 34290 37492 34302
rect 37548 34020 37604 34030
rect 37772 34020 37828 34638
rect 39452 34242 39508 36318
rect 39852 36092 40116 36102
rect 39908 36036 39956 36092
rect 40012 36036 40060 36092
rect 39852 36026 40116 36036
rect 40124 35924 40180 35934
rect 40124 35698 40180 35868
rect 40124 35646 40126 35698
rect 40178 35646 40180 35698
rect 40124 35634 40180 35646
rect 40236 35252 40292 37996
rect 41132 37940 41188 39200
rect 41132 37884 41524 37940
rect 41468 36594 41524 37884
rect 41468 36542 41470 36594
rect 41522 36542 41524 36594
rect 41468 36530 41524 36542
rect 42588 36482 42644 36494
rect 42588 36430 42590 36482
rect 42642 36430 42644 36482
rect 42588 36260 42644 36430
rect 42588 36194 42644 36204
rect 43036 36260 43092 36270
rect 43036 36166 43092 36204
rect 42700 36148 42756 36158
rect 40572 35924 40628 35934
rect 40572 35830 40628 35868
rect 42700 35810 42756 36092
rect 42700 35758 42702 35810
rect 42754 35758 42756 35810
rect 42700 35746 42756 35758
rect 43596 35812 43652 39200
rect 46060 37940 46116 39200
rect 46060 37884 46452 37940
rect 46396 36594 46452 37884
rect 46396 36542 46398 36594
rect 46450 36542 46452 36594
rect 46396 36530 46452 36542
rect 48524 36596 48580 39200
rect 49512 36876 49776 36886
rect 49568 36820 49616 36876
rect 49672 36820 49720 36876
rect 49512 36810 49776 36820
rect 48524 36530 48580 36540
rect 48972 36596 49028 36606
rect 48972 36502 49028 36540
rect 50988 36594 51044 39200
rect 50988 36542 50990 36594
rect 51042 36542 51044 36594
rect 50988 36530 51044 36542
rect 52220 36820 52276 36830
rect 43820 36484 43876 36494
rect 43820 36370 43876 36428
rect 47516 36484 47572 36494
rect 49868 36484 49924 36494
rect 47516 36482 47684 36484
rect 47516 36430 47518 36482
rect 47570 36430 47684 36482
rect 47516 36428 47684 36430
rect 47516 36418 47572 36428
rect 43820 36318 43822 36370
rect 43874 36318 43876 36370
rect 43820 36306 43876 36318
rect 44156 36370 44212 36382
rect 44156 36318 44158 36370
rect 44210 36318 44212 36370
rect 43932 35812 43988 35822
rect 43596 35810 43988 35812
rect 43596 35758 43934 35810
rect 43986 35758 43988 35810
rect 43596 35756 43988 35758
rect 43932 35746 43988 35756
rect 41804 35700 41860 35710
rect 39788 34916 39844 34926
rect 39676 34914 39844 34916
rect 39676 34862 39790 34914
rect 39842 34862 39844 34914
rect 39676 34860 39844 34862
rect 39676 34356 39732 34860
rect 39788 34850 39844 34860
rect 39852 34524 40116 34534
rect 39908 34468 39956 34524
rect 40012 34468 40060 34524
rect 39852 34458 40116 34468
rect 39676 34290 39732 34300
rect 39788 34356 39844 34366
rect 40236 34356 40292 35196
rect 41468 35698 41860 35700
rect 41468 35646 41806 35698
rect 41858 35646 41860 35698
rect 41468 35644 41860 35646
rect 39788 34354 40292 34356
rect 39788 34302 39790 34354
rect 39842 34302 40292 34354
rect 39788 34300 40292 34302
rect 40348 34914 40404 34926
rect 40348 34862 40350 34914
rect 40402 34862 40404 34914
rect 39788 34290 39844 34300
rect 40348 34244 40404 34862
rect 40460 34916 40516 34926
rect 40460 34822 40516 34860
rect 41356 34916 41412 34926
rect 41356 34822 41412 34860
rect 41468 34690 41524 35644
rect 41804 35634 41860 35644
rect 44156 35700 44212 36318
rect 44156 35634 44212 35644
rect 44380 36260 44436 36270
rect 42028 35586 42084 35598
rect 42028 35534 42030 35586
rect 42082 35534 42084 35586
rect 42028 34916 42084 35534
rect 42028 34850 42084 34860
rect 42588 35026 42644 35038
rect 42588 34974 42590 35026
rect 42642 34974 42644 35026
rect 41468 34638 41470 34690
rect 41522 34638 41524 34690
rect 40460 34356 40516 34366
rect 40460 34262 40516 34300
rect 40684 34356 40740 34366
rect 40684 34262 40740 34300
rect 39452 34190 39454 34242
rect 39506 34190 39508 34242
rect 39452 34178 39508 34190
rect 40124 34242 40404 34244
rect 40124 34190 40350 34242
rect 40402 34190 40404 34242
rect 40124 34188 40404 34190
rect 37548 34018 37828 34020
rect 37548 33966 37550 34018
rect 37602 33966 37828 34018
rect 37548 33964 37828 33966
rect 37548 33954 37604 33964
rect 37212 33814 37268 33852
rect 38668 33908 38724 33918
rect 34972 33458 35252 33460
rect 34972 33406 34974 33458
rect 35026 33406 35252 33458
rect 34972 33404 35252 33406
rect 37884 33458 37940 33470
rect 37884 33406 37886 33458
rect 37938 33406 37940 33458
rect 34972 33394 35028 33404
rect 37324 33348 37380 33358
rect 36876 33124 36932 33134
rect 36876 33030 36932 33068
rect 34188 32786 34356 32788
rect 34188 32734 34190 32786
rect 34242 32734 34356 32786
rect 34188 32732 34356 32734
rect 34188 32722 34244 32732
rect 33852 32432 33908 32508
rect 37324 32562 37380 33292
rect 37884 32676 37940 33406
rect 37996 33346 38052 33358
rect 37996 33294 37998 33346
rect 38050 33294 38052 33346
rect 37996 33124 38052 33294
rect 37996 33058 38052 33068
rect 38556 33124 38612 33134
rect 38556 32786 38612 33068
rect 38556 32734 38558 32786
rect 38610 32734 38612 32786
rect 38556 32722 38612 32734
rect 38668 32786 38724 33852
rect 40124 33458 40180 34188
rect 40348 34178 40404 34188
rect 41468 34244 41524 34638
rect 41468 34178 41524 34188
rect 41692 34690 41748 34702
rect 41692 34638 41694 34690
rect 41746 34638 41748 34690
rect 41692 34244 41748 34638
rect 41692 34178 41748 34188
rect 42476 34356 42532 34366
rect 42588 34356 42644 34974
rect 44044 34914 44100 34926
rect 44044 34862 44046 34914
rect 44098 34862 44100 34914
rect 42476 34354 42644 34356
rect 42476 34302 42478 34354
rect 42530 34302 42644 34354
rect 42476 34300 42644 34302
rect 42812 34802 42868 34814
rect 42812 34750 42814 34802
rect 42866 34750 42868 34802
rect 42812 34356 42868 34750
rect 42252 33908 42308 33918
rect 42252 33814 42308 33852
rect 40124 33406 40126 33458
rect 40178 33406 40180 33458
rect 40124 33394 40180 33406
rect 42476 33460 42532 34300
rect 42812 34290 42868 34300
rect 43484 34692 43540 34702
rect 43484 34354 43540 34636
rect 43484 34302 43486 34354
rect 43538 34302 43540 34354
rect 43484 34290 43540 34302
rect 43596 34356 43652 34366
rect 43148 34130 43204 34142
rect 43148 34078 43150 34130
rect 43202 34078 43204 34130
rect 42588 34020 42644 34030
rect 43148 34020 43204 34078
rect 43596 34130 43652 34300
rect 43932 34244 43988 34254
rect 43932 34150 43988 34188
rect 43596 34078 43598 34130
rect 43650 34078 43652 34130
rect 43596 34066 43652 34078
rect 42588 34018 43204 34020
rect 42588 33966 42590 34018
rect 42642 33966 43204 34018
rect 42588 33964 43204 33966
rect 42588 33954 42644 33964
rect 43484 33906 43540 33918
rect 43484 33854 43486 33906
rect 43538 33854 43540 33906
rect 42812 33796 42868 33806
rect 42812 33570 42868 33740
rect 42812 33518 42814 33570
rect 42866 33518 42868 33570
rect 42812 33506 42868 33518
rect 42588 33460 42644 33470
rect 42476 33458 42644 33460
rect 42476 33406 42590 33458
rect 42642 33406 42644 33458
rect 42476 33404 42644 33406
rect 39340 33348 39396 33358
rect 39340 33254 39396 33292
rect 38668 32734 38670 32786
rect 38722 32734 38724 32786
rect 38668 32722 38724 32734
rect 39228 33124 39284 33134
rect 39228 32786 39284 33068
rect 39852 32956 40116 32966
rect 39908 32900 39956 32956
rect 40012 32900 40060 32956
rect 39852 32890 40116 32900
rect 39228 32734 39230 32786
rect 39282 32734 39284 32786
rect 39228 32722 39284 32734
rect 42364 32788 42420 32798
rect 42476 32788 42532 33404
rect 42588 33394 42644 33404
rect 43148 33348 43204 33358
rect 43148 33254 43204 33292
rect 43484 33348 43540 33854
rect 44044 33908 44100 34862
rect 44044 33842 44100 33852
rect 43484 33282 43540 33292
rect 43932 33458 43988 33470
rect 43932 33406 43934 33458
rect 43986 33406 43988 33458
rect 42364 32786 42532 32788
rect 42364 32734 42366 32786
rect 42418 32734 42532 32786
rect 42364 32732 42532 32734
rect 43932 33236 43988 33406
rect 44268 33348 44324 33358
rect 44268 33254 44324 33292
rect 42364 32722 42420 32732
rect 37324 32510 37326 32562
rect 37378 32510 37380 32562
rect 37100 32452 37156 32462
rect 37100 32358 37156 32396
rect 37324 32004 37380 32510
rect 33740 31838 33742 31890
rect 33794 31838 33796 31890
rect 33740 31826 33796 31838
rect 37100 31892 37380 31948
rect 37548 32620 37940 32676
rect 37548 32452 37604 32620
rect 38108 32564 38164 32574
rect 33516 31490 33572 31500
rect 35532 31106 35588 31118
rect 35532 31054 35534 31106
rect 35586 31054 35588 31106
rect 32284 30884 32340 30894
rect 32732 30884 32788 30894
rect 33852 30884 33908 30894
rect 32284 30882 32788 30884
rect 32284 30830 32286 30882
rect 32338 30830 32734 30882
rect 32786 30830 32788 30882
rect 32284 30828 32788 30830
rect 32060 30772 32116 30782
rect 32060 30678 32116 30716
rect 32284 30324 32340 30828
rect 32732 30818 32788 30828
rect 33740 30882 33908 30884
rect 33740 30830 33854 30882
rect 33906 30830 33908 30882
rect 33740 30828 33908 30830
rect 33740 30324 33796 30828
rect 33852 30818 33908 30828
rect 34412 30884 34468 30894
rect 34972 30884 35028 30894
rect 34412 30882 35028 30884
rect 34412 30830 34414 30882
rect 34466 30830 34974 30882
rect 35026 30830 35028 30882
rect 34412 30828 35028 30830
rect 32284 30258 32340 30268
rect 33516 30268 33740 30324
rect 31836 30158 31838 30210
rect 31890 30158 31892 30210
rect 31836 30146 31892 30158
rect 31612 29968 31668 30044
rect 32172 30100 32228 30110
rect 32172 30006 32228 30044
rect 32732 30098 32788 30110
rect 32732 30046 32734 30098
rect 32786 30046 32788 30098
rect 30604 29820 31108 29876
rect 29820 29764 29876 29774
rect 29820 29650 29876 29708
rect 29820 29598 29822 29650
rect 29874 29598 29876 29650
rect 29820 29586 29876 29598
rect 30192 29036 30456 29046
rect 30248 28980 30296 29036
rect 30352 28980 30400 29036
rect 30192 28970 30456 28980
rect 30604 28754 30660 29820
rect 32732 29652 32788 30046
rect 32284 29596 32788 29652
rect 32844 29986 32900 29998
rect 32844 29934 32846 29986
rect 32898 29934 32900 29986
rect 30604 28702 30606 28754
rect 30658 28702 30660 28754
rect 30604 28690 30660 28702
rect 32060 29316 32116 29326
rect 32284 29316 32340 29596
rect 32844 29540 32900 29934
rect 32060 29314 32340 29316
rect 32060 29262 32062 29314
rect 32114 29262 32340 29314
rect 32396 29484 32900 29540
rect 33068 29986 33124 29998
rect 33068 29934 33070 29986
rect 33122 29934 33124 29986
rect 33068 29540 33124 29934
rect 33404 29988 33460 29998
rect 33516 29988 33572 30268
rect 33740 30192 33796 30268
rect 33852 30324 33908 30334
rect 34412 30324 34468 30828
rect 34972 30818 35028 30828
rect 33852 30322 34468 30324
rect 33852 30270 33854 30322
rect 33906 30270 34468 30322
rect 33852 30268 34468 30270
rect 34524 30660 34580 30670
rect 34524 30324 34580 30604
rect 33852 30258 33908 30268
rect 33404 29986 33572 29988
rect 33404 29934 33406 29986
rect 33458 29934 33572 29986
rect 33404 29932 33572 29934
rect 33404 29922 33460 29932
rect 32396 29428 32452 29484
rect 33068 29474 33124 29484
rect 32396 29296 32452 29372
rect 32732 29316 32788 29326
rect 32060 29260 32340 29262
rect 32060 28754 32116 29260
rect 32732 29222 32788 29260
rect 32060 28702 32062 28754
rect 32114 28702 32116 28754
rect 32060 28690 32116 28702
rect 32396 28754 32452 28766
rect 32396 28702 32398 28754
rect 32450 28702 32452 28754
rect 29708 28644 29764 28654
rect 29708 28550 29764 28588
rect 29932 28642 29988 28654
rect 29932 28590 29934 28642
rect 29986 28590 29988 28642
rect 29932 28532 29988 28590
rect 29932 28466 29988 28476
rect 31052 28644 31108 28654
rect 30716 27972 30772 27982
rect 30604 27916 30716 27972
rect 30044 27860 30100 27870
rect 30044 27766 30100 27804
rect 30192 27468 30456 27478
rect 30248 27412 30296 27468
rect 30352 27412 30400 27468
rect 30192 27402 30456 27412
rect 30604 27188 30660 27916
rect 30716 27878 30772 27916
rect 30828 27860 30884 27870
rect 30828 27766 30884 27804
rect 30716 27636 30772 27646
rect 30716 27542 30772 27580
rect 30940 27188 30996 27198
rect 30604 27186 30996 27188
rect 30604 27134 30942 27186
rect 30994 27134 30996 27186
rect 30604 27132 30996 27134
rect 30940 26964 30996 27132
rect 30940 26898 30996 26908
rect 29820 26292 29876 26302
rect 29820 26198 29876 26236
rect 30940 26292 30996 26302
rect 30940 26198 30996 26236
rect 29708 26178 29764 26190
rect 29708 26126 29710 26178
rect 29762 26126 29764 26178
rect 29708 25620 29764 26126
rect 30492 26178 30548 26190
rect 30492 26126 30494 26178
rect 30546 26126 30548 26178
rect 29708 25554 29764 25564
rect 29820 26068 29876 26078
rect 29596 23314 29652 23324
rect 29708 23828 29764 23838
rect 29708 21698 29764 23772
rect 29820 23266 29876 26012
rect 30492 26068 30548 26126
rect 30492 26002 30548 26012
rect 30192 25900 30456 25910
rect 30248 25844 30296 25900
rect 30352 25844 30400 25900
rect 30192 25834 30456 25844
rect 30940 25396 30996 25406
rect 30604 24836 30660 24846
rect 30492 24724 30548 24734
rect 30492 24630 30548 24668
rect 30044 24610 30100 24622
rect 30044 24558 30046 24610
rect 30098 24558 30100 24610
rect 30044 23828 30100 24558
rect 30192 24332 30456 24342
rect 30248 24276 30296 24332
rect 30352 24276 30400 24332
rect 30192 24266 30456 24276
rect 30604 23938 30660 24780
rect 30940 24834 30996 25340
rect 30940 24782 30942 24834
rect 30994 24782 30996 24834
rect 30940 24770 30996 24782
rect 30604 23886 30606 23938
rect 30658 23886 30660 23938
rect 30604 23874 30660 23886
rect 30716 24724 30772 24734
rect 30044 23762 30100 23772
rect 30268 23828 30324 23838
rect 30268 23734 30324 23772
rect 30380 23716 30436 23726
rect 30380 23622 30436 23660
rect 30716 23716 30772 24668
rect 31052 24500 31108 28588
rect 31612 28644 31668 28654
rect 31612 28550 31668 28588
rect 32396 28532 32452 28702
rect 32508 28644 32564 28654
rect 32508 28550 32564 28588
rect 31164 28418 31220 28430
rect 31164 28366 31166 28418
rect 31218 28366 31220 28418
rect 31164 27860 31220 28366
rect 31164 27794 31220 27804
rect 31612 27858 31668 27870
rect 31612 27806 31614 27858
rect 31666 27806 31668 27858
rect 31612 27636 31668 27806
rect 31612 27570 31668 27580
rect 31724 27860 31780 27870
rect 31388 27076 31444 27086
rect 31388 26402 31444 27020
rect 31500 26964 31556 26974
rect 31500 26870 31556 26908
rect 31724 26964 31780 27804
rect 32060 27746 32116 27758
rect 32060 27694 32062 27746
rect 32114 27694 32116 27746
rect 31724 26870 31780 26908
rect 31836 27186 31892 27198
rect 31836 27134 31838 27186
rect 31890 27134 31892 27186
rect 31388 26350 31390 26402
rect 31442 26350 31444 26402
rect 31388 26338 31444 26350
rect 31836 26292 31892 27134
rect 32060 27076 32116 27694
rect 32396 27746 32452 28476
rect 32396 27694 32398 27746
rect 32450 27694 32452 27746
rect 32396 27682 32452 27694
rect 32060 26944 32116 27020
rect 32396 26964 32452 26974
rect 32396 26870 32452 26908
rect 31948 26292 32004 26302
rect 31836 26290 32004 26292
rect 31836 26238 31950 26290
rect 32002 26238 32004 26290
rect 31836 26236 32004 26238
rect 31948 26226 32004 26236
rect 32284 26292 32340 26302
rect 32284 26198 32340 26236
rect 32508 26290 32564 26302
rect 32508 26238 32510 26290
rect 32562 26238 32564 26290
rect 32396 26180 32452 26190
rect 32396 26086 32452 26124
rect 32508 26068 32564 26238
rect 32508 26002 32564 26012
rect 33068 25508 33124 25518
rect 33068 25394 33124 25452
rect 33068 25342 33070 25394
rect 33122 25342 33124 25394
rect 33068 25330 33124 25342
rect 33180 25396 33236 25406
rect 33180 25302 33236 25340
rect 32844 25282 32900 25294
rect 32844 25230 32846 25282
rect 32898 25230 32900 25282
rect 32732 24836 32788 24846
rect 32732 24742 32788 24780
rect 32844 24834 32900 25230
rect 32844 24782 32846 24834
rect 32898 24782 32900 24834
rect 32844 24770 32900 24782
rect 32508 24724 32564 24734
rect 32508 24630 32564 24668
rect 31052 24434 31108 24444
rect 32844 24612 32900 24622
rect 30716 23650 30772 23660
rect 32620 23716 32676 23726
rect 32620 23622 32676 23660
rect 29820 23214 29822 23266
rect 29874 23214 29876 23266
rect 29820 23202 29876 23214
rect 30192 22764 30456 22774
rect 30248 22708 30296 22764
rect 30352 22708 30400 22764
rect 30192 22698 30456 22708
rect 30716 22708 30772 22718
rect 29708 21646 29710 21698
rect 29762 21646 29764 21698
rect 29708 21634 29764 21646
rect 30604 22148 30660 22158
rect 30192 21196 30456 21206
rect 30248 21140 30296 21196
rect 30352 21140 30400 21196
rect 30192 21130 30456 21140
rect 30604 21028 30660 22092
rect 30716 21700 30772 22652
rect 32060 22372 32116 22382
rect 30716 21634 30772 21644
rect 31948 22370 32116 22372
rect 31948 22318 32062 22370
rect 32114 22318 32116 22370
rect 31948 22316 32116 22318
rect 31948 21698 32004 22316
rect 32060 22306 32116 22316
rect 32508 22372 32564 22382
rect 32508 22370 32788 22372
rect 32508 22318 32510 22370
rect 32562 22318 32788 22370
rect 32508 22316 32788 22318
rect 32508 22306 32564 22316
rect 31948 21646 31950 21698
rect 32002 21646 32004 21698
rect 30604 20962 30660 20972
rect 30268 20914 30324 20926
rect 30268 20862 30270 20914
rect 30322 20862 30324 20914
rect 29708 20692 29764 20702
rect 29596 20578 29652 20590
rect 29596 20526 29598 20578
rect 29650 20526 29652 20578
rect 29596 20356 29652 20526
rect 29596 20290 29652 20300
rect 29708 20242 29764 20636
rect 29708 20190 29710 20242
rect 29762 20190 29764 20242
rect 29708 20178 29764 20190
rect 29596 20018 29652 20030
rect 29596 19966 29598 20018
rect 29650 19966 29652 20018
rect 29596 19908 29652 19966
rect 29932 20020 29988 20030
rect 30268 20020 30324 20862
rect 30604 20690 30660 20702
rect 30604 20638 30606 20690
rect 30658 20638 30660 20690
rect 30380 20020 30436 20030
rect 29932 20018 30436 20020
rect 29932 19966 29934 20018
rect 29986 19966 30382 20018
rect 30434 19966 30436 20018
rect 29932 19964 30436 19966
rect 29932 19954 29988 19964
rect 30380 19954 30436 19964
rect 29596 19842 29652 19852
rect 30604 19796 30660 20638
rect 31948 20578 32004 21646
rect 32732 21698 32788 22316
rect 32732 21646 32734 21698
rect 32786 21646 32788 21698
rect 32060 21588 32116 21598
rect 32620 21588 32676 21598
rect 32060 21586 32676 21588
rect 32060 21534 32062 21586
rect 32114 21534 32622 21586
rect 32674 21534 32676 21586
rect 32060 21532 32676 21534
rect 32060 21522 32116 21532
rect 32620 21522 32676 21532
rect 31948 20526 31950 20578
rect 32002 20526 32004 20578
rect 31948 20514 32004 20526
rect 32060 20690 32116 20702
rect 32060 20638 32062 20690
rect 32114 20638 32116 20690
rect 30828 20244 30884 20254
rect 30192 19628 30456 19638
rect 30248 19572 30296 19628
rect 30352 19572 30400 19628
rect 30192 19562 30456 19572
rect 30604 19460 30660 19740
rect 30268 19404 30660 19460
rect 30716 20018 30772 20030
rect 30716 19966 30718 20018
rect 30770 19966 30772 20018
rect 30716 19460 30772 19966
rect 30828 20018 30884 20188
rect 30828 19966 30830 20018
rect 30882 19966 30884 20018
rect 30828 19954 30884 19966
rect 31052 20018 31108 20030
rect 31052 19966 31054 20018
rect 31106 19966 31108 20018
rect 30940 19906 30996 19918
rect 30940 19854 30942 19906
rect 30994 19854 30996 19906
rect 30828 19460 30884 19470
rect 30716 19458 30884 19460
rect 30716 19406 30830 19458
rect 30882 19406 30884 19458
rect 30716 19404 30884 19406
rect 30268 19346 30324 19404
rect 30828 19394 30884 19404
rect 30268 19294 30270 19346
rect 30322 19294 30324 19346
rect 30268 19282 30324 19294
rect 30492 19234 30548 19246
rect 30492 19182 30494 19234
rect 30546 19182 30548 19234
rect 30492 19124 30548 19182
rect 30940 19236 30996 19854
rect 30940 19170 30996 19180
rect 30492 19058 30548 19068
rect 29708 19012 29764 19022
rect 29596 19010 29764 19012
rect 29596 18958 29710 19010
rect 29762 18958 29764 19010
rect 29596 18956 29764 18958
rect 29596 18900 29652 18956
rect 29708 18946 29764 18956
rect 29596 17444 29652 18844
rect 29596 17350 29652 17388
rect 29932 18564 29988 18574
rect 29260 16706 29316 16716
rect 29596 16772 29652 16782
rect 28588 16594 28644 16604
rect 29596 15986 29652 16716
rect 29596 15934 29598 15986
rect 29650 15934 29652 15986
rect 28812 15876 28868 15886
rect 28924 15876 28980 15886
rect 28812 15874 28924 15876
rect 28812 15822 28814 15874
rect 28866 15822 28924 15874
rect 28812 15820 28924 15822
rect 28812 15810 28868 15820
rect 28140 15486 28142 15538
rect 28194 15486 28196 15538
rect 28140 15474 28196 15486
rect 28028 15314 28084 15326
rect 28028 15262 28030 15314
rect 28082 15262 28084 15314
rect 28028 14754 28084 15262
rect 28252 15314 28308 15326
rect 28252 15262 28254 15314
rect 28306 15262 28308 15314
rect 28252 15148 28308 15262
rect 28028 14702 28030 14754
rect 28082 14702 28084 14754
rect 28028 14690 28084 14702
rect 28140 15092 28308 15148
rect 28700 15314 28756 15326
rect 28700 15262 28702 15314
rect 28754 15262 28756 15314
rect 28028 14530 28084 14542
rect 28028 14478 28030 14530
rect 28082 14478 28084 14530
rect 28028 14308 28084 14478
rect 28028 13636 28084 14252
rect 28140 13748 28196 15092
rect 28700 14754 28756 15262
rect 28700 14702 28702 14754
rect 28754 14702 28756 14754
rect 28700 14690 28756 14702
rect 28812 14420 28868 14430
rect 28700 14308 28756 14318
rect 28700 14214 28756 14252
rect 28140 13654 28196 13692
rect 28812 13748 28868 14364
rect 28812 13682 28868 13692
rect 28028 13542 28084 13580
rect 28924 13300 28980 15820
rect 29596 15204 29652 15934
rect 29708 16548 29764 16558
rect 29708 15876 29764 16492
rect 29708 15782 29764 15820
rect 29932 15874 29988 18508
rect 31052 18564 31108 19966
rect 31052 18498 31108 18508
rect 31164 19908 31220 19918
rect 30156 18452 30212 18462
rect 30156 18358 30212 18396
rect 30604 18340 30660 18350
rect 30192 18060 30456 18070
rect 30248 18004 30296 18060
rect 30352 18004 30400 18060
rect 30192 17994 30456 18004
rect 30492 17668 30548 17678
rect 30604 17668 30660 18284
rect 31164 18004 31220 19852
rect 32060 19572 32116 20638
rect 32732 20580 32788 21646
rect 32732 20514 32788 20524
rect 31724 19516 32116 19572
rect 31724 19234 31780 19516
rect 31724 19182 31726 19234
rect 31778 19182 31780 19234
rect 31388 19122 31444 19134
rect 31724 19124 31780 19182
rect 31388 19070 31390 19122
rect 31442 19070 31444 19122
rect 31388 18900 31444 19070
rect 31612 19068 31724 19124
rect 31500 19012 31556 19022
rect 31500 18918 31556 18956
rect 31388 18834 31444 18844
rect 31388 18676 31444 18686
rect 31388 18582 31444 18620
rect 31276 18562 31332 18574
rect 31276 18510 31278 18562
rect 31330 18510 31332 18562
rect 31276 18340 31332 18510
rect 31276 18274 31332 18284
rect 31164 17948 31332 18004
rect 30492 17666 30660 17668
rect 30492 17614 30494 17666
rect 30546 17614 30660 17666
rect 30492 17612 30660 17614
rect 31164 17778 31220 17790
rect 31164 17726 31166 17778
rect 31218 17726 31220 17778
rect 30492 17602 30548 17612
rect 30156 17554 30212 17566
rect 30156 17502 30158 17554
rect 30210 17502 30212 17554
rect 30156 17444 30212 17502
rect 30156 17378 30212 17388
rect 30268 17442 30324 17454
rect 30268 17390 30270 17442
rect 30322 17390 30324 17442
rect 30268 17108 30324 17390
rect 30156 16882 30212 16894
rect 30156 16830 30158 16882
rect 30210 16830 30212 16882
rect 30156 16772 30212 16830
rect 30156 16706 30212 16716
rect 30268 16660 30324 17052
rect 30492 17108 30548 17118
rect 31164 17108 31220 17726
rect 30492 17106 31220 17108
rect 30492 17054 30494 17106
rect 30546 17054 31220 17106
rect 30492 17052 31220 17054
rect 30492 17042 30548 17052
rect 30828 16884 30884 16894
rect 30268 16604 30660 16660
rect 30192 16492 30456 16502
rect 30248 16436 30296 16492
rect 30352 16436 30400 16492
rect 30192 16426 30456 16436
rect 30268 16212 30324 16222
rect 30268 16118 30324 16156
rect 29932 15822 29934 15874
rect 29986 15822 29988 15874
rect 29932 15428 29988 15822
rect 30604 15876 30660 16604
rect 30828 16212 30884 16828
rect 31164 16882 31220 17052
rect 31164 16830 31166 16882
rect 31218 16830 31220 16882
rect 31164 16818 31220 16830
rect 30828 16098 30884 16156
rect 30828 16046 30830 16098
rect 30882 16046 30884 16098
rect 30828 16034 30884 16046
rect 30940 15876 30996 15886
rect 30604 15874 30996 15876
rect 30604 15822 30942 15874
rect 30994 15822 30996 15874
rect 30604 15820 30996 15822
rect 30492 15540 30548 15550
rect 30604 15540 30660 15820
rect 30940 15810 30996 15820
rect 31164 15876 31220 15886
rect 31164 15782 31220 15820
rect 30492 15538 30660 15540
rect 30492 15486 30494 15538
rect 30546 15486 30660 15538
rect 30492 15484 30660 15486
rect 30492 15474 30548 15484
rect 29932 15362 29988 15372
rect 29596 15138 29652 15148
rect 30044 15204 30100 15214
rect 30044 15110 30100 15148
rect 30716 15204 30772 15214
rect 30192 14924 30456 14934
rect 30248 14868 30296 14924
rect 30352 14868 30400 14924
rect 30192 14858 30456 14868
rect 30156 13860 30212 13870
rect 30156 13766 30212 13804
rect 29484 13748 29540 13758
rect 29484 13654 29540 13692
rect 30192 13356 30456 13366
rect 30248 13300 30296 13356
rect 30352 13300 30400 13356
rect 30192 13290 30456 13300
rect 28924 13234 28980 13244
rect 28476 13188 28532 13198
rect 28028 12740 28084 12750
rect 28028 12646 28084 12684
rect 27916 12180 27972 12218
rect 27916 12114 27972 12124
rect 28364 12068 28420 12078
rect 27916 11954 27972 11966
rect 27916 11902 27918 11954
rect 27970 11902 27972 11954
rect 27916 11396 27972 11902
rect 27916 11330 27972 11340
rect 28140 11170 28196 11182
rect 28140 11118 28142 11170
rect 28194 11118 28196 11170
rect 28140 10836 28196 11118
rect 28140 10770 28196 10780
rect 25676 10670 25678 10722
rect 25730 10670 25732 10722
rect 25676 10658 25732 10670
rect 27692 10668 27860 10724
rect 27020 10500 27076 10510
rect 26796 10388 26852 10398
rect 26796 9940 26852 10332
rect 26908 9940 26964 9950
rect 26796 9938 26964 9940
rect 26796 9886 26910 9938
rect 26962 9886 26964 9938
rect 26796 9884 26964 9886
rect 26908 9874 26964 9884
rect 27020 9940 27076 10444
rect 26012 9826 26068 9838
rect 26012 9774 26014 9826
rect 26066 9774 26068 9826
rect 25900 9268 25956 9278
rect 25900 9174 25956 9212
rect 26012 9156 26068 9774
rect 26124 9828 26180 9838
rect 26236 9828 26292 9838
rect 26180 9826 26292 9828
rect 26180 9774 26238 9826
rect 26290 9774 26292 9826
rect 26180 9772 26292 9774
rect 26124 9266 26180 9772
rect 26236 9762 26292 9772
rect 26124 9214 26126 9266
rect 26178 9214 26180 9266
rect 26124 9202 26180 9214
rect 26236 9268 26292 9278
rect 26236 9174 26292 9212
rect 27020 9266 27076 9884
rect 27020 9214 27022 9266
rect 27074 9214 27076 9266
rect 26012 9090 26068 9100
rect 26348 9156 26404 9166
rect 26348 9062 26404 9100
rect 26908 8260 26964 8270
rect 26908 8166 26964 8204
rect 26348 8148 26404 8158
rect 26348 8054 26404 8092
rect 27020 8146 27076 9214
rect 27692 8930 27748 10668
rect 28252 10610 28308 10622
rect 28252 10558 28254 10610
rect 28306 10558 28308 10610
rect 27804 10498 27860 10510
rect 27804 10446 27806 10498
rect 27858 10446 27860 10498
rect 27804 9940 27860 10446
rect 27804 9874 27860 9884
rect 28252 9828 28308 10558
rect 28140 9602 28196 9614
rect 28140 9550 28142 9602
rect 28194 9550 28196 9602
rect 28140 9044 28196 9550
rect 28140 8950 28196 8988
rect 27692 8878 27694 8930
rect 27746 8878 27748 8930
rect 27020 8094 27022 8146
rect 27074 8094 27076 8146
rect 26684 7812 26740 7822
rect 26684 7700 26740 7756
rect 26572 7698 26740 7700
rect 26572 7646 26686 7698
rect 26738 7646 26740 7698
rect 26572 7644 26740 7646
rect 27020 7700 27076 8094
rect 27244 8148 27300 8158
rect 27132 7700 27188 7710
rect 27020 7698 27188 7700
rect 27020 7646 27134 7698
rect 27186 7646 27188 7698
rect 27020 7644 27188 7646
rect 26348 7588 26404 7598
rect 25564 7532 25732 7588
rect 25340 7298 25396 7308
rect 25564 7362 25620 7374
rect 25564 7310 25566 7362
rect 25618 7310 25620 7362
rect 25116 6692 25172 6702
rect 25116 6466 25172 6636
rect 25116 6414 25118 6466
rect 25170 6414 25172 6466
rect 25116 6020 25172 6414
rect 25116 5954 25172 5964
rect 25228 6580 25284 6590
rect 25004 3490 25060 3500
rect 24780 2818 24836 2828
rect 25228 1204 25284 6524
rect 25564 6580 25620 7310
rect 25564 6514 25620 6524
rect 25676 6244 25732 7532
rect 26012 7362 26068 7374
rect 26012 7310 26014 7362
rect 26066 7310 26068 7362
rect 26012 6692 26068 7310
rect 26012 6626 26068 6636
rect 26348 6692 26404 7532
rect 26572 6804 26628 7644
rect 26684 7634 26740 7644
rect 27132 7634 27188 7644
rect 27244 6916 27300 8092
rect 27692 8036 27748 8878
rect 27692 7970 27748 7980
rect 28028 8148 28084 8158
rect 28028 7474 28084 8092
rect 28252 7588 28308 9772
rect 28364 8484 28420 12012
rect 28476 10724 28532 13132
rect 30716 13188 30772 15148
rect 29260 12852 29316 12862
rect 28588 12180 28644 12190
rect 28588 12066 28644 12124
rect 28588 12014 28590 12066
rect 28642 12014 28644 12066
rect 28588 12002 28644 12014
rect 28812 12178 28868 12190
rect 28812 12126 28814 12178
rect 28866 12126 28868 12178
rect 28812 11170 28868 12126
rect 28812 11118 28814 11170
rect 28866 11118 28868 11170
rect 28812 10836 28868 11118
rect 28812 10770 28868 10780
rect 28476 10658 28532 10668
rect 28812 9940 28868 9950
rect 28476 9828 28532 9838
rect 28476 9734 28532 9772
rect 28812 9266 28868 9884
rect 29260 9380 29316 12796
rect 29596 12850 29652 12862
rect 29596 12798 29598 12850
rect 29650 12798 29652 12850
rect 29596 12740 29652 12798
rect 29596 12674 29652 12684
rect 29708 12738 29764 12750
rect 29708 12686 29710 12738
rect 29762 12686 29764 12738
rect 29708 12180 29764 12686
rect 29708 12114 29764 12124
rect 29932 12738 29988 12750
rect 29932 12686 29934 12738
rect 29986 12686 29988 12738
rect 29708 11956 29764 11966
rect 29708 11506 29764 11900
rect 29708 11454 29710 11506
rect 29762 11454 29764 11506
rect 29708 11442 29764 11454
rect 29596 11396 29652 11406
rect 29596 11302 29652 11340
rect 29932 11284 29988 12686
rect 30044 12740 30100 12750
rect 30044 12178 30100 12684
rect 30268 12740 30324 12750
rect 30268 12646 30324 12684
rect 30044 12126 30046 12178
rect 30098 12126 30100 12178
rect 30044 12114 30100 12126
rect 30192 11788 30456 11798
rect 30248 11732 30296 11788
rect 30352 11732 30400 11788
rect 30192 11722 30456 11732
rect 30044 11284 30100 11294
rect 29932 11282 30100 11284
rect 29932 11230 30046 11282
rect 30098 11230 30100 11282
rect 29932 11228 30100 11230
rect 30044 11218 30100 11228
rect 29820 11170 29876 11182
rect 29820 11118 29822 11170
rect 29874 11118 29876 11170
rect 29820 10836 29876 11118
rect 29820 10770 29876 10780
rect 29932 11060 29988 11070
rect 29484 10610 29540 10622
rect 29484 10558 29486 10610
rect 29538 10558 29540 10610
rect 29372 10498 29428 10510
rect 29372 10446 29374 10498
rect 29426 10446 29428 10498
rect 29372 9716 29428 10446
rect 29484 9940 29540 10558
rect 29820 10500 29876 10510
rect 29820 10406 29876 10444
rect 29484 9884 29764 9940
rect 29596 9716 29652 9726
rect 29372 9714 29652 9716
rect 29372 9662 29598 9714
rect 29650 9662 29652 9714
rect 29372 9660 29652 9662
rect 28812 9214 28814 9266
rect 28866 9214 28868 9266
rect 28812 9202 28868 9214
rect 29036 9324 29540 9380
rect 28700 9044 28756 9054
rect 28700 8950 28756 8988
rect 28812 8820 28868 8830
rect 28588 8764 28812 8820
rect 28364 8428 28532 8484
rect 28364 8258 28420 8270
rect 28364 8206 28366 8258
rect 28418 8206 28420 8258
rect 28364 7700 28420 8206
rect 28476 8260 28532 8428
rect 28588 8370 28644 8764
rect 28812 8726 28868 8764
rect 28588 8318 28590 8370
rect 28642 8318 28644 8370
rect 28588 8306 28644 8318
rect 28476 8036 28532 8204
rect 28812 8260 28868 8270
rect 28812 8166 28868 8204
rect 28476 7980 28980 8036
rect 28700 7700 28756 7710
rect 28364 7698 28756 7700
rect 28364 7646 28702 7698
rect 28754 7646 28756 7698
rect 28364 7644 28756 7646
rect 28252 7532 28532 7588
rect 28028 7422 28030 7474
rect 28082 7422 28084 7474
rect 28028 7410 28084 7422
rect 28252 7364 28308 7374
rect 28140 7362 28308 7364
rect 28140 7310 28254 7362
rect 28306 7310 28308 7362
rect 28140 7308 28308 7310
rect 27020 6860 27300 6916
rect 27692 7250 27748 7262
rect 27692 7198 27694 7250
rect 27746 7198 27748 7250
rect 26572 6748 26964 6804
rect 26348 6690 26852 6692
rect 26348 6638 26350 6690
rect 26402 6638 26852 6690
rect 26348 6636 26852 6638
rect 26348 6626 26404 6636
rect 26796 6578 26852 6636
rect 26796 6526 26798 6578
rect 26850 6526 26852 6578
rect 26796 6514 26852 6526
rect 25788 6468 25844 6478
rect 25788 6374 25844 6412
rect 26908 6466 26964 6748
rect 26908 6414 26910 6466
rect 26962 6414 26964 6466
rect 25676 6188 25844 6244
rect 25676 6020 25732 6030
rect 25676 5794 25732 5964
rect 25676 5742 25678 5794
rect 25730 5742 25732 5794
rect 25564 5682 25620 5694
rect 25564 5630 25566 5682
rect 25618 5630 25620 5682
rect 25452 5346 25508 5358
rect 25452 5294 25454 5346
rect 25506 5294 25508 5346
rect 25452 5236 25508 5294
rect 25452 5170 25508 5180
rect 25564 5122 25620 5630
rect 25564 5070 25566 5122
rect 25618 5070 25620 5122
rect 25564 5058 25620 5070
rect 25452 5012 25508 5022
rect 25452 3666 25508 4956
rect 25676 4676 25732 5742
rect 25676 4610 25732 4620
rect 25676 4340 25732 4350
rect 25676 4246 25732 4284
rect 25452 3614 25454 3666
rect 25506 3614 25508 3666
rect 25452 3602 25508 3614
rect 25788 3332 25844 6188
rect 26236 5794 26292 5806
rect 26236 5742 26238 5794
rect 26290 5742 26292 5794
rect 26236 4788 26292 5742
rect 26684 5794 26740 5806
rect 26684 5742 26686 5794
rect 26738 5742 26740 5794
rect 26124 4564 26180 4574
rect 26236 4564 26292 4732
rect 26460 5682 26516 5694
rect 26460 5630 26462 5682
rect 26514 5630 26516 5682
rect 26460 5122 26516 5630
rect 26684 5460 26740 5742
rect 26684 5394 26740 5404
rect 26908 5236 26964 6414
rect 27020 6468 27076 6860
rect 27692 6804 27748 7198
rect 27804 6804 27860 6814
rect 27692 6802 27860 6804
rect 27692 6750 27806 6802
rect 27858 6750 27860 6802
rect 27692 6748 27860 6750
rect 27804 6738 27860 6748
rect 28140 6804 28196 7308
rect 28252 7298 28308 7308
rect 28140 6738 28196 6748
rect 28252 7028 28308 7038
rect 27132 6692 27188 6702
rect 27580 6692 27636 6702
rect 27132 6690 27636 6692
rect 27132 6638 27134 6690
rect 27186 6638 27582 6690
rect 27634 6638 27636 6690
rect 27132 6636 27636 6638
rect 27132 6626 27188 6636
rect 27020 6412 27188 6468
rect 26460 5070 26462 5122
rect 26514 5070 26516 5122
rect 26348 4564 26404 4574
rect 26236 4562 26404 4564
rect 26236 4510 26350 4562
rect 26402 4510 26404 4562
rect 26236 4508 26404 4510
rect 26124 4470 26180 4508
rect 26348 4498 26404 4508
rect 26012 4340 26068 4350
rect 26012 4246 26068 4284
rect 26236 4228 26292 4238
rect 26236 4134 26292 4172
rect 25900 3556 25956 3566
rect 25900 3462 25956 3500
rect 25788 3266 25844 3276
rect 26124 3444 26180 3454
rect 25228 1138 25284 1148
rect 23996 924 24500 980
rect 23996 800 24052 924
rect 26124 800 26180 3388
rect 26348 3444 26404 3482
rect 26348 3378 26404 3388
rect 26460 2100 26516 5070
rect 26796 5180 26964 5236
rect 27020 6244 27076 6254
rect 26796 3388 26852 5180
rect 27020 5124 27076 6188
rect 27132 5906 27188 6412
rect 27132 5854 27134 5906
rect 27186 5854 27188 5906
rect 27132 5842 27188 5854
rect 27580 5908 27636 6636
rect 28252 6690 28308 6972
rect 28252 6638 28254 6690
rect 28306 6638 28308 6690
rect 28252 6626 28308 6638
rect 28140 6580 28196 6590
rect 28140 6486 28196 6524
rect 28028 6468 28084 6478
rect 28028 6374 28084 6412
rect 28140 5908 28196 5918
rect 27580 5906 28196 5908
rect 27580 5854 28142 5906
rect 28194 5854 28196 5906
rect 27580 5852 28196 5854
rect 28140 5842 28196 5852
rect 27468 5796 27524 5806
rect 27468 5346 27524 5740
rect 27468 5294 27470 5346
rect 27522 5294 27524 5346
rect 27468 5234 27524 5294
rect 27468 5182 27470 5234
rect 27522 5182 27524 5234
rect 27468 5170 27524 5182
rect 27916 5460 27972 5470
rect 27916 5234 27972 5404
rect 27916 5182 27918 5234
rect 27970 5182 27972 5234
rect 26684 3332 26852 3388
rect 26908 5068 27076 5124
rect 26684 3330 26740 3332
rect 26684 3278 26686 3330
rect 26738 3278 26740 3330
rect 26684 3266 26740 3278
rect 26460 2034 26516 2044
rect 26908 1316 26964 5068
rect 27916 5012 27972 5182
rect 28364 5124 28420 5134
rect 28364 5030 28420 5068
rect 27916 4946 27972 4956
rect 27020 4898 27076 4910
rect 28476 4900 28532 7532
rect 28588 7028 28644 7644
rect 28700 7634 28756 7644
rect 28924 7698 28980 7980
rect 28924 7646 28926 7698
rect 28978 7646 28980 7698
rect 28588 6962 28644 6972
rect 28924 6804 28980 7646
rect 29036 7586 29092 9324
rect 29484 9266 29540 9324
rect 29484 9214 29486 9266
rect 29538 9214 29540 9266
rect 29484 9156 29540 9214
rect 29484 9090 29540 9100
rect 29596 8372 29652 9660
rect 29708 9602 29764 9884
rect 29932 9826 29988 11004
rect 30716 10948 30772 13132
rect 30828 12292 30884 12302
rect 30828 12198 30884 12236
rect 30492 10892 30772 10948
rect 30492 10722 30548 10892
rect 30492 10670 30494 10722
rect 30546 10670 30548 10722
rect 30492 10658 30548 10670
rect 30604 10722 30660 10734
rect 30604 10670 30606 10722
rect 30658 10670 30660 10722
rect 30192 10220 30456 10230
rect 30248 10164 30296 10220
rect 30352 10164 30400 10220
rect 30192 10154 30456 10164
rect 29932 9774 29934 9826
rect 29986 9774 29988 9826
rect 30268 9940 30324 9950
rect 30604 9940 30660 10670
rect 30716 10612 30772 10892
rect 31052 11170 31108 11182
rect 31052 11118 31054 11170
rect 31106 11118 31108 11170
rect 30828 10836 30884 10846
rect 30828 10742 30884 10780
rect 31052 10836 31108 11118
rect 31052 10770 31108 10780
rect 31276 10612 31332 17948
rect 31612 17666 31668 19068
rect 31724 19058 31780 19068
rect 32172 19012 32228 19022
rect 32172 18918 32228 18956
rect 32172 18452 32228 18462
rect 31612 17614 31614 17666
rect 31666 17614 31668 17666
rect 31612 17602 31668 17614
rect 32060 18338 32116 18350
rect 32060 18286 32062 18338
rect 32114 18286 32116 18338
rect 31724 17554 31780 17566
rect 31724 17502 31726 17554
rect 31778 17502 31780 17554
rect 31724 16548 31780 17502
rect 31948 17108 32004 17118
rect 32060 17108 32116 18286
rect 32172 17778 32228 18396
rect 32284 18340 32340 18350
rect 32284 18246 32340 18284
rect 32172 17726 32174 17778
rect 32226 17726 32228 17778
rect 32172 17714 32228 17726
rect 32620 18226 32676 18238
rect 32620 18174 32622 18226
rect 32674 18174 32676 18226
rect 32508 17668 32564 17678
rect 32620 17668 32676 18174
rect 32508 17666 32676 17668
rect 32508 17614 32510 17666
rect 32562 17614 32676 17666
rect 32508 17612 32676 17614
rect 32508 17602 32564 17612
rect 32844 17556 32900 24556
rect 32956 22372 33012 22382
rect 33404 22372 33460 22382
rect 32956 22278 33012 22316
rect 33068 22370 33460 22372
rect 33068 22318 33406 22370
rect 33458 22318 33460 22370
rect 33068 22316 33460 22318
rect 32956 21812 33012 21822
rect 33068 21812 33124 22316
rect 33404 22306 33460 22316
rect 32956 21810 33124 21812
rect 32956 21758 32958 21810
rect 33010 21758 33124 21810
rect 32956 21756 33124 21758
rect 32956 21746 33012 21756
rect 33516 20188 33572 29932
rect 33964 30100 34020 30110
rect 33964 29650 34020 30044
rect 33964 29598 33966 29650
rect 34018 29598 34020 29650
rect 33964 29586 34020 29598
rect 34076 29988 34132 30268
rect 34412 30100 34468 30110
rect 34524 30100 34580 30268
rect 34748 30322 34804 30334
rect 34748 30270 34750 30322
rect 34802 30270 34804 30322
rect 34748 30212 34804 30270
rect 35420 30324 35476 30334
rect 35420 30230 35476 30268
rect 34748 30146 34804 30156
rect 35308 30212 35364 30222
rect 35308 30118 35364 30156
rect 34412 30098 34580 30100
rect 34412 30046 34414 30098
rect 34466 30046 34580 30098
rect 34412 30044 34580 30046
rect 34412 30034 34468 30044
rect 33628 29540 33684 29550
rect 33628 29446 33684 29484
rect 33740 29540 33796 29550
rect 33740 29538 33908 29540
rect 33740 29486 33742 29538
rect 33794 29486 33908 29538
rect 33740 29484 33908 29486
rect 33740 29474 33796 29484
rect 33740 28868 33796 28878
rect 33852 28868 33908 29484
rect 33740 28866 33908 28868
rect 33740 28814 33742 28866
rect 33794 28814 33908 28866
rect 33740 28812 33908 28814
rect 33740 28802 33796 28812
rect 33740 28644 33796 28654
rect 33628 28532 33684 28542
rect 33628 28438 33684 28476
rect 33740 28530 33796 28588
rect 33740 28478 33742 28530
rect 33794 28478 33796 28530
rect 33740 28466 33796 28478
rect 34076 28308 34132 29932
rect 34636 29988 34692 29998
rect 34636 29894 34692 29932
rect 35532 29986 35588 31054
rect 37100 31106 37156 31892
rect 37548 31890 37604 32396
rect 37660 32562 38164 32564
rect 37660 32510 38110 32562
rect 38162 32510 38164 32562
rect 37660 32508 38164 32510
rect 37660 32450 37716 32508
rect 38108 32498 38164 32508
rect 38780 32562 38836 32574
rect 38780 32510 38782 32562
rect 38834 32510 38836 32562
rect 37660 32398 37662 32450
rect 37714 32398 37716 32450
rect 37660 32386 37716 32398
rect 38108 32228 38164 32238
rect 37772 32004 37828 32042
rect 37772 31938 37828 31948
rect 37548 31838 37550 31890
rect 37602 31838 37604 31890
rect 37548 31826 37604 31838
rect 38108 31890 38164 32172
rect 38780 32228 38836 32510
rect 42252 32452 42308 32462
rect 38780 32162 38836 32172
rect 41804 32450 42308 32452
rect 41804 32398 42254 32450
rect 42306 32398 42308 32450
rect 41804 32396 42308 32398
rect 38108 31838 38110 31890
rect 38162 31838 38164 31890
rect 38108 31826 38164 31838
rect 40124 31892 40180 31902
rect 40124 31890 40292 31892
rect 40124 31838 40126 31890
rect 40178 31838 40292 31890
rect 40124 31836 40292 31838
rect 40124 31826 40180 31836
rect 39676 31778 39732 31790
rect 39676 31726 39678 31778
rect 39730 31726 39732 31778
rect 37100 31054 37102 31106
rect 37154 31054 37156 31106
rect 37100 31042 37156 31054
rect 39004 31556 39060 31566
rect 39676 31556 39732 31726
rect 39004 31554 39732 31556
rect 39004 31502 39006 31554
rect 39058 31502 39732 31554
rect 39004 31500 39732 31502
rect 36428 30994 36484 31006
rect 36428 30942 36430 30994
rect 36482 30942 36484 30994
rect 36428 30660 36484 30942
rect 37884 30772 37940 30782
rect 36484 30604 36708 30660
rect 36428 30594 36484 30604
rect 35980 30212 36036 30222
rect 36316 30212 36372 30222
rect 35980 30210 36372 30212
rect 35980 30158 35982 30210
rect 36034 30158 36318 30210
rect 36370 30158 36372 30210
rect 35980 30156 36372 30158
rect 35980 30146 36036 30156
rect 36316 30146 36372 30156
rect 36652 30212 36708 30604
rect 36652 30080 36708 30156
rect 37436 30212 37492 30222
rect 37436 30118 37492 30156
rect 35532 29934 35534 29986
rect 35586 29934 35588 29986
rect 35532 29316 35588 29934
rect 36092 29988 36148 29998
rect 36092 29650 36148 29932
rect 36540 29988 36596 29998
rect 36540 29894 36596 29932
rect 36092 29598 36094 29650
rect 36146 29598 36148 29650
rect 36092 29586 36148 29598
rect 37884 29538 37940 30716
rect 39004 30100 39060 31500
rect 39852 31388 40116 31398
rect 39908 31332 39956 31388
rect 40012 31332 40060 31388
rect 39852 31322 40116 31332
rect 39340 31108 39396 31118
rect 39340 30994 39396 31052
rect 39340 30942 39342 30994
rect 39394 30942 39396 30994
rect 39116 30884 39172 30894
rect 39116 30324 39172 30828
rect 39340 30772 39396 30942
rect 39676 30996 39732 31006
rect 39676 30882 39732 30940
rect 39676 30830 39678 30882
rect 39730 30830 39732 30882
rect 39676 30818 39732 30830
rect 40236 30884 40292 31836
rect 41804 31890 41860 32396
rect 42252 32386 42308 32396
rect 41804 31838 41806 31890
rect 41858 31838 41860 31890
rect 41804 31826 41860 31838
rect 43932 31892 43988 33180
rect 44380 33012 44436 36204
rect 45052 36258 45108 36270
rect 45052 36206 45054 36258
rect 45106 36206 45108 36258
rect 44940 35698 44996 35710
rect 44940 35646 44942 35698
rect 44994 35646 44996 35698
rect 44716 35252 44772 35262
rect 44716 35026 44772 35196
rect 44716 34974 44718 35026
rect 44770 34974 44772 35026
rect 44716 34962 44772 34974
rect 44940 34916 44996 35646
rect 44940 34850 44996 34860
rect 45052 34244 45108 36206
rect 45276 36260 45332 36270
rect 45276 36166 45332 36204
rect 45388 36258 45444 36270
rect 45388 36206 45390 36258
rect 45442 36206 45444 36258
rect 45388 35924 45444 36206
rect 45500 36258 45556 36270
rect 45500 36206 45502 36258
rect 45554 36206 45556 36258
rect 45500 36148 45556 36206
rect 45500 36082 45556 36092
rect 47180 36260 47236 36270
rect 45388 35868 46116 35924
rect 45612 35700 45668 35710
rect 45612 35606 45668 35644
rect 46060 35698 46116 35868
rect 46060 35646 46062 35698
rect 46114 35646 46116 35698
rect 46060 35634 46116 35646
rect 47180 35700 47236 36204
rect 46508 35586 46564 35598
rect 46508 35534 46510 35586
rect 46562 35534 46564 35586
rect 46172 35476 46228 35486
rect 46172 35026 46228 35420
rect 46508 35252 46564 35534
rect 46508 35186 46564 35196
rect 47180 35138 47236 35644
rect 47180 35086 47182 35138
rect 47234 35086 47236 35138
rect 47180 35074 47236 35086
rect 47628 36260 47684 36428
rect 49196 36482 49924 36484
rect 49196 36430 49870 36482
rect 49922 36430 49924 36482
rect 49196 36428 49924 36430
rect 47964 36260 48020 36270
rect 47628 36258 48020 36260
rect 47628 36206 47966 36258
rect 48018 36206 48020 36258
rect 47628 36204 48020 36206
rect 46172 34974 46174 35026
rect 46226 34974 46228 35026
rect 45052 34178 45108 34188
rect 45388 34916 45444 34926
rect 45388 34690 45444 34860
rect 46172 34916 46228 34974
rect 46172 34850 46228 34860
rect 47180 34916 47236 34926
rect 46620 34804 46676 34814
rect 46620 34710 46676 34748
rect 45388 34638 45390 34690
rect 45442 34638 45444 34690
rect 44716 33234 44772 33246
rect 44716 33182 44718 33234
rect 44770 33182 44772 33234
rect 44716 33124 44772 33182
rect 44716 33058 44772 33068
rect 44044 31892 44100 31902
rect 43932 31890 44100 31892
rect 43932 31838 44046 31890
rect 44098 31838 44100 31890
rect 43932 31836 44100 31838
rect 44044 31826 44100 31836
rect 40460 31780 40516 31790
rect 40460 31108 40516 31724
rect 41020 31780 41076 31790
rect 41020 31686 41076 31724
rect 43596 31778 43652 31790
rect 43596 31726 43598 31778
rect 43650 31726 43652 31778
rect 40460 30994 40516 31052
rect 42028 31108 42084 31118
rect 42028 31014 42084 31052
rect 43596 31108 43652 31726
rect 43596 31014 43652 31052
rect 43820 31778 43876 31790
rect 43820 31726 43822 31778
rect 43874 31726 43876 31778
rect 40460 30942 40462 30994
rect 40514 30942 40516 30994
rect 40460 30930 40516 30942
rect 40796 30996 40852 31006
rect 41580 30996 41636 31006
rect 41804 30996 41860 31006
rect 40796 30994 41636 30996
rect 40796 30942 40798 30994
rect 40850 30942 41582 30994
rect 41634 30942 41636 30994
rect 40796 30940 41636 30942
rect 40796 30930 40852 30940
rect 41580 30930 41636 30940
rect 41692 30994 41860 30996
rect 41692 30942 41806 30994
rect 41858 30942 41860 30994
rect 41692 30940 41860 30942
rect 40236 30790 40292 30828
rect 39340 30706 39396 30716
rect 39116 30258 39172 30268
rect 39004 30034 39060 30044
rect 41692 30100 41748 30940
rect 41804 30930 41860 30940
rect 42140 30996 42196 31006
rect 43820 30996 43876 31726
rect 44380 31444 44436 32956
rect 44380 31378 44436 31388
rect 44492 32676 44548 32686
rect 45388 32676 45444 34638
rect 47180 33684 47236 34860
rect 47516 34804 47572 34814
rect 47516 34710 47572 34748
rect 47180 33460 47236 33628
rect 47292 33460 47348 33470
rect 47180 33458 47348 33460
rect 47180 33406 47294 33458
rect 47346 33406 47348 33458
rect 47180 33404 47348 33406
rect 47292 33394 47348 33404
rect 45612 33348 45668 33358
rect 45500 33236 45556 33246
rect 45500 33142 45556 33180
rect 45612 33234 45668 33292
rect 45612 33182 45614 33234
rect 45666 33182 45668 33234
rect 45612 33170 45668 33182
rect 45836 33236 45892 33246
rect 45836 33142 45892 33180
rect 46060 33236 46116 33246
rect 47628 33236 47684 36204
rect 47964 36194 48020 36204
rect 47852 36036 47908 36046
rect 47852 35698 47908 35980
rect 48300 36036 48356 36046
rect 47852 35646 47854 35698
rect 47906 35646 47908 35698
rect 47852 35634 47908 35646
rect 48076 35700 48132 35710
rect 48076 35606 48132 35644
rect 48188 35252 48244 35262
rect 48188 35138 48244 35196
rect 48188 35086 48190 35138
rect 48242 35086 48244 35138
rect 48188 35074 48244 35086
rect 48300 35138 48356 35980
rect 48300 35086 48302 35138
rect 48354 35086 48356 35138
rect 48300 35074 48356 35086
rect 48524 35700 48580 35710
rect 48524 35138 48580 35644
rect 48524 35086 48526 35138
rect 48578 35086 48580 35138
rect 48524 35074 48580 35086
rect 48748 35586 48804 35598
rect 48748 35534 48750 35586
rect 48802 35534 48804 35586
rect 48748 34916 48804 35534
rect 48748 34850 48804 34860
rect 47740 34804 47796 34814
rect 47740 33460 47796 34748
rect 48636 34804 48692 34814
rect 48636 34710 48692 34748
rect 49196 34690 49252 36428
rect 49868 36418 49924 36428
rect 51884 36482 51940 36494
rect 51884 36430 51886 36482
rect 51938 36430 51940 36482
rect 49756 36036 49812 36046
rect 49756 35922 49812 35980
rect 49756 35870 49758 35922
rect 49810 35870 49812 35922
rect 49756 35858 49812 35870
rect 51436 35698 51492 35710
rect 51436 35646 51438 35698
rect 51490 35646 51492 35698
rect 50540 35588 50596 35598
rect 51436 35588 51492 35646
rect 50540 35586 51492 35588
rect 50540 35534 50542 35586
rect 50594 35534 51492 35586
rect 50540 35532 51492 35534
rect 51884 35588 51940 36430
rect 52220 35924 52276 36764
rect 53452 36596 53508 39200
rect 55916 39060 55972 39200
rect 56252 39060 56308 39228
rect 55916 39004 56308 39060
rect 53452 36530 53508 36540
rect 53676 37716 53732 37726
rect 53676 36484 53732 37660
rect 54348 36596 54404 36606
rect 54348 36502 54404 36540
rect 56812 36594 56868 39228
rect 58352 39200 58464 40000
rect 60816 39200 60928 40000
rect 61180 39228 61796 39284
rect 56812 36542 56814 36594
rect 56866 36542 56868 36594
rect 56812 36530 56868 36542
rect 57708 37492 57764 37502
rect 53564 36482 53732 36484
rect 53564 36430 53678 36482
rect 53730 36430 53732 36482
rect 53564 36428 53732 36430
rect 52108 35812 52164 35822
rect 52108 35718 52164 35756
rect 49532 35476 49588 35486
rect 49308 35474 49588 35476
rect 49308 35422 49534 35474
rect 49586 35422 49588 35474
rect 49308 35420 49588 35422
rect 49308 35252 49364 35420
rect 49532 35410 49588 35420
rect 49868 35474 49924 35486
rect 49868 35422 49870 35474
rect 49922 35422 49924 35474
rect 49512 35308 49776 35318
rect 49568 35252 49616 35308
rect 49672 35252 49720 35308
rect 49512 35242 49776 35252
rect 49308 35186 49364 35196
rect 49756 34804 49812 34814
rect 49756 34710 49812 34748
rect 49196 34638 49198 34690
rect 49250 34638 49252 34690
rect 48412 33684 48468 33694
rect 47740 33458 48244 33460
rect 47740 33406 47742 33458
rect 47794 33406 48244 33458
rect 47740 33404 48244 33406
rect 47740 33394 47796 33404
rect 48188 33346 48244 33404
rect 48188 33294 48190 33346
rect 48242 33294 48244 33346
rect 48188 33282 48244 33294
rect 48412 33346 48468 33628
rect 48412 33294 48414 33346
rect 48466 33294 48468 33346
rect 48412 33282 48468 33294
rect 45388 32620 45556 32676
rect 44492 31332 44548 32620
rect 44492 31266 44548 31276
rect 45388 32450 45444 32462
rect 45388 32398 45390 32450
rect 45442 32398 45444 32450
rect 45388 31780 45444 32398
rect 44156 31220 44212 31230
rect 44156 31126 44212 31164
rect 42140 30902 42196 30940
rect 43708 30994 43876 30996
rect 43708 30942 43822 30994
rect 43874 30942 43876 30994
rect 43708 30940 43876 30942
rect 41692 30006 41748 30044
rect 42140 30772 42196 30782
rect 40908 29988 40964 29998
rect 39852 29820 40116 29830
rect 39908 29764 39956 29820
rect 40012 29764 40060 29820
rect 39852 29754 40116 29764
rect 40460 29652 40516 29662
rect 40460 29558 40516 29596
rect 37884 29486 37886 29538
rect 37938 29486 37940 29538
rect 37884 29474 37940 29486
rect 37324 29426 37380 29438
rect 40124 29428 40180 29438
rect 37324 29374 37326 29426
rect 37378 29374 37380 29426
rect 35532 29250 35588 29260
rect 37100 29314 37156 29326
rect 37100 29262 37102 29314
rect 37154 29262 37156 29314
rect 35756 29204 35812 29214
rect 34300 28644 34356 28654
rect 34300 28550 34356 28588
rect 33628 28252 34132 28308
rect 35196 28420 35252 28430
rect 33628 24612 33684 28252
rect 35084 27748 35140 27758
rect 35196 27748 35252 28364
rect 35644 28420 35700 28430
rect 35644 28326 35700 28364
rect 35756 28084 35812 29148
rect 36876 28644 36932 28654
rect 36876 28550 36932 28588
rect 36540 28530 36596 28542
rect 36540 28478 36542 28530
rect 36594 28478 36596 28530
rect 35756 28018 35812 28028
rect 36092 28420 36148 28430
rect 35084 27746 35252 27748
rect 35084 27694 35086 27746
rect 35138 27694 35252 27746
rect 35084 27692 35252 27694
rect 35084 27682 35140 27692
rect 34636 27188 34692 27198
rect 34636 27094 34692 27132
rect 34300 27074 34356 27086
rect 34300 27022 34302 27074
rect 34354 27022 34356 27074
rect 33628 24546 33684 24556
rect 33740 26850 33796 26862
rect 33740 26798 33742 26850
rect 33794 26798 33796 26850
rect 33740 26180 33796 26798
rect 34300 26516 34356 27022
rect 34860 27074 34916 27086
rect 34860 27022 34862 27074
rect 34914 27022 34916 27074
rect 34300 26450 34356 26460
rect 34412 26962 34468 26974
rect 34412 26910 34414 26962
rect 34466 26910 34468 26962
rect 34412 26292 34468 26910
rect 34748 26292 34804 26302
rect 34188 26290 34804 26292
rect 34188 26238 34750 26290
rect 34802 26238 34804 26290
rect 34188 26236 34804 26238
rect 33852 26180 33908 26190
rect 34188 26180 34244 26236
rect 34748 26226 34804 26236
rect 33740 26178 34244 26180
rect 33740 26126 33854 26178
rect 33906 26126 34244 26178
rect 33740 26124 34244 26126
rect 34860 26180 34916 27022
rect 34972 26180 35028 26190
rect 34860 26178 35028 26180
rect 34860 26126 34974 26178
rect 35026 26126 35028 26178
rect 34860 26124 35028 26126
rect 32844 17490 32900 17500
rect 33180 20132 33236 20142
rect 32844 17332 32900 17342
rect 32732 17220 32788 17230
rect 32060 17052 32340 17108
rect 31836 16996 31892 17006
rect 31836 16882 31892 16940
rect 31836 16830 31838 16882
rect 31890 16830 31892 16882
rect 31836 16818 31892 16830
rect 31724 16492 31892 16548
rect 31724 16324 31780 16334
rect 31724 15876 31780 16268
rect 31836 15876 31892 16492
rect 31948 16100 32004 17052
rect 32060 16882 32116 16894
rect 32060 16830 32062 16882
rect 32114 16830 32116 16882
rect 32060 16212 32116 16830
rect 32172 16212 32228 16222
rect 32060 16210 32228 16212
rect 32060 16158 32174 16210
rect 32226 16158 32228 16210
rect 32060 16156 32228 16158
rect 31948 15968 32004 16044
rect 32172 16100 32228 16156
rect 32172 16034 32228 16044
rect 32060 15988 32116 15998
rect 32060 15876 32116 15932
rect 31836 15820 32116 15876
rect 31724 15538 31780 15820
rect 32284 15764 32340 17052
rect 32732 17106 32788 17164
rect 32732 17054 32734 17106
rect 32786 17054 32788 17106
rect 32508 16996 32564 17006
rect 32508 16902 32564 16940
rect 32732 16660 32788 17054
rect 32844 16994 32900 17276
rect 32844 16942 32846 16994
rect 32898 16942 32900 16994
rect 32844 16884 32900 16942
rect 32844 16818 32900 16828
rect 32732 16594 32788 16604
rect 32396 15988 32452 15998
rect 32620 15988 32676 15998
rect 32452 15932 32564 15988
rect 32396 15922 32452 15932
rect 32508 15876 32564 15932
rect 32620 15894 32676 15932
rect 31724 15486 31726 15538
rect 31778 15486 31780 15538
rect 31724 15474 31780 15486
rect 31948 15708 32340 15764
rect 32396 15764 32452 15774
rect 31948 15538 32004 15708
rect 31948 15486 31950 15538
rect 32002 15486 32004 15538
rect 31948 15428 32004 15486
rect 31948 15362 32004 15372
rect 31836 15316 31892 15326
rect 31836 15222 31892 15260
rect 32396 15314 32452 15708
rect 32396 15262 32398 15314
rect 32450 15262 32452 15314
rect 32396 15250 32452 15262
rect 32172 15204 32228 15214
rect 32172 15110 32228 15148
rect 32396 14756 32452 14766
rect 32396 14530 32452 14700
rect 32508 14642 32564 15820
rect 32508 14590 32510 14642
rect 32562 14590 32564 14642
rect 32508 14578 32564 14590
rect 32396 14478 32398 14530
rect 32450 14478 32452 14530
rect 32396 14466 32452 14478
rect 32620 13748 32676 13758
rect 32172 13074 32228 13086
rect 32172 13022 32174 13074
rect 32226 13022 32228 13074
rect 31500 12740 31556 12750
rect 31500 12180 31556 12684
rect 32172 12740 32228 13022
rect 32620 12962 32676 13692
rect 32620 12910 32622 12962
rect 32674 12910 32676 12962
rect 32620 12898 32676 12910
rect 32732 13524 32788 13534
rect 32172 12674 32228 12684
rect 31500 12114 31556 12124
rect 31836 10836 31892 10846
rect 30716 10556 30996 10612
rect 30324 9884 30660 9940
rect 30940 9940 30996 10556
rect 31276 10546 31332 10556
rect 31500 10610 31556 10622
rect 31500 10558 31502 10610
rect 31554 10558 31556 10610
rect 30268 9808 30324 9884
rect 30940 9808 30996 9884
rect 29932 9762 29988 9774
rect 29708 9550 29710 9602
rect 29762 9550 29764 9602
rect 29708 9268 29764 9550
rect 29708 9202 29764 9212
rect 30828 9268 30884 9278
rect 31388 9268 31444 9278
rect 31500 9268 31556 10558
rect 31836 10498 31892 10780
rect 31836 10446 31838 10498
rect 31890 10446 31892 10498
rect 31836 10434 31892 10446
rect 32284 10724 32340 10734
rect 30828 9266 31556 9268
rect 30828 9214 30830 9266
rect 30882 9214 31390 9266
rect 31442 9214 31556 9266
rect 30828 9212 31556 9214
rect 32284 9938 32340 10668
rect 32396 10612 32452 10622
rect 32396 10518 32452 10556
rect 32284 9886 32286 9938
rect 32338 9886 32340 9938
rect 32284 9268 32340 9886
rect 32732 9716 32788 13468
rect 32844 12628 32900 12638
rect 32844 10500 32900 12572
rect 33180 12292 33236 20076
rect 33404 20132 33572 20188
rect 33628 23938 33684 23950
rect 33628 23886 33630 23938
rect 33682 23886 33684 23938
rect 33628 23716 33684 23886
rect 33292 17442 33348 17454
rect 33292 17390 33294 17442
rect 33346 17390 33348 17442
rect 33292 17220 33348 17390
rect 33292 17154 33348 17164
rect 33404 13860 33460 20132
rect 33516 19572 33572 19582
rect 33516 19012 33572 19516
rect 33516 18946 33572 18956
rect 33628 18452 33684 23660
rect 33740 22596 33796 26124
rect 33852 26114 33908 26124
rect 34300 26068 34356 26078
rect 33852 25506 33908 25518
rect 33852 25454 33854 25506
rect 33906 25454 33908 25506
rect 33852 25396 33908 25454
rect 34300 25508 34356 26012
rect 34748 25620 34804 25630
rect 34860 25620 34916 26124
rect 34972 26114 35028 26124
rect 34748 25618 34916 25620
rect 34748 25566 34750 25618
rect 34802 25566 34916 25618
rect 34748 25564 34916 25566
rect 34748 25554 34804 25564
rect 34300 25376 34356 25452
rect 33852 25330 33908 25340
rect 33852 24724 33908 24734
rect 33852 24630 33908 24668
rect 34076 24724 34132 24734
rect 34076 24050 34132 24668
rect 34524 24724 34580 24734
rect 34524 24630 34580 24668
rect 34636 24612 34692 24622
rect 34636 24518 34692 24556
rect 34076 23998 34078 24050
rect 34130 23998 34132 24050
rect 34076 23986 34132 23998
rect 33964 23940 34020 23950
rect 33964 23846 34020 23884
rect 34636 23940 34692 23950
rect 34636 23266 34692 23884
rect 34748 23716 34804 23726
rect 34748 23492 34804 23660
rect 34972 23716 35028 23726
rect 34972 23622 35028 23660
rect 34748 23436 35140 23492
rect 35084 23378 35140 23436
rect 35084 23326 35086 23378
rect 35138 23326 35140 23378
rect 35084 23314 35140 23326
rect 34636 23214 34638 23266
rect 34690 23214 34692 23266
rect 34636 23202 34692 23214
rect 34076 23156 34132 23166
rect 33740 22530 33796 22540
rect 33852 23100 34076 23156
rect 33852 22370 33908 23100
rect 34076 23062 34132 23100
rect 34188 23042 34244 23054
rect 34188 22990 34190 23042
rect 34242 22990 34244 23042
rect 33852 22318 33854 22370
rect 33906 22318 33908 22370
rect 33852 22306 33908 22318
rect 34076 22372 34132 22382
rect 34188 22372 34244 22990
rect 34132 22316 34244 22372
rect 34076 22240 34132 22316
rect 33964 22146 34020 22158
rect 33964 22094 33966 22146
rect 34018 22094 34020 22146
rect 33964 21700 34020 22094
rect 33964 21634 34020 21644
rect 34972 21028 35028 21038
rect 34972 20934 35028 20972
rect 33852 20804 33908 20814
rect 34412 20804 34468 20814
rect 33740 20802 34468 20804
rect 33740 20750 33854 20802
rect 33906 20750 34414 20802
rect 34466 20750 34468 20802
rect 33740 20748 34468 20750
rect 33740 20018 33796 20748
rect 33852 20738 33908 20748
rect 34412 20738 34468 20748
rect 34636 20802 34692 20814
rect 34636 20750 34638 20802
rect 34690 20750 34692 20802
rect 33740 19966 33742 20018
rect 33794 19966 33796 20018
rect 33740 19684 33796 19966
rect 34300 19908 34356 19918
rect 33740 19618 33796 19628
rect 33852 19906 34356 19908
rect 33852 19854 34302 19906
rect 34354 19854 34356 19906
rect 33852 19852 34356 19854
rect 33852 19234 33908 19852
rect 34300 19842 34356 19852
rect 34636 19908 34692 20750
rect 35196 20132 35252 27692
rect 35532 27748 35588 27758
rect 35532 27654 35588 27692
rect 36092 27748 36148 28364
rect 36428 28308 36484 28318
rect 36540 28308 36596 28478
rect 36652 28420 36708 28430
rect 36652 28326 36708 28364
rect 37100 28420 37156 29262
rect 36484 28252 36596 28308
rect 36092 27682 36148 27692
rect 36316 27858 36372 27870
rect 36316 27806 36318 27858
rect 36370 27806 36372 27858
rect 36316 27748 36372 27806
rect 36316 27682 36372 27692
rect 36428 27746 36484 28252
rect 36428 27694 36430 27746
rect 36482 27694 36484 27746
rect 36428 27682 36484 27694
rect 36316 27300 36372 27310
rect 36316 27206 36372 27244
rect 37100 27300 37156 28364
rect 37212 27972 37268 27982
rect 37324 27972 37380 29374
rect 39676 29426 40180 29428
rect 39676 29374 40126 29426
rect 40178 29374 40180 29426
rect 39676 29372 40180 29374
rect 37996 29316 38052 29326
rect 37436 28644 37492 28654
rect 37436 28550 37492 28588
rect 37996 28530 38052 29260
rect 37996 28478 37998 28530
rect 38050 28478 38052 28530
rect 37996 28466 38052 28478
rect 38556 29314 38612 29326
rect 38556 29262 38558 29314
rect 38610 29262 38612 29314
rect 38556 29204 38612 29262
rect 39116 29316 39172 29326
rect 39116 29222 39172 29260
rect 39676 29314 39732 29372
rect 40124 29362 40180 29372
rect 40572 29428 40628 29438
rect 40572 29334 40628 29372
rect 40684 29426 40740 29438
rect 40684 29374 40686 29426
rect 40738 29374 40740 29426
rect 39676 29262 39678 29314
rect 39730 29262 39732 29314
rect 39676 29250 39732 29262
rect 37884 28418 37940 28430
rect 37884 28366 37886 28418
rect 37938 28366 37940 28418
rect 37884 27972 37940 28366
rect 38108 28420 38164 28430
rect 38108 28326 38164 28364
rect 38556 28196 38612 29148
rect 39340 29204 39396 29214
rect 39340 28756 39396 29148
rect 40572 28868 40628 28878
rect 40684 28868 40740 29374
rect 40572 28866 40740 28868
rect 40572 28814 40574 28866
rect 40626 28814 40740 28866
rect 40572 28812 40740 28814
rect 40796 29428 40852 29438
rect 40572 28802 40628 28812
rect 39340 28690 39396 28700
rect 40012 28756 40068 28766
rect 40012 28662 40068 28700
rect 40236 28532 40292 28542
rect 37212 27970 37940 27972
rect 37212 27918 37214 27970
rect 37266 27918 37940 27970
rect 37212 27916 37940 27918
rect 37996 28140 38612 28196
rect 39852 28252 40116 28262
rect 39908 28196 39956 28252
rect 40012 28196 40060 28252
rect 39852 28186 40116 28196
rect 37212 27906 37268 27916
rect 37100 27234 37156 27244
rect 35644 27186 35700 27198
rect 35644 27134 35646 27186
rect 35698 27134 35700 27186
rect 35420 26404 35476 26414
rect 35644 26404 35700 27134
rect 35420 26402 35700 26404
rect 35420 26350 35422 26402
rect 35474 26350 35700 26402
rect 35420 26348 35700 26350
rect 35420 26338 35476 26348
rect 35644 26292 35700 26348
rect 35644 26226 35700 26236
rect 35980 27074 36036 27086
rect 35980 27022 35982 27074
rect 36034 27022 36036 27074
rect 35980 26180 36036 27022
rect 36652 26852 36708 26862
rect 36540 26516 36596 26526
rect 36540 26422 36596 26460
rect 36204 26292 36260 26302
rect 36204 26198 36260 26236
rect 35980 26086 36036 26124
rect 35420 24836 35476 24846
rect 35420 24742 35476 24780
rect 35308 24724 35364 24734
rect 35308 24630 35364 24668
rect 35420 24498 35476 24510
rect 35420 24446 35422 24498
rect 35474 24446 35476 24498
rect 35420 23938 35476 24446
rect 35420 23886 35422 23938
rect 35474 23886 35476 23938
rect 35420 23874 35476 23886
rect 35756 24276 35812 24286
rect 35756 23938 35812 24220
rect 35756 23886 35758 23938
rect 35810 23886 35812 23938
rect 35756 23874 35812 23886
rect 35532 23716 35588 23726
rect 35532 23622 35588 23660
rect 36204 23044 36260 23054
rect 36204 22036 36260 22988
rect 36652 22260 36708 26796
rect 37772 24836 37828 24846
rect 37996 24836 38052 28140
rect 40124 27858 40180 27870
rect 40124 27806 40126 27858
rect 40178 27806 40180 27858
rect 39340 27746 39396 27758
rect 39340 27694 39342 27746
rect 39394 27694 39396 27746
rect 39228 27300 39284 27310
rect 39228 27186 39284 27244
rect 39228 27134 39230 27186
rect 39282 27134 39284 27186
rect 39228 27122 39284 27134
rect 38556 27076 38612 27086
rect 38556 26982 38612 27020
rect 39004 27076 39060 27086
rect 38668 26740 38724 26750
rect 38668 26402 38724 26684
rect 38668 26350 38670 26402
rect 38722 26350 38724 26402
rect 38668 26338 38724 26350
rect 38332 26292 38388 26330
rect 38332 26226 38388 26236
rect 38332 26068 38388 26078
rect 38332 25974 38388 26012
rect 38668 25844 38724 25854
rect 38668 25618 38724 25788
rect 38668 25566 38670 25618
rect 38722 25566 38724 25618
rect 38668 25554 38724 25566
rect 39004 25620 39060 27020
rect 39340 26908 39396 27694
rect 39900 27746 39956 27758
rect 39900 27694 39902 27746
rect 39954 27694 39956 27746
rect 39900 27636 39956 27694
rect 39676 27300 39732 27310
rect 39676 27206 39732 27244
rect 39900 27188 39956 27580
rect 40124 27748 40180 27806
rect 40124 27300 40180 27692
rect 40124 27234 40180 27244
rect 39900 27122 39956 27132
rect 39788 27076 39844 27086
rect 39788 26982 39844 27020
rect 39900 26962 39956 26974
rect 39900 26910 39902 26962
rect 39954 26910 39956 26962
rect 39116 26850 39172 26862
rect 39340 26852 39508 26908
rect 39116 26798 39118 26850
rect 39170 26798 39172 26850
rect 39116 26740 39172 26798
rect 39116 26674 39172 26684
rect 39452 26628 39508 26852
rect 39676 26852 39732 26862
rect 39564 26628 39620 26638
rect 39452 26572 39564 26628
rect 39452 26180 39508 26190
rect 39116 25620 39172 25630
rect 39004 25618 39172 25620
rect 39004 25566 39118 25618
rect 39170 25566 39172 25618
rect 39004 25564 39172 25566
rect 39116 25508 39172 25564
rect 39116 25442 39172 25452
rect 39340 25508 39396 25518
rect 38108 25284 38164 25294
rect 39228 25284 39284 25294
rect 38108 25282 38276 25284
rect 38108 25230 38110 25282
rect 38162 25230 38276 25282
rect 38108 25228 38276 25230
rect 38108 25218 38164 25228
rect 37772 24834 38052 24836
rect 37772 24782 37774 24834
rect 37826 24782 38052 24834
rect 37772 24780 38052 24782
rect 37772 24770 37828 24780
rect 37100 24722 37156 24734
rect 37100 24670 37102 24722
rect 37154 24670 37156 24722
rect 37100 24612 37156 24670
rect 37100 24546 37156 24556
rect 37660 24722 37716 24734
rect 37660 24670 37662 24722
rect 37714 24670 37716 24722
rect 37660 24052 37716 24670
rect 37996 24612 38052 24622
rect 37660 23996 37940 24052
rect 36876 23716 36932 23726
rect 36764 23154 36820 23166
rect 36764 23102 36766 23154
rect 36818 23102 36820 23154
rect 36764 23044 36820 23102
rect 36764 22978 36820 22988
rect 36540 22204 36708 22260
rect 36428 22148 36484 22158
rect 35756 21700 35812 21710
rect 35756 20802 35812 21644
rect 36092 21586 36148 21598
rect 36092 21534 36094 21586
rect 36146 21534 36148 21586
rect 36092 20916 36148 21534
rect 35756 20750 35758 20802
rect 35810 20750 35812 20802
rect 35756 20738 35812 20750
rect 35980 20914 36148 20916
rect 35980 20862 36094 20914
rect 36146 20862 36148 20914
rect 35980 20860 36148 20862
rect 35196 20066 35252 20076
rect 35868 20580 35924 20590
rect 35308 20018 35364 20030
rect 35308 19966 35310 20018
rect 35362 19966 35364 20018
rect 34636 19842 34692 19852
rect 35196 19908 35252 19918
rect 34412 19794 34468 19806
rect 34412 19742 34414 19794
rect 34466 19742 34468 19794
rect 33852 19182 33854 19234
rect 33906 19182 33908 19234
rect 33852 18676 33908 19182
rect 34076 19236 34132 19246
rect 34076 19142 34132 19180
rect 33852 18610 33908 18620
rect 34412 18564 34468 19742
rect 35196 19348 35252 19852
rect 35308 19684 35364 19966
rect 35308 19618 35364 19628
rect 35532 19684 35588 19694
rect 35308 19348 35364 19358
rect 35196 19346 35364 19348
rect 35196 19294 35310 19346
rect 35362 19294 35364 19346
rect 35196 19292 35364 19294
rect 35308 19282 35364 19292
rect 34636 19236 34692 19246
rect 34636 18674 34692 19180
rect 34748 19124 34804 19134
rect 34748 19030 34804 19068
rect 34636 18622 34638 18674
rect 34690 18622 34692 18674
rect 34636 18610 34692 18622
rect 34524 18564 34580 18574
rect 34412 18562 34580 18564
rect 34412 18510 34526 18562
rect 34578 18510 34580 18562
rect 34412 18508 34580 18510
rect 34524 18498 34580 18508
rect 34748 18564 34804 18574
rect 33628 18396 33796 18452
rect 33628 18228 33684 18238
rect 33628 17780 33684 18172
rect 33628 17648 33684 17724
rect 33516 17332 33572 17342
rect 33516 17106 33572 17276
rect 33516 17054 33518 17106
rect 33570 17054 33572 17106
rect 33516 17042 33572 17054
rect 33740 16100 33796 18396
rect 34748 18228 34804 18508
rect 34860 18452 34916 18462
rect 35196 18452 35252 18462
rect 34860 18450 35252 18452
rect 34860 18398 34862 18450
rect 34914 18398 35198 18450
rect 35250 18398 35252 18450
rect 34860 18396 35252 18398
rect 34860 18386 34916 18396
rect 35196 18386 35252 18396
rect 34748 18172 34916 18228
rect 34188 18116 34244 18126
rect 34188 17778 34244 18060
rect 34188 17726 34190 17778
rect 34242 17726 34244 17778
rect 34188 17714 34244 17726
rect 34524 17780 34580 17790
rect 34524 17686 34580 17724
rect 33852 16212 33908 16222
rect 33852 16210 34244 16212
rect 33852 16158 33854 16210
rect 33906 16158 34244 16210
rect 33852 16156 34244 16158
rect 33852 16146 33908 16156
rect 33628 16044 33796 16100
rect 33516 15988 33572 15998
rect 33516 14530 33572 15932
rect 33516 14478 33518 14530
rect 33570 14478 33572 14530
rect 33516 14466 33572 14478
rect 33628 14532 33684 16044
rect 33740 15876 33796 15886
rect 33740 15782 33796 15820
rect 34188 15538 34244 16156
rect 34412 15988 34468 15998
rect 34412 15894 34468 15932
rect 34524 15876 34580 15886
rect 34524 15782 34580 15820
rect 34748 15874 34804 15886
rect 34748 15822 34750 15874
rect 34802 15822 34804 15874
rect 34188 15486 34190 15538
rect 34242 15486 34244 15538
rect 34188 15474 34244 15486
rect 34300 15764 34356 15774
rect 34300 15538 34356 15708
rect 34300 15486 34302 15538
rect 34354 15486 34356 15538
rect 34300 15474 34356 15486
rect 34412 15314 34468 15326
rect 34412 15262 34414 15314
rect 34466 15262 34468 15314
rect 33628 14466 33684 14476
rect 33852 15092 33908 15102
rect 33404 13794 33460 13804
rect 33180 12226 33236 12236
rect 33404 12068 33460 12078
rect 32956 10724 33012 10734
rect 32956 10722 33348 10724
rect 32956 10670 32958 10722
rect 33010 10670 33348 10722
rect 32956 10668 33348 10670
rect 32956 10658 33012 10668
rect 32844 10434 32900 10444
rect 33180 10500 33236 10510
rect 32956 10276 33012 10286
rect 30828 9202 30884 9212
rect 31388 9202 31444 9212
rect 32284 9202 32340 9212
rect 32620 9660 32788 9716
rect 32844 9940 32900 9950
rect 30044 9156 30100 9166
rect 29932 9044 29988 9054
rect 29932 8932 29988 8988
rect 29820 8930 29988 8932
rect 29820 8878 29934 8930
rect 29986 8878 29988 8930
rect 29820 8876 29988 8878
rect 29596 8306 29652 8316
rect 29708 8820 29764 8830
rect 29036 7534 29038 7586
rect 29090 7534 29092 7586
rect 29036 7522 29092 7534
rect 29484 8034 29540 8046
rect 29484 7982 29486 8034
rect 29538 7982 29540 8034
rect 29484 7588 29540 7982
rect 29596 7700 29652 7710
rect 29708 7700 29764 8764
rect 29596 7698 29764 7700
rect 29596 7646 29598 7698
rect 29650 7646 29764 7698
rect 29596 7644 29764 7646
rect 29596 7634 29652 7644
rect 29484 7522 29540 7532
rect 29820 7588 29876 8876
rect 29932 8866 29988 8876
rect 30044 8372 30100 9100
rect 30604 9156 30660 9166
rect 30604 9062 30660 9100
rect 30492 9044 30548 9054
rect 30492 8950 30548 8988
rect 31500 9044 31556 9054
rect 31500 8950 31556 8988
rect 31612 9042 31668 9054
rect 31612 8990 31614 9042
rect 31666 8990 31668 9042
rect 30192 8652 30456 8662
rect 30248 8596 30296 8652
rect 30352 8596 30400 8652
rect 30192 8586 30456 8596
rect 30156 8372 30212 8382
rect 30044 8370 30212 8372
rect 30044 8318 30158 8370
rect 30210 8318 30212 8370
rect 30044 8316 30212 8318
rect 29932 7700 29988 7710
rect 30044 7700 30100 8316
rect 30156 8306 30212 8316
rect 31388 8260 31444 8270
rect 31388 8166 31444 8204
rect 31612 8148 31668 8990
rect 31724 9042 31780 9054
rect 32060 9044 32116 9054
rect 32508 9044 32564 9054
rect 31724 8990 31726 9042
rect 31778 8990 31780 9042
rect 31724 8260 31780 8990
rect 31948 9042 32564 9044
rect 31948 8990 32062 9042
rect 32114 8990 32510 9042
rect 32562 8990 32564 9042
rect 31948 8988 32564 8990
rect 31948 8596 32004 8988
rect 32060 8978 32116 8988
rect 32508 8978 32564 8988
rect 31724 8194 31780 8204
rect 31836 8540 32004 8596
rect 31836 8258 31892 8540
rect 31836 8206 31838 8258
rect 31890 8206 31892 8258
rect 31836 8194 31892 8206
rect 31612 8082 31668 8092
rect 32284 8146 32340 8158
rect 32284 8094 32286 8146
rect 32338 8094 32340 8146
rect 29932 7698 30100 7700
rect 29932 7646 29934 7698
rect 29986 7646 30100 7698
rect 29932 7644 30100 7646
rect 30716 8034 30772 8046
rect 30716 7982 30718 8034
rect 30770 7982 30772 8034
rect 29932 7634 29988 7644
rect 29820 7522 29876 7532
rect 30716 7364 30772 7982
rect 31612 7586 31668 7598
rect 31612 7534 31614 7586
rect 31666 7534 31668 7586
rect 31164 7476 31220 7486
rect 30940 7364 30996 7374
rect 30716 7308 30940 7364
rect 30192 7084 30456 7094
rect 30248 7028 30296 7084
rect 30352 7028 30400 7084
rect 30192 7018 30456 7028
rect 28924 6738 28980 6748
rect 29484 6804 29540 6814
rect 29484 6710 29540 6748
rect 27020 4846 27022 4898
rect 27074 4846 27076 4898
rect 27020 4338 27076 4846
rect 28364 4844 28532 4900
rect 28812 6692 28868 6702
rect 28812 6466 28868 6636
rect 30044 6468 30100 6478
rect 28812 6414 28814 6466
rect 28866 6414 28868 6466
rect 28812 5906 28868 6414
rect 29932 6466 30100 6468
rect 29932 6414 30046 6466
rect 30098 6414 30100 6466
rect 29932 6412 30100 6414
rect 28812 5854 28814 5906
rect 28866 5854 28868 5906
rect 28812 5346 28868 5854
rect 28812 5294 28814 5346
rect 28866 5294 28868 5346
rect 27692 4788 27748 4798
rect 27244 4676 27300 4686
rect 27244 4562 27300 4620
rect 27244 4510 27246 4562
rect 27298 4510 27300 4562
rect 27244 4498 27300 4510
rect 27692 4450 27748 4732
rect 28140 4788 28196 4798
rect 27692 4398 27694 4450
rect 27746 4398 27748 4450
rect 27692 4386 27748 4398
rect 27804 4676 27860 4686
rect 27020 4286 27022 4338
rect 27074 4286 27076 4338
rect 27020 4116 27076 4286
rect 27356 4340 27412 4350
rect 27356 4246 27412 4284
rect 27468 4338 27524 4350
rect 27468 4286 27470 4338
rect 27522 4286 27524 4338
rect 27020 3388 27076 4060
rect 27244 3668 27300 3678
rect 27468 3668 27524 4286
rect 27804 4004 27860 4620
rect 27244 3666 27524 3668
rect 27244 3614 27246 3666
rect 27298 3614 27524 3666
rect 27244 3612 27524 3614
rect 27692 3668 27748 3678
rect 27804 3668 27860 3948
rect 27692 3666 27860 3668
rect 27692 3614 27694 3666
rect 27746 3614 27860 3666
rect 27692 3612 27860 3614
rect 28140 3666 28196 4732
rect 28140 3614 28142 3666
rect 28194 3614 28196 3666
rect 27020 3332 27188 3388
rect 27132 2996 27188 3332
rect 27132 2930 27188 2940
rect 27244 1540 27300 3612
rect 27692 3602 27748 3612
rect 28140 3602 28196 3614
rect 27244 1474 27300 1484
rect 28252 3556 28308 3566
rect 26908 1250 26964 1260
rect 28252 800 28308 3500
rect 28364 3332 28420 4844
rect 28364 3266 28420 3276
rect 28476 4114 28532 4126
rect 28476 4062 28478 4114
rect 28530 4062 28532 4114
rect 28476 3220 28532 4062
rect 28588 3444 28644 3482
rect 28588 3378 28644 3388
rect 28476 3154 28532 3164
rect 28812 1316 28868 5294
rect 29708 5908 29764 5918
rect 29708 5460 29764 5852
rect 28924 5122 28980 5134
rect 28924 5070 28926 5122
rect 28978 5070 28980 5122
rect 28924 5012 28980 5070
rect 28924 4946 28980 4956
rect 29148 5124 29204 5134
rect 29148 4338 29204 5068
rect 29148 4286 29150 4338
rect 29202 4286 29204 4338
rect 29148 4274 29204 4286
rect 29708 5122 29764 5404
rect 29708 5070 29710 5122
rect 29762 5070 29764 5122
rect 29260 3556 29316 3566
rect 29260 3462 29316 3500
rect 29596 3332 29652 3342
rect 29596 3238 29652 3276
rect 29708 2324 29764 5070
rect 29820 5236 29876 5246
rect 29820 5010 29876 5180
rect 29820 4958 29822 5010
rect 29874 4958 29876 5010
rect 29820 2548 29876 4958
rect 29932 4452 29988 6412
rect 30044 6402 30100 6412
rect 30604 6466 30660 6478
rect 30604 6414 30606 6466
rect 30658 6414 30660 6466
rect 30604 6356 30660 6414
rect 30044 5908 30100 5918
rect 30044 5814 30100 5852
rect 30380 5796 30436 5806
rect 30380 5702 30436 5740
rect 30192 5516 30456 5526
rect 30248 5460 30296 5516
rect 30352 5460 30400 5516
rect 30192 5450 30456 5460
rect 29932 4386 29988 4396
rect 30044 5236 30100 5246
rect 30044 5122 30100 5180
rect 30044 5070 30046 5122
rect 30098 5070 30100 5122
rect 30044 3780 30100 5070
rect 30492 5124 30548 5134
rect 30492 5030 30548 5068
rect 30156 4452 30212 4462
rect 30156 4338 30212 4396
rect 30156 4286 30158 4338
rect 30210 4286 30212 4338
rect 30156 4274 30212 4286
rect 30604 4226 30660 6300
rect 30828 5684 30884 7308
rect 30940 7270 30996 7308
rect 31164 6690 31220 7420
rect 31500 7474 31556 7486
rect 31500 7422 31502 7474
rect 31554 7422 31556 7474
rect 31500 6804 31556 7422
rect 31500 6738 31556 6748
rect 31164 6638 31166 6690
rect 31218 6638 31220 6690
rect 31164 6626 31220 6638
rect 31612 6692 31668 7534
rect 31836 7476 31892 7486
rect 32172 7476 32228 7486
rect 31836 7474 32228 7476
rect 31836 7422 31838 7474
rect 31890 7422 32174 7474
rect 32226 7422 32228 7474
rect 31836 7420 32228 7422
rect 31836 7410 31892 7420
rect 32172 7410 32228 7420
rect 32060 6804 32116 6814
rect 32284 6804 32340 8094
rect 32620 7700 32676 9660
rect 32732 9268 32788 9278
rect 32732 9174 32788 9212
rect 32844 9154 32900 9884
rect 32844 9102 32846 9154
rect 32898 9102 32900 9154
rect 32844 8596 32900 9102
rect 32844 8530 32900 8540
rect 32732 7700 32788 7710
rect 32620 7698 32788 7700
rect 32620 7646 32734 7698
rect 32786 7646 32788 7698
rect 32620 7644 32788 7646
rect 32732 7634 32788 7644
rect 32620 7476 32676 7486
rect 32620 7382 32676 7420
rect 32844 7474 32900 7486
rect 32844 7422 32846 7474
rect 32898 7422 32900 7474
rect 32116 6748 32340 6804
rect 32508 6916 32564 6926
rect 32844 6916 32900 7422
rect 32508 6914 32900 6916
rect 32508 6862 32510 6914
rect 32562 6862 32900 6914
rect 32508 6860 32900 6862
rect 32060 6710 32116 6748
rect 31612 6626 31668 6636
rect 32396 6692 32452 6702
rect 32396 6598 32452 6636
rect 31052 6580 31108 6590
rect 31052 6486 31108 6524
rect 32060 6580 32116 6590
rect 30940 5908 30996 5918
rect 30940 5814 30996 5852
rect 32060 5906 32116 6524
rect 32060 5854 32062 5906
rect 32114 5854 32116 5906
rect 32060 5842 32116 5854
rect 32508 5906 32564 6860
rect 32508 5854 32510 5906
rect 32562 5854 32564 5906
rect 32508 5842 32564 5854
rect 32732 5908 32788 5918
rect 32732 5814 32788 5852
rect 30828 5628 30996 5684
rect 30828 5012 30884 5022
rect 30828 4918 30884 4956
rect 30716 4898 30772 4910
rect 30716 4846 30718 4898
rect 30770 4846 30772 4898
rect 30716 4788 30772 4846
rect 30716 4722 30772 4732
rect 30604 4174 30606 4226
rect 30658 4174 30660 4226
rect 30604 4162 30660 4174
rect 30192 3948 30456 3958
rect 30248 3892 30296 3948
rect 30352 3892 30400 3948
rect 30192 3882 30456 3892
rect 30044 3714 30100 3724
rect 29820 2482 29876 2492
rect 30156 3668 30212 3678
rect 30156 2436 30212 3612
rect 30156 2370 30212 2380
rect 30604 3444 30660 3482
rect 29708 2258 29764 2268
rect 30604 2212 30660 3388
rect 30940 3442 30996 5628
rect 32284 5236 32340 5246
rect 32284 5142 32340 5180
rect 32956 5010 33012 10220
rect 33180 9714 33236 10444
rect 33180 9662 33182 9714
rect 33234 9662 33236 9714
rect 33068 8596 33124 8606
rect 33068 8260 33124 8540
rect 33180 8484 33236 9662
rect 33292 9604 33348 10668
rect 33404 10388 33460 12012
rect 33740 11396 33796 11406
rect 33404 10322 33460 10332
rect 33516 11394 33796 11396
rect 33516 11342 33742 11394
rect 33794 11342 33796 11394
rect 33516 11340 33796 11342
rect 33516 9826 33572 11340
rect 33740 11330 33796 11340
rect 33852 10836 33908 15036
rect 34412 14756 34468 15262
rect 34748 15314 34804 15822
rect 34860 15876 34916 18172
rect 35308 18116 35364 18126
rect 35196 17780 35252 17790
rect 35196 17554 35252 17724
rect 35308 17666 35364 18060
rect 35308 17614 35310 17666
rect 35362 17614 35364 17666
rect 35308 17602 35364 17614
rect 35196 17502 35198 17554
rect 35250 17502 35252 17554
rect 35196 17490 35252 17502
rect 34972 17442 35028 17454
rect 34972 17390 34974 17442
rect 35026 17390 35028 17442
rect 34972 17108 35028 17390
rect 34972 17042 35028 17052
rect 35196 17220 35252 17230
rect 34972 16882 35028 16894
rect 34972 16830 34974 16882
rect 35026 16830 35028 16882
rect 34972 16324 35028 16830
rect 34972 16258 35028 16268
rect 35084 16770 35140 16782
rect 35084 16718 35086 16770
rect 35138 16718 35140 16770
rect 35084 16098 35140 16718
rect 35084 16046 35086 16098
rect 35138 16046 35140 16098
rect 35084 16034 35140 16046
rect 35196 15876 35252 17164
rect 35420 16212 35476 16222
rect 35420 16098 35476 16156
rect 35420 16046 35422 16098
rect 35474 16046 35476 16098
rect 35420 16034 35476 16046
rect 35308 15876 35364 15886
rect 35532 15876 35588 19628
rect 35868 19236 35924 20524
rect 35980 20130 36036 20860
rect 36092 20850 36148 20860
rect 36204 20916 36260 21980
rect 36204 20850 36260 20860
rect 36316 22146 36484 22148
rect 36316 22094 36430 22146
rect 36482 22094 36484 22146
rect 36316 22092 36484 22094
rect 36316 21476 36372 22092
rect 36428 22082 36484 22092
rect 36540 21812 36596 22204
rect 36764 22148 36820 22158
rect 36764 22054 36820 22092
rect 35980 20078 35982 20130
rect 36034 20078 36036 20130
rect 35980 20066 36036 20078
rect 36092 20692 36148 20702
rect 36092 19684 36148 20636
rect 36316 20188 36372 21420
rect 36092 19618 36148 19628
rect 36204 20132 36372 20188
rect 36428 21756 36596 21812
rect 36652 22036 36708 22046
rect 36652 21810 36708 21980
rect 36652 21758 36654 21810
rect 36706 21758 36708 21810
rect 36092 19348 36148 19358
rect 35644 19234 35924 19236
rect 35644 19182 35870 19234
rect 35922 19182 35924 19234
rect 35644 19180 35924 19182
rect 35644 18674 35700 19180
rect 35868 19170 35924 19180
rect 35980 19346 36148 19348
rect 35980 19294 36094 19346
rect 36146 19294 36148 19346
rect 35980 19292 36148 19294
rect 35980 19124 36036 19292
rect 36092 19282 36148 19292
rect 35644 18622 35646 18674
rect 35698 18622 35700 18674
rect 35644 18610 35700 18622
rect 35868 18676 35924 18686
rect 35980 18676 36036 19068
rect 35868 18674 36036 18676
rect 35868 18622 35870 18674
rect 35922 18622 36036 18674
rect 35868 18620 36036 18622
rect 35868 18610 35924 18620
rect 35756 18338 35812 18350
rect 35756 18286 35758 18338
rect 35810 18286 35812 18338
rect 34860 15820 35140 15876
rect 34748 15262 34750 15314
rect 34802 15262 34804 15314
rect 34748 15250 34804 15262
rect 34412 14690 34468 14700
rect 34860 14868 34916 14878
rect 33964 14532 34020 14542
rect 34748 14532 34804 14542
rect 33964 14418 34020 14476
rect 33964 14366 33966 14418
rect 34018 14366 34020 14418
rect 33964 12962 34020 14366
rect 34636 14530 34804 14532
rect 34636 14478 34750 14530
rect 34802 14478 34804 14530
rect 34636 14476 34804 14478
rect 33964 12910 33966 12962
rect 34018 12910 34020 12962
rect 33964 12898 34020 12910
rect 34076 13636 34132 13646
rect 34076 12740 34132 13580
rect 34636 13636 34692 14476
rect 34748 14466 34804 14476
rect 34748 14308 34804 14318
rect 34748 13746 34804 14252
rect 34748 13694 34750 13746
rect 34802 13694 34804 13746
rect 34748 13682 34804 13694
rect 34860 13748 34916 14812
rect 34972 14532 35028 14542
rect 34972 14438 35028 14476
rect 35084 13970 35140 15820
rect 35196 15874 35364 15876
rect 35196 15822 35310 15874
rect 35362 15822 35364 15874
rect 35196 15820 35364 15822
rect 35196 15538 35252 15820
rect 35308 15810 35364 15820
rect 35420 15820 35588 15876
rect 35644 18228 35700 18238
rect 35196 15486 35198 15538
rect 35250 15486 35252 15538
rect 35196 15474 35252 15486
rect 35308 14308 35364 14318
rect 35308 14214 35364 14252
rect 35084 13918 35086 13970
rect 35138 13918 35140 13970
rect 35084 13906 35140 13918
rect 34860 13654 34916 13692
rect 35308 13748 35364 13758
rect 35308 13654 35364 13692
rect 34636 13570 34692 13580
rect 34076 12674 34132 12684
rect 34188 12850 34244 12862
rect 34188 12798 34190 12850
rect 34242 12798 34244 12850
rect 34188 12178 34244 12798
rect 34748 12292 34804 12302
rect 34748 12198 34804 12236
rect 34188 12126 34190 12178
rect 34242 12126 34244 12178
rect 34188 11394 34244 12126
rect 34412 12066 34468 12078
rect 34412 12014 34414 12066
rect 34466 12014 34468 12066
rect 34300 11508 34356 11518
rect 34300 11414 34356 11452
rect 34188 11342 34190 11394
rect 34242 11342 34244 11394
rect 34188 11330 34244 11342
rect 34412 11394 34468 12014
rect 35420 11732 35476 15820
rect 35644 15538 35700 18172
rect 35644 15486 35646 15538
rect 35698 15486 35700 15538
rect 35644 14756 35700 15486
rect 35756 14868 35812 18286
rect 36204 18004 36260 20132
rect 36428 19348 36484 21756
rect 36652 21746 36708 21758
rect 36540 21588 36596 21598
rect 36540 21026 36596 21532
rect 36540 20974 36542 21026
rect 36594 20974 36596 21026
rect 36540 20962 36596 20974
rect 36652 21586 36708 21598
rect 36652 21534 36654 21586
rect 36706 21534 36708 21586
rect 36652 21028 36708 21534
rect 36652 20962 36708 20972
rect 36764 19348 36820 19358
rect 36428 19346 36820 19348
rect 36428 19294 36766 19346
rect 36818 19294 36820 19346
rect 36428 19292 36820 19294
rect 35868 17948 36260 18004
rect 36428 18900 36484 18910
rect 35868 17108 35924 17948
rect 36428 17668 36484 18844
rect 36540 18562 36596 19292
rect 36764 19282 36820 19292
rect 36652 18676 36708 18686
rect 36652 18582 36708 18620
rect 36540 18510 36542 18562
rect 36594 18510 36596 18562
rect 36540 18498 36596 18510
rect 36652 18226 36708 18238
rect 36652 18174 36654 18226
rect 36706 18174 36708 18226
rect 36316 17666 36484 17668
rect 36316 17614 36430 17666
rect 36482 17614 36484 17666
rect 36316 17612 36484 17614
rect 35980 17556 36036 17566
rect 36316 17556 36372 17612
rect 36428 17602 36484 17612
rect 36540 17780 36596 17790
rect 35980 17554 36372 17556
rect 35980 17502 35982 17554
rect 36034 17502 36372 17554
rect 35980 17500 36372 17502
rect 36540 17554 36596 17724
rect 36540 17502 36542 17554
rect 36594 17502 36596 17554
rect 35980 17490 36036 17500
rect 36540 17490 36596 17502
rect 36652 17220 36708 18174
rect 36764 17668 36820 17678
rect 36764 17574 36820 17612
rect 36540 17164 36708 17220
rect 35868 17052 36148 17108
rect 35868 16884 35924 16894
rect 35868 16790 35924 16828
rect 35868 16212 35924 16222
rect 35868 16118 35924 16156
rect 35756 14802 35812 14812
rect 35644 14690 35700 14700
rect 35980 14532 36036 14542
rect 35756 14306 35812 14318
rect 35756 14254 35758 14306
rect 35810 14254 35812 14306
rect 35756 13636 35812 14254
rect 35980 13746 36036 14476
rect 35980 13694 35982 13746
rect 36034 13694 36036 13746
rect 35980 13682 36036 13694
rect 35756 13542 35812 13580
rect 35644 13300 35700 13310
rect 35532 12740 35588 12750
rect 35532 11956 35588 12684
rect 35532 11890 35588 11900
rect 35420 11666 35476 11676
rect 34412 11342 34414 11394
rect 34466 11342 34468 11394
rect 33852 10780 34132 10836
rect 33516 9774 33518 9826
rect 33570 9774 33572 9826
rect 33516 9762 33572 9774
rect 33852 10610 33908 10622
rect 33852 10558 33854 10610
rect 33906 10558 33908 10610
rect 33852 9604 33908 10558
rect 33964 10500 34020 10510
rect 33964 10406 34020 10444
rect 33292 9602 33908 9604
rect 33292 9550 33294 9602
rect 33346 9550 33854 9602
rect 33906 9550 33908 9602
rect 33292 9548 33908 9550
rect 33292 9538 33348 9548
rect 33180 8428 33348 8484
rect 33180 8260 33236 8270
rect 33068 8258 33236 8260
rect 33068 8206 33182 8258
rect 33234 8206 33236 8258
rect 33068 8204 33236 8206
rect 33180 8194 33236 8204
rect 32956 4958 32958 5010
rect 33010 4958 33012 5010
rect 32956 4946 33012 4958
rect 31164 4900 31220 4910
rect 31164 4564 31220 4844
rect 31276 4900 31332 4910
rect 31948 4900 32004 4910
rect 31276 4898 31444 4900
rect 31276 4846 31278 4898
rect 31330 4846 31444 4898
rect 31276 4844 31444 4846
rect 31276 4834 31332 4844
rect 31388 4788 31444 4844
rect 31948 4806 32004 4844
rect 32172 4900 32228 4910
rect 32844 4900 32900 4910
rect 31276 4564 31332 4574
rect 31164 4508 31276 4564
rect 31276 4432 31332 4508
rect 31388 4228 31444 4732
rect 31388 4162 31444 4172
rect 31948 4564 32004 4574
rect 31948 3666 32004 4508
rect 31948 3614 31950 3666
rect 32002 3614 32004 3666
rect 31948 3602 32004 3614
rect 32172 4338 32228 4844
rect 32172 4286 32174 4338
rect 32226 4286 32228 4338
rect 32172 3668 32228 4286
rect 32732 4898 32900 4900
rect 32732 4846 32846 4898
rect 32898 4846 32900 4898
rect 32732 4844 32900 4846
rect 32732 4340 32788 4844
rect 32844 4834 32900 4844
rect 33068 4900 33124 4910
rect 33068 4806 33124 4844
rect 32844 4452 32900 4462
rect 33292 4452 33348 8428
rect 33404 7924 33460 9548
rect 33852 9538 33908 9548
rect 34076 9380 34132 10780
rect 33852 9324 34132 9380
rect 33852 9266 33908 9324
rect 33852 9214 33854 9266
rect 33906 9214 33908 9266
rect 33852 9202 33908 9214
rect 34076 9268 34132 9324
rect 34076 9202 34132 9212
rect 34188 10500 34244 10510
rect 34188 9044 34244 10444
rect 34412 10386 34468 11342
rect 35532 11620 35588 11630
rect 35532 11394 35588 11564
rect 35532 11342 35534 11394
rect 35586 11342 35588 11394
rect 35532 11330 35588 11342
rect 34972 11172 35028 11182
rect 34972 10724 35028 11116
rect 35644 11172 35700 13244
rect 35980 12852 36036 12862
rect 35980 12738 36036 12796
rect 35980 12686 35982 12738
rect 36034 12686 36036 12738
rect 35980 12068 36036 12686
rect 35980 11974 36036 12012
rect 35644 11078 35700 11116
rect 35868 11170 35924 11182
rect 35868 11118 35870 11170
rect 35922 11118 35924 11170
rect 34972 10658 35028 10668
rect 34412 10334 34414 10386
rect 34466 10334 34468 10386
rect 34412 10322 34468 10334
rect 35420 10612 35476 10622
rect 35420 10052 35476 10556
rect 35868 10610 35924 11118
rect 36092 11060 36148 17052
rect 36540 16882 36596 17164
rect 36876 17108 36932 23660
rect 37772 23716 37828 23726
rect 37884 23716 37940 23996
rect 37996 23938 38052 24556
rect 38108 24052 38164 24062
rect 38108 23958 38164 23996
rect 37996 23886 37998 23938
rect 38050 23886 38052 23938
rect 37996 23874 38052 23886
rect 38220 23716 38276 25228
rect 38892 24722 38948 24734
rect 38892 24670 38894 24722
rect 38946 24670 38948 24722
rect 38780 24610 38836 24622
rect 38780 24558 38782 24610
rect 38834 24558 38836 24610
rect 38780 23938 38836 24558
rect 38780 23886 38782 23938
rect 38834 23886 38836 23938
rect 38780 23828 38836 23886
rect 37884 23714 38276 23716
rect 37884 23662 38222 23714
rect 38274 23662 38276 23714
rect 37884 23660 38276 23662
rect 37772 23622 37828 23660
rect 37212 23268 37268 23278
rect 37212 23042 37268 23212
rect 37212 22990 37214 23042
rect 37266 22990 37268 23042
rect 36988 22148 37044 22158
rect 36988 17220 37044 22092
rect 37212 20188 37268 22990
rect 38108 23044 38164 23054
rect 38220 23044 38276 23660
rect 38108 23042 38276 23044
rect 38108 22990 38110 23042
rect 38162 22990 38276 23042
rect 38108 22988 38276 22990
rect 38108 22978 38164 22988
rect 37660 22370 37716 22382
rect 37884 22372 37940 22382
rect 37660 22318 37662 22370
rect 37714 22318 37716 22370
rect 37660 22148 37716 22318
rect 37660 22082 37716 22092
rect 37772 22370 37940 22372
rect 37772 22318 37886 22370
rect 37938 22318 37940 22370
rect 37772 22316 37940 22318
rect 37324 21586 37380 21598
rect 37324 21534 37326 21586
rect 37378 21534 37380 21586
rect 37324 21476 37380 21534
rect 37772 21588 37828 22316
rect 37884 22306 37940 22316
rect 37996 22148 38052 22158
rect 37996 21810 38052 22092
rect 37996 21758 37998 21810
rect 38050 21758 38052 21810
rect 37996 21746 38052 21758
rect 37884 21700 37940 21710
rect 37884 21606 37940 21644
rect 37772 21494 37828 21532
rect 37324 21410 37380 21420
rect 38108 20916 38164 20926
rect 38108 20822 38164 20860
rect 37772 20578 37828 20590
rect 37772 20526 37774 20578
rect 37826 20526 37828 20578
rect 37772 20468 37828 20526
rect 37772 20402 37828 20412
rect 38220 20188 38276 22988
rect 38556 23772 38836 23828
rect 38892 24052 38948 24670
rect 38892 23826 38948 23996
rect 39116 23940 39172 23950
rect 39228 23940 39284 25228
rect 39116 23938 39284 23940
rect 39116 23886 39118 23938
rect 39170 23886 39284 23938
rect 39116 23884 39284 23886
rect 39116 23874 39172 23884
rect 38892 23774 38894 23826
rect 38946 23774 38948 23826
rect 38556 22482 38612 23772
rect 38892 23762 38948 23774
rect 38668 23156 38724 23166
rect 38668 23062 38724 23100
rect 38556 22430 38558 22482
rect 38610 22430 38612 22482
rect 38556 22418 38612 22430
rect 38444 22148 38500 22158
rect 38444 21810 38500 22092
rect 38444 21758 38446 21810
rect 38498 21758 38500 21810
rect 38444 21746 38500 21758
rect 39340 21700 39396 25452
rect 39452 24834 39508 26124
rect 39564 25844 39620 26572
rect 39564 25778 39620 25788
rect 39676 25506 39732 26796
rect 39900 26852 39956 26910
rect 39900 26786 39956 26796
rect 39852 26684 40116 26694
rect 39908 26628 39956 26684
rect 40012 26628 40060 26684
rect 39852 26618 40116 26628
rect 39900 26404 39956 26414
rect 39788 26292 39844 26302
rect 39788 25618 39844 26236
rect 39900 26290 39956 26348
rect 39900 26238 39902 26290
rect 39954 26238 39956 26290
rect 39900 26226 39956 26238
rect 40236 26178 40292 28476
rect 40796 27970 40852 29372
rect 40908 28866 40964 29932
rect 41356 29988 41412 29998
rect 41356 29894 41412 29932
rect 41804 29428 41860 29438
rect 41804 29334 41860 29372
rect 40908 28814 40910 28866
rect 40962 28814 40964 28866
rect 40908 28756 40964 28814
rect 40908 28690 40964 28700
rect 41132 29316 41188 29326
rect 41132 28754 41188 29260
rect 41692 29316 41748 29326
rect 41692 29222 41748 29260
rect 41132 28702 41134 28754
rect 41186 28702 41188 28754
rect 41132 28690 41188 28702
rect 42140 28082 42196 30716
rect 43148 29988 43204 29998
rect 43148 29426 43204 29932
rect 43708 29538 43764 30940
rect 43820 30930 43876 30940
rect 45388 30882 45444 31724
rect 45388 30830 45390 30882
rect 45442 30830 45444 30882
rect 45388 30772 45444 30830
rect 45388 30706 45444 30716
rect 44716 30322 44772 30334
rect 44716 30270 44718 30322
rect 44770 30270 44772 30322
rect 44716 30212 44772 30270
rect 44716 30146 44772 30156
rect 44380 30098 44436 30110
rect 44380 30046 44382 30098
rect 44434 30046 44436 30098
rect 43820 29988 43876 29998
rect 44380 29988 44436 30046
rect 43820 29986 44436 29988
rect 43820 29934 43822 29986
rect 43874 29934 44436 29986
rect 43820 29932 44436 29934
rect 43820 29922 43876 29932
rect 43708 29486 43710 29538
rect 43762 29486 43764 29538
rect 43708 29474 43764 29486
rect 43148 29374 43150 29426
rect 43202 29374 43204 29426
rect 43148 29362 43204 29374
rect 44380 29314 44436 29932
rect 44604 29986 44660 29998
rect 44604 29934 44606 29986
rect 44658 29934 44660 29986
rect 44380 29262 44382 29314
rect 44434 29262 44436 29314
rect 44380 28532 44436 29262
rect 44380 28466 44436 28476
rect 44492 29876 44548 29886
rect 42140 28030 42142 28082
rect 42194 28030 42196 28082
rect 42140 28018 42196 28030
rect 40796 27918 40798 27970
rect 40850 27918 40852 27970
rect 40796 27906 40852 27918
rect 41580 27748 41636 27758
rect 41580 27654 41636 27692
rect 41804 27636 41860 27646
rect 41804 27542 41860 27580
rect 41692 27524 41748 27534
rect 40796 27188 40852 27198
rect 40572 27074 40628 27086
rect 40572 27022 40574 27074
rect 40626 27022 40628 27074
rect 40572 26908 40628 27022
rect 40236 26126 40238 26178
rect 40290 26126 40292 26178
rect 40236 26114 40292 26126
rect 40348 26852 40628 26908
rect 39788 25566 39790 25618
rect 39842 25566 39844 25618
rect 39788 25554 39844 25566
rect 40348 25844 40404 26852
rect 39676 25454 39678 25506
rect 39730 25454 39732 25506
rect 39676 25396 39732 25454
rect 39900 25508 39956 25518
rect 39900 25414 39956 25452
rect 40124 25508 40180 25518
rect 40124 25414 40180 25452
rect 39676 25330 39732 25340
rect 40348 25394 40404 25788
rect 40796 25618 40852 27132
rect 41244 27188 41300 27198
rect 41244 27074 41300 27132
rect 41244 27022 41246 27074
rect 41298 27022 41300 27074
rect 41244 27010 41300 27022
rect 41692 26852 41748 27468
rect 42252 27412 42308 27422
rect 42140 27188 42196 27198
rect 42140 27094 42196 27132
rect 41692 26758 41748 26796
rect 41916 26404 41972 26414
rect 41916 26310 41972 26348
rect 40796 25566 40798 25618
rect 40850 25566 40852 25618
rect 40796 25508 40852 25566
rect 40796 25442 40852 25452
rect 41468 26290 41524 26302
rect 41468 26238 41470 26290
rect 41522 26238 41524 26290
rect 40348 25342 40350 25394
rect 40402 25342 40404 25394
rect 39852 25116 40116 25126
rect 39908 25060 39956 25116
rect 40012 25060 40060 25116
rect 39852 25050 40116 25060
rect 39452 24782 39454 24834
rect 39506 24782 39508 24834
rect 39452 24770 39508 24782
rect 39564 24052 39620 24062
rect 40348 24052 40404 25342
rect 41244 25396 41300 25406
rect 41244 25302 41300 25340
rect 41468 25284 41524 26238
rect 42028 26292 42084 26302
rect 42028 26198 42084 26236
rect 42140 26290 42196 26302
rect 42140 26238 42142 26290
rect 42194 26238 42196 26290
rect 42140 26180 42196 26238
rect 42140 26114 42196 26124
rect 41468 25218 41524 25228
rect 42028 25284 42084 25294
rect 40460 24164 40516 24174
rect 41020 24164 41076 24174
rect 40460 24162 41972 24164
rect 40460 24110 40462 24162
rect 40514 24110 41022 24162
rect 41074 24110 41972 24162
rect 40460 24108 41972 24110
rect 40460 24098 40516 24108
rect 41020 24098 41076 24108
rect 39564 24050 40404 24052
rect 39564 23998 39566 24050
rect 39618 23998 40404 24050
rect 39564 23996 40404 23998
rect 39564 23986 39620 23996
rect 40348 23940 40404 23996
rect 40348 23884 40516 23940
rect 40124 23828 40180 23838
rect 40124 23826 40292 23828
rect 40124 23774 40126 23826
rect 40178 23774 40292 23826
rect 40124 23772 40292 23774
rect 40124 23762 40180 23772
rect 39852 23548 40116 23558
rect 39908 23492 39956 23548
rect 40012 23492 40060 23548
rect 39852 23482 40116 23492
rect 40236 23380 40292 23772
rect 40124 23324 40292 23380
rect 40348 23714 40404 23726
rect 40348 23662 40350 23714
rect 40402 23662 40404 23714
rect 39564 23156 39620 23166
rect 39564 23062 39620 23100
rect 39452 23042 39508 23054
rect 39452 22990 39454 23042
rect 39506 22990 39508 23042
rect 39452 22932 39508 22990
rect 40124 22932 40180 23324
rect 40236 23156 40292 23166
rect 40348 23156 40404 23662
rect 40460 23378 40516 23884
rect 41916 23938 41972 24108
rect 42028 24050 42084 25228
rect 42028 23998 42030 24050
rect 42082 23998 42084 24050
rect 42028 23986 42084 23998
rect 41916 23886 41918 23938
rect 41970 23886 41972 23938
rect 41916 23874 41972 23886
rect 41132 23828 41188 23838
rect 41132 23734 41188 23772
rect 41244 23716 41300 23726
rect 41692 23716 41748 23726
rect 41244 23714 41692 23716
rect 41244 23662 41246 23714
rect 41298 23662 41692 23714
rect 41244 23660 41692 23662
rect 41244 23650 41300 23660
rect 40460 23326 40462 23378
rect 40514 23326 40516 23378
rect 40460 23314 40516 23326
rect 41692 23378 41748 23660
rect 42140 23716 42196 23726
rect 42140 23622 42196 23660
rect 41692 23326 41694 23378
rect 41746 23326 41748 23378
rect 41692 23314 41748 23326
rect 42252 23380 42308 27356
rect 44492 27188 44548 29820
rect 44604 29652 44660 29934
rect 44604 29586 44660 29596
rect 45276 29652 45332 29662
rect 45276 29426 45332 29596
rect 45500 29540 45556 32620
rect 46060 31780 46116 33180
rect 47404 33180 47684 33236
rect 46620 32674 46676 32686
rect 46620 32622 46622 32674
rect 46674 32622 46676 32674
rect 46508 32564 46564 32574
rect 46172 32452 46228 32462
rect 46172 32450 46452 32452
rect 46172 32398 46174 32450
rect 46226 32398 46452 32450
rect 46172 32396 46452 32398
rect 46172 32386 46228 32396
rect 46172 31780 46228 31790
rect 46060 31778 46228 31780
rect 46060 31726 46174 31778
rect 46226 31726 46228 31778
rect 46060 31724 46228 31726
rect 46172 31714 46228 31724
rect 46396 31778 46452 32396
rect 46508 31890 46564 32508
rect 46508 31838 46510 31890
rect 46562 31838 46564 31890
rect 46508 31826 46564 31838
rect 46396 31726 46398 31778
rect 46450 31726 46452 31778
rect 46396 31220 46452 31726
rect 46620 31780 46676 32622
rect 46620 31714 46676 31724
rect 46956 31780 47012 31790
rect 46844 31668 46900 31678
rect 46844 31574 46900 31612
rect 46620 31554 46676 31566
rect 46620 31502 46622 31554
rect 46674 31502 46676 31554
rect 46396 31154 46452 31164
rect 46508 31220 46564 31230
rect 46620 31220 46676 31502
rect 46508 31218 46676 31220
rect 46508 31166 46510 31218
rect 46562 31166 46676 31218
rect 46508 31164 46676 31166
rect 46508 31154 46564 31164
rect 45948 30882 46004 30894
rect 45948 30830 45950 30882
rect 46002 30830 46004 30882
rect 45948 30772 46004 30830
rect 45948 30706 46004 30716
rect 46172 30884 46228 30894
rect 46172 30436 46228 30828
rect 45500 29474 45556 29484
rect 45948 30380 46228 30436
rect 46956 30884 47012 31724
rect 47292 31668 47348 31678
rect 47292 31574 47348 31612
rect 45948 29538 46004 30380
rect 46060 30212 46116 30222
rect 46060 30118 46116 30156
rect 46956 30210 47012 30828
rect 46956 30158 46958 30210
rect 47010 30158 47012 30210
rect 46956 30146 47012 30158
rect 47180 30100 47236 30110
rect 47180 30006 47236 30044
rect 45948 29486 45950 29538
rect 46002 29486 46004 29538
rect 45948 29474 46004 29486
rect 46284 29986 46340 29998
rect 46284 29934 46286 29986
rect 46338 29934 46340 29986
rect 45276 29374 45278 29426
rect 45330 29374 45332 29426
rect 45276 29362 45332 29374
rect 45052 29314 45108 29326
rect 45052 29262 45054 29314
rect 45106 29262 45108 29314
rect 45052 28532 45108 29262
rect 45052 28466 45108 28476
rect 45388 28756 45444 28766
rect 46284 28756 46340 29934
rect 46508 29540 46564 29550
rect 46508 29446 46564 29484
rect 46844 29428 46900 29438
rect 46844 29334 46900 29372
rect 46396 28756 46452 28766
rect 46284 28754 46452 28756
rect 46284 28702 46398 28754
rect 46450 28702 46452 28754
rect 46284 28700 46452 28702
rect 45052 27972 45108 27982
rect 45052 27858 45108 27916
rect 45052 27806 45054 27858
rect 45106 27806 45108 27858
rect 45052 27794 45108 27806
rect 45276 27860 45332 27870
rect 45276 27766 45332 27804
rect 45388 27746 45444 28700
rect 46396 28644 46452 28700
rect 46396 28578 46452 28588
rect 46620 28756 46676 28766
rect 46620 28642 46676 28700
rect 46620 28590 46622 28642
rect 46674 28590 46676 28642
rect 46620 28578 46676 28590
rect 47292 28530 47348 28542
rect 47292 28478 47294 28530
rect 47346 28478 47348 28530
rect 47292 28196 47348 28478
rect 47292 28130 47348 28140
rect 45724 27972 45780 27982
rect 45388 27694 45390 27746
rect 45442 27694 45444 27746
rect 45388 27682 45444 27694
rect 45500 27860 45556 27870
rect 44492 27122 44548 27132
rect 44716 27188 44772 27198
rect 44716 27094 44772 27132
rect 45500 27188 45556 27804
rect 44044 27074 44100 27086
rect 44044 27022 44046 27074
rect 44098 27022 44100 27074
rect 43260 26740 43316 26750
rect 43148 26516 43204 26526
rect 43148 26422 43204 26460
rect 42588 24722 42644 24734
rect 42588 24670 42590 24722
rect 42642 24670 42644 24722
rect 42364 24276 42420 24286
rect 42588 24276 42644 24670
rect 42420 24220 42644 24276
rect 42700 24610 42756 24622
rect 42700 24558 42702 24610
rect 42754 24558 42756 24610
rect 42364 23826 42420 24220
rect 42364 23774 42366 23826
rect 42418 23774 42420 23826
rect 42364 23762 42420 23774
rect 42700 23828 42756 24558
rect 42700 23762 42756 23772
rect 42252 23314 42308 23324
rect 40292 23100 40404 23156
rect 40572 23154 40628 23166
rect 40572 23102 40574 23154
rect 40626 23102 40628 23154
rect 40236 23062 40292 23100
rect 39452 22876 40180 22932
rect 40124 22594 40180 22876
rect 40572 22708 40628 23102
rect 40908 23156 40964 23166
rect 40572 22642 40628 22652
rect 40796 22930 40852 22942
rect 40796 22878 40798 22930
rect 40850 22878 40852 22930
rect 40124 22542 40126 22594
rect 40178 22542 40180 22594
rect 40124 22530 40180 22542
rect 40796 22484 40852 22878
rect 40572 22482 40852 22484
rect 40572 22430 40798 22482
rect 40850 22430 40852 22482
rect 40572 22428 40852 22430
rect 40348 22372 40404 22382
rect 39852 21980 40116 21990
rect 39908 21924 39956 21980
rect 40012 21924 40060 21980
rect 39852 21914 40116 21924
rect 40348 21810 40404 22316
rect 40348 21758 40350 21810
rect 40402 21758 40404 21810
rect 40348 21746 40404 21758
rect 39340 21644 39732 21700
rect 39004 21476 39060 21486
rect 39452 21476 39508 21486
rect 39004 21474 39396 21476
rect 39004 21422 39006 21474
rect 39058 21422 39396 21474
rect 39004 21420 39396 21422
rect 39004 21410 39060 21420
rect 38668 20916 38724 20926
rect 38668 20802 38724 20860
rect 39228 20916 39284 20926
rect 39228 20822 39284 20860
rect 38668 20750 38670 20802
rect 38722 20750 38724 20802
rect 38668 20738 38724 20750
rect 39340 20802 39396 21420
rect 39340 20750 39342 20802
rect 39394 20750 39396 20802
rect 38892 20578 38948 20590
rect 38892 20526 38894 20578
rect 38946 20526 38948 20578
rect 37212 20132 37604 20188
rect 37100 19906 37156 19918
rect 37100 19854 37102 19906
rect 37154 19854 37156 19906
rect 37100 19684 37156 19854
rect 37100 18676 37156 19628
rect 37548 19458 37604 20132
rect 38108 20132 38164 20142
rect 38220 20132 38388 20188
rect 37548 19406 37550 19458
rect 37602 19406 37604 19458
rect 37100 18610 37156 18620
rect 37212 19124 37268 19134
rect 36988 17164 37156 17220
rect 36540 16830 36542 16882
rect 36594 16830 36596 16882
rect 36540 16818 36596 16830
rect 36652 17052 36932 17108
rect 36204 14756 36260 14766
rect 36204 14642 36260 14700
rect 36204 14590 36206 14642
rect 36258 14590 36260 14642
rect 36204 14578 36260 14590
rect 36316 13748 36372 13758
rect 36316 13634 36372 13692
rect 36316 13582 36318 13634
rect 36370 13582 36372 13634
rect 36316 13570 36372 13582
rect 36652 13186 36708 17052
rect 36988 16996 37044 17006
rect 36876 16940 36988 16996
rect 36876 16882 36932 16940
rect 36988 16930 37044 16940
rect 36876 16830 36878 16882
rect 36930 16830 36932 16882
rect 36876 16818 36932 16830
rect 36652 13134 36654 13186
rect 36706 13134 36708 13186
rect 36652 13122 36708 13134
rect 36540 12852 36596 12862
rect 36540 12758 36596 12796
rect 36652 12740 36708 12750
rect 36652 12646 36708 12684
rect 37100 12628 37156 17164
rect 37212 16212 37268 19068
rect 37548 18674 37604 19406
rect 37548 18622 37550 18674
rect 37602 18622 37604 18674
rect 37548 18610 37604 18622
rect 37660 20020 37716 20030
rect 37660 19346 37716 19964
rect 37660 19294 37662 19346
rect 37714 19294 37716 19346
rect 37660 18676 37716 19294
rect 38108 19346 38164 20076
rect 38108 19294 38110 19346
rect 38162 19294 38164 19346
rect 38108 19282 38164 19294
rect 37660 18610 37716 18620
rect 37996 18340 38052 18350
rect 37996 18246 38052 18284
rect 37772 17778 37828 17790
rect 37772 17726 37774 17778
rect 37826 17726 37828 17778
rect 37548 17668 37604 17678
rect 37548 16882 37604 17612
rect 37548 16830 37550 16882
rect 37602 16830 37604 16882
rect 37548 16818 37604 16830
rect 37772 16884 37828 17726
rect 37884 17668 37940 17678
rect 37884 17574 37940 17612
rect 37772 16790 37828 16828
rect 37884 16772 37940 16782
rect 37884 16658 37940 16716
rect 37884 16606 37886 16658
rect 37938 16606 37940 16658
rect 37884 16594 37940 16606
rect 37212 16146 37268 16156
rect 37660 16100 37716 16110
rect 37660 15876 37716 16044
rect 37548 15874 37716 15876
rect 37548 15822 37662 15874
rect 37714 15822 37716 15874
rect 37548 15820 37716 15822
rect 37548 15316 37604 15820
rect 37660 15810 37716 15820
rect 37548 15250 37604 15260
rect 38220 15202 38276 15214
rect 38220 15150 38222 15202
rect 38274 15150 38276 15202
rect 38220 14644 38276 15150
rect 37996 14642 38276 14644
rect 37996 14590 38222 14642
rect 38274 14590 38276 14642
rect 37996 14588 38276 14590
rect 37660 14308 37716 14318
rect 37548 14306 37716 14308
rect 37548 14254 37662 14306
rect 37714 14254 37716 14306
rect 37548 14252 37716 14254
rect 37324 13860 37380 13870
rect 37212 13636 37268 13646
rect 37324 13636 37380 13804
rect 37548 13860 37604 14252
rect 37660 14242 37716 14252
rect 37772 14308 37828 14318
rect 37660 13972 37716 13982
rect 37772 13972 37828 14252
rect 37660 13970 37828 13972
rect 37660 13918 37662 13970
rect 37714 13918 37828 13970
rect 37660 13916 37828 13918
rect 37660 13906 37716 13916
rect 37548 13794 37604 13804
rect 37884 13860 37940 13870
rect 37884 13766 37940 13804
rect 37996 13858 38052 14588
rect 38220 14578 38276 14588
rect 37996 13806 37998 13858
rect 38050 13806 38052 13858
rect 37996 13794 38052 13806
rect 37212 13634 37380 13636
rect 37212 13582 37214 13634
rect 37266 13582 37380 13634
rect 37212 13580 37380 13582
rect 37212 13570 37268 13580
rect 37100 12562 37156 12572
rect 37212 12740 37268 12750
rect 37212 12402 37268 12684
rect 37212 12350 37214 12402
rect 37266 12350 37268 12402
rect 37212 12338 37268 12350
rect 36204 11620 36260 11630
rect 36204 11506 36260 11564
rect 36204 11454 36206 11506
rect 36258 11454 36260 11506
rect 36204 11442 36260 11454
rect 36092 10994 36148 11004
rect 35868 10558 35870 10610
rect 35922 10558 35924 10610
rect 35756 10388 35812 10398
rect 35532 10052 35588 10062
rect 35420 10050 35588 10052
rect 35420 9998 35534 10050
rect 35586 9998 35588 10050
rect 35420 9996 35588 9998
rect 35532 9986 35588 9996
rect 35644 10052 35700 10062
rect 34748 9716 34804 9726
rect 34300 9380 34356 9390
rect 34300 9266 34356 9324
rect 34300 9214 34302 9266
rect 34354 9214 34356 9266
rect 34300 9202 34356 9214
rect 34188 8978 34244 8988
rect 34748 8372 34804 9660
rect 34972 9716 35028 9726
rect 34972 9622 35028 9660
rect 34860 9380 34916 9390
rect 34860 9156 34916 9324
rect 34972 9268 35028 9278
rect 34972 9174 35028 9212
rect 35308 9268 35364 9278
rect 34860 9024 34916 9100
rect 35196 9042 35252 9054
rect 35196 8990 35198 9042
rect 35250 8990 35252 9042
rect 34860 8372 34916 8382
rect 34748 8370 34916 8372
rect 34748 8318 34862 8370
rect 34914 8318 34916 8370
rect 34748 8316 34916 8318
rect 34860 8306 34916 8316
rect 33404 7858 33460 7868
rect 35196 7364 35252 8990
rect 35308 8370 35364 9212
rect 35644 9044 35700 9996
rect 35756 9938 35812 10332
rect 35756 9886 35758 9938
rect 35810 9886 35812 9938
rect 35756 9874 35812 9886
rect 35868 9826 35924 10558
rect 36316 10500 36372 10510
rect 36316 10406 36372 10444
rect 36876 10498 36932 10510
rect 36876 10446 36878 10498
rect 36930 10446 36932 10498
rect 36876 9940 36932 10446
rect 35868 9774 35870 9826
rect 35922 9774 35924 9826
rect 35868 9762 35924 9774
rect 36428 9884 37044 9940
rect 36428 9826 36484 9884
rect 36428 9774 36430 9826
rect 36482 9774 36484 9826
rect 36428 9762 36484 9774
rect 35756 9716 35812 9726
rect 35756 9266 35812 9660
rect 36540 9716 36596 9726
rect 36540 9622 36596 9660
rect 36764 9604 36820 9614
rect 36764 9602 36932 9604
rect 36764 9550 36766 9602
rect 36818 9550 36932 9602
rect 36764 9548 36932 9550
rect 36764 9538 36820 9548
rect 35756 9214 35758 9266
rect 35810 9214 35812 9266
rect 35756 9202 35812 9214
rect 36428 9492 36484 9502
rect 36428 9154 36484 9436
rect 36540 9268 36596 9278
rect 36540 9174 36596 9212
rect 36428 9102 36430 9154
rect 36482 9102 36484 9154
rect 36428 9090 36484 9102
rect 35980 9044 36036 9054
rect 35644 9042 35812 9044
rect 35644 8990 35646 9042
rect 35698 8990 35812 9042
rect 35644 8988 35812 8990
rect 35644 8978 35700 8988
rect 35308 8318 35310 8370
rect 35362 8318 35364 8370
rect 35308 8306 35364 8318
rect 35756 8484 35812 8988
rect 35980 9042 36372 9044
rect 35980 8990 35982 9042
rect 36034 8990 36372 9042
rect 35980 8988 36372 8990
rect 35980 8978 36036 8988
rect 36316 8484 36372 8988
rect 36540 8820 36596 8830
rect 36540 8726 36596 8764
rect 36428 8484 36484 8494
rect 36316 8482 36484 8484
rect 36316 8430 36430 8482
rect 36482 8430 36484 8482
rect 36316 8428 36484 8430
rect 35756 8370 35812 8428
rect 35756 8318 35758 8370
rect 35810 8318 35812 8370
rect 35756 8306 35812 8318
rect 36204 8258 36260 8270
rect 36204 8206 36206 8258
rect 36258 8206 36260 8258
rect 36204 7588 36260 8206
rect 36428 7812 36484 8428
rect 36764 8260 36820 8270
rect 36764 8166 36820 8204
rect 36876 8148 36932 9548
rect 36988 9044 37044 9884
rect 37212 9604 37268 9614
rect 37212 9268 37268 9548
rect 37324 9380 37380 13580
rect 38332 13186 38388 20132
rect 38668 20020 38724 20030
rect 38668 19926 38724 19964
rect 38892 19908 38948 20526
rect 39116 20578 39172 20590
rect 39116 20526 39118 20578
rect 39170 20526 39172 20578
rect 39116 20468 39172 20526
rect 39116 20402 39172 20412
rect 39116 19908 39172 19918
rect 38892 19906 39172 19908
rect 38892 19854 39118 19906
rect 39170 19854 39172 19906
rect 38892 19852 39172 19854
rect 38444 19458 38500 19470
rect 38444 19406 38446 19458
rect 38498 19406 38500 19458
rect 38444 18562 38500 19406
rect 38668 19236 38724 19246
rect 38444 18510 38446 18562
rect 38498 18510 38500 18562
rect 38444 18498 38500 18510
rect 38556 19180 38668 19236
rect 38556 18228 38612 19180
rect 38668 19170 38724 19180
rect 39004 19236 39060 19246
rect 39004 19142 39060 19180
rect 38668 19010 38724 19022
rect 38668 18958 38670 19010
rect 38722 18958 38724 19010
rect 38668 18452 38724 18958
rect 39116 18900 39172 19852
rect 39116 18834 39172 18844
rect 38892 18676 38948 18686
rect 38892 18582 38948 18620
rect 39228 18676 39284 18686
rect 38668 18358 38724 18396
rect 39004 18562 39060 18574
rect 39004 18510 39006 18562
rect 39058 18510 39060 18562
rect 38892 18338 38948 18350
rect 38892 18286 38894 18338
rect 38946 18286 38948 18338
rect 38556 18172 38724 18228
rect 38556 17554 38612 17566
rect 38556 17502 38558 17554
rect 38610 17502 38612 17554
rect 38556 16212 38612 17502
rect 38668 17106 38724 18172
rect 38892 17668 38948 18286
rect 39004 18340 39060 18510
rect 39004 18274 39060 18284
rect 38892 17602 38948 17612
rect 38668 17054 38670 17106
rect 38722 17054 38724 17106
rect 38668 17042 38724 17054
rect 39228 17444 39284 18620
rect 39340 18116 39396 20750
rect 39452 20356 39508 21420
rect 39452 20290 39508 20300
rect 39676 20244 39732 21644
rect 40124 21698 40180 21710
rect 40124 21646 40126 21698
rect 40178 21646 40180 21698
rect 40012 21586 40068 21598
rect 40012 21534 40014 21586
rect 40066 21534 40068 21586
rect 40012 21252 40068 21534
rect 40124 21476 40180 21646
rect 40124 21410 40180 21420
rect 40460 21362 40516 21374
rect 40460 21310 40462 21362
rect 40514 21310 40516 21362
rect 40460 21252 40516 21310
rect 40012 21196 40516 21252
rect 39900 20690 39956 20702
rect 39900 20638 39902 20690
rect 39954 20638 39956 20690
rect 39900 20580 39956 20638
rect 39900 20514 39956 20524
rect 39852 20412 40116 20422
rect 39908 20356 39956 20412
rect 40012 20356 40060 20412
rect 39852 20346 40116 20356
rect 39788 20244 39844 20254
rect 39676 20242 39844 20244
rect 39676 20190 39790 20242
rect 39842 20190 39844 20242
rect 39676 20188 39844 20190
rect 39564 20132 39620 20142
rect 39564 20038 39620 20076
rect 39676 20020 39732 20188
rect 39788 20178 39844 20188
rect 39564 19124 39620 19134
rect 39340 18050 39396 18060
rect 39452 19122 39620 19124
rect 39452 19070 39566 19122
rect 39618 19070 39620 19122
rect 39452 19068 39620 19070
rect 39452 18452 39508 19068
rect 39564 19058 39620 19068
rect 39676 19122 39732 19964
rect 39900 20018 39956 20030
rect 39900 19966 39902 20018
rect 39954 19966 39956 20018
rect 39900 19348 39956 19966
rect 39900 19282 39956 19292
rect 39676 19070 39678 19122
rect 39730 19070 39732 19122
rect 39676 19058 39732 19070
rect 39900 19012 39956 19050
rect 39900 18946 39956 18956
rect 40236 18900 40292 21196
rect 40348 20802 40404 20814
rect 40348 20750 40350 20802
rect 40402 20750 40404 20802
rect 40348 20132 40404 20750
rect 40348 20066 40404 20076
rect 40572 20130 40628 22428
rect 40796 22418 40852 22428
rect 40908 22372 40964 23100
rect 41916 23156 41972 23166
rect 41916 23062 41972 23100
rect 41020 22932 41076 22942
rect 41580 22932 41636 22942
rect 41020 22930 41636 22932
rect 41020 22878 41022 22930
rect 41074 22878 41582 22930
rect 41634 22878 41636 22930
rect 41020 22876 41636 22878
rect 41020 22866 41076 22876
rect 41580 22866 41636 22876
rect 40908 22240 40964 22316
rect 41580 22708 41636 22718
rect 41580 22148 41636 22652
rect 42476 22372 42532 22382
rect 41580 22146 41748 22148
rect 41580 22094 41582 22146
rect 41634 22094 41748 22146
rect 41580 22092 41748 22094
rect 41580 22082 41636 22092
rect 40684 21474 40740 21486
rect 40684 21422 40686 21474
rect 40738 21422 40740 21474
rect 40684 21362 40740 21422
rect 40684 21310 40686 21362
rect 40738 21310 40740 21362
rect 40684 21298 40740 21310
rect 41580 21028 41636 21038
rect 40684 21026 41636 21028
rect 40684 20974 41582 21026
rect 41634 20974 41636 21026
rect 40684 20972 41636 20974
rect 40684 20914 40740 20972
rect 40684 20862 40686 20914
rect 40738 20862 40740 20914
rect 40684 20850 40740 20862
rect 40572 20078 40574 20130
rect 40626 20078 40628 20130
rect 40460 19460 40516 19470
rect 40572 19460 40628 20078
rect 40908 20244 40964 20254
rect 40684 20020 40740 20030
rect 40684 19926 40740 19964
rect 40460 19458 40628 19460
rect 40460 19406 40462 19458
rect 40514 19406 40628 19458
rect 40460 19404 40628 19406
rect 40796 19794 40852 19806
rect 40796 19742 40798 19794
rect 40850 19742 40852 19794
rect 40460 19394 40516 19404
rect 40460 19236 40516 19246
rect 40516 19180 40740 19236
rect 40348 19124 40404 19134
rect 40348 19030 40404 19068
rect 40460 19122 40516 19180
rect 40460 19070 40462 19122
rect 40514 19070 40516 19122
rect 40460 19058 40516 19070
rect 39852 18844 40116 18854
rect 39908 18788 39956 18844
rect 40012 18788 40060 18844
rect 39852 18778 40116 18788
rect 40124 18676 40180 18686
rect 40236 18676 40292 18844
rect 40180 18620 40292 18676
rect 40572 19012 40628 19022
rect 40124 18610 40180 18620
rect 39340 17668 39396 17678
rect 39340 17574 39396 17612
rect 39228 17106 39284 17388
rect 39228 17054 39230 17106
rect 39282 17054 39284 17106
rect 39228 17042 39284 17054
rect 39452 17108 39508 18396
rect 40460 18452 40516 18462
rect 40460 18338 40516 18396
rect 40572 18450 40628 18956
rect 40572 18398 40574 18450
rect 40626 18398 40628 18450
rect 40572 18386 40628 18398
rect 40460 18286 40462 18338
rect 40514 18286 40516 18338
rect 40460 18274 40516 18286
rect 39788 18228 39844 18238
rect 39788 18134 39844 18172
rect 39676 17780 39732 17790
rect 39676 17686 39732 17724
rect 40236 17554 40292 17566
rect 40236 17502 40238 17554
rect 40290 17502 40292 17554
rect 39452 16884 39508 17052
rect 39564 17442 39620 17454
rect 39564 17390 39566 17442
rect 39618 17390 39620 17442
rect 39564 16996 39620 17390
rect 40236 17332 40292 17502
rect 40348 17444 40404 17454
rect 40348 17350 40404 17388
rect 40572 17444 40628 17454
rect 40572 17350 40628 17388
rect 39852 17276 40116 17286
rect 39908 17220 39956 17276
rect 40012 17220 40060 17276
rect 40236 17266 40292 17276
rect 39852 17210 40116 17220
rect 40684 17106 40740 19180
rect 40796 18452 40852 19742
rect 40796 18386 40852 18396
rect 40908 17668 40964 20188
rect 41580 20130 41636 20972
rect 41580 20078 41582 20130
rect 41634 20078 41636 20130
rect 41580 20066 41636 20078
rect 41020 19348 41076 19358
rect 41020 19010 41076 19292
rect 41580 19124 41636 19134
rect 41580 19030 41636 19068
rect 41020 18958 41022 19010
rect 41074 18958 41076 19010
rect 41020 18788 41076 18958
rect 41020 18722 41076 18732
rect 41692 18788 41748 22092
rect 42476 21698 42532 22316
rect 43036 22260 43092 22270
rect 43036 22166 43092 22204
rect 42476 21646 42478 21698
rect 42530 21646 42532 21698
rect 42476 21634 42532 21646
rect 42140 21586 42196 21598
rect 42140 21534 42142 21586
rect 42194 21534 42196 21586
rect 42028 21474 42084 21486
rect 42028 21422 42030 21474
rect 42082 21422 42084 21474
rect 41916 20916 41972 20926
rect 41916 20822 41972 20860
rect 41804 20132 41860 20142
rect 41804 20038 41860 20076
rect 41916 19908 41972 19918
rect 42028 19908 42084 21422
rect 42140 20690 42196 21534
rect 42140 20638 42142 20690
rect 42194 20638 42196 20690
rect 42140 20020 42196 20638
rect 42140 19954 42196 19964
rect 41916 19906 42084 19908
rect 41916 19854 41918 19906
rect 41970 19854 42084 19906
rect 41916 19852 42084 19854
rect 41916 19842 41972 19852
rect 42700 19348 42756 19358
rect 42700 19254 42756 19292
rect 42364 19122 42420 19134
rect 42364 19070 42366 19122
rect 42418 19070 42420 19122
rect 41692 18722 41748 18732
rect 41916 18788 41972 18798
rect 41580 18452 41636 18462
rect 40908 17612 41076 17668
rect 40908 17442 40964 17454
rect 40908 17390 40910 17442
rect 40962 17390 40964 17442
rect 40908 17332 40964 17390
rect 40908 17266 40964 17276
rect 40684 17054 40686 17106
rect 40738 17054 40740 17106
rect 40684 17042 40740 17054
rect 40908 17108 40964 17118
rect 40908 17014 40964 17052
rect 39564 16940 39732 16996
rect 39452 16828 39620 16884
rect 39564 16770 39620 16828
rect 39564 16718 39566 16770
rect 39618 16718 39620 16770
rect 39564 16706 39620 16718
rect 38780 16658 38836 16670
rect 38780 16606 38782 16658
rect 38834 16606 38836 16658
rect 38556 16156 38724 16212
rect 38444 16100 38500 16110
rect 38444 16006 38500 16044
rect 38668 15876 38724 16156
rect 38668 15810 38724 15820
rect 38780 15314 38836 16606
rect 39676 16658 39732 16940
rect 40124 16884 40180 16894
rect 40572 16884 40628 16894
rect 40124 16882 40628 16884
rect 40124 16830 40126 16882
rect 40178 16830 40574 16882
rect 40626 16830 40628 16882
rect 40124 16828 40628 16830
rect 40124 16818 40180 16828
rect 39676 16606 39678 16658
rect 39730 16606 39732 16658
rect 39004 16098 39060 16110
rect 39004 16046 39006 16098
rect 39058 16046 39060 16098
rect 39004 15876 39060 16046
rect 39004 15810 39060 15820
rect 39116 16100 39172 16110
rect 39116 15986 39172 16044
rect 39116 15934 39118 15986
rect 39170 15934 39172 15986
rect 38780 15262 38782 15314
rect 38834 15262 38836 15314
rect 38780 15250 38836 15262
rect 38892 15764 38948 15774
rect 38892 15204 38948 15708
rect 39116 15314 39172 15934
rect 39564 15988 39620 15998
rect 39564 15540 39620 15932
rect 39676 15986 39732 16606
rect 40572 16660 40628 16828
rect 40572 16594 40628 16604
rect 40460 16436 40516 16446
rect 40124 16212 40180 16222
rect 39900 16100 39956 16110
rect 39900 16006 39956 16044
rect 40124 16098 40180 16156
rect 40124 16046 40126 16098
rect 40178 16046 40180 16098
rect 40124 16034 40180 16046
rect 40236 16210 40292 16222
rect 40236 16158 40238 16210
rect 40290 16158 40292 16210
rect 40236 16100 40292 16158
rect 40236 16044 40404 16100
rect 39676 15934 39678 15986
rect 39730 15934 39732 15986
rect 39676 15922 39732 15934
rect 40236 15876 40292 15886
rect 40236 15782 40292 15820
rect 39852 15708 40116 15718
rect 39908 15652 39956 15708
rect 40012 15652 40060 15708
rect 40348 15652 40404 16044
rect 39852 15642 40116 15652
rect 40236 15596 40404 15652
rect 39676 15540 39732 15550
rect 39564 15538 39732 15540
rect 39564 15486 39678 15538
rect 39730 15486 39732 15538
rect 39564 15484 39732 15486
rect 39676 15474 39732 15484
rect 39116 15262 39118 15314
rect 39170 15262 39172 15314
rect 39116 15250 39172 15262
rect 38444 14530 38500 14542
rect 38444 14478 38446 14530
rect 38498 14478 38500 14530
rect 38444 13860 38500 14478
rect 38444 13794 38500 13804
rect 38892 13746 38948 15148
rect 39788 14980 39844 14990
rect 39788 14754 39844 14924
rect 39788 14702 39790 14754
rect 39842 14702 39844 14754
rect 39788 14690 39844 14702
rect 40236 14644 40292 15596
rect 40236 14578 40292 14588
rect 38892 13694 38894 13746
rect 38946 13694 38948 13746
rect 38892 13682 38948 13694
rect 39116 14532 39172 14542
rect 39116 14418 39172 14476
rect 39116 14366 39118 14418
rect 39170 14366 39172 14418
rect 39116 13634 39172 14366
rect 39900 14420 39956 14430
rect 39788 14308 39844 14346
rect 39900 14326 39956 14364
rect 40348 14420 40404 14430
rect 40348 14326 40404 14364
rect 39788 14242 39844 14252
rect 39852 14140 40116 14150
rect 39908 14084 39956 14140
rect 40012 14084 40060 14140
rect 39852 14074 40116 14084
rect 39676 13748 39732 13758
rect 39676 13654 39732 13692
rect 40236 13746 40292 13758
rect 40236 13694 40238 13746
rect 40290 13694 40292 13746
rect 39116 13582 39118 13634
rect 39170 13582 39172 13634
rect 39116 13570 39172 13582
rect 39900 13636 39956 13646
rect 38332 13134 38334 13186
rect 38386 13134 38388 13186
rect 38332 13122 38388 13134
rect 37884 13074 37940 13086
rect 37884 13022 37886 13074
rect 37938 13022 37940 13074
rect 37772 12962 37828 12974
rect 37772 12910 37774 12962
rect 37826 12910 37828 12962
rect 37772 12740 37828 12910
rect 37884 12852 37940 13022
rect 39900 12962 39956 13580
rect 39900 12910 39902 12962
rect 39954 12910 39956 12962
rect 39900 12852 39956 12910
rect 37884 12786 37940 12796
rect 39676 12796 39956 12852
rect 37772 12674 37828 12684
rect 39228 12180 39284 12190
rect 39116 12178 39284 12180
rect 39116 12126 39230 12178
rect 39282 12126 39284 12178
rect 39116 12124 39284 12126
rect 38556 12066 38612 12078
rect 38556 12014 38558 12066
rect 38610 12014 38612 12066
rect 38556 11172 38612 12014
rect 38556 11106 38612 11116
rect 39116 11172 39172 12124
rect 39228 12114 39284 12124
rect 38332 10612 38388 10622
rect 38220 10610 38388 10612
rect 38220 10558 38334 10610
rect 38386 10558 38388 10610
rect 38220 10556 38388 10558
rect 37436 9604 37492 9614
rect 37436 9510 37492 9548
rect 38220 9604 38276 10556
rect 38332 10546 38388 10556
rect 38668 10500 38724 10510
rect 38556 10444 38668 10500
rect 38556 9826 38612 10444
rect 38668 10406 38724 10444
rect 39116 10276 39172 11116
rect 39564 12066 39620 12078
rect 39564 12014 39566 12066
rect 39618 12014 39620 12066
rect 39564 11284 39620 12014
rect 39676 11954 39732 12796
rect 39852 12572 40116 12582
rect 39908 12516 39956 12572
rect 40012 12516 40060 12572
rect 39852 12506 40116 12516
rect 40236 12404 40292 13694
rect 40348 13748 40404 13758
rect 40348 12962 40404 13692
rect 40348 12910 40350 12962
rect 40402 12910 40404 12962
rect 40348 12898 40404 12910
rect 39676 11902 39678 11954
rect 39730 11902 39732 11954
rect 39676 11890 39732 11902
rect 40012 12348 40292 12404
rect 40348 12516 40404 12526
rect 40012 11394 40068 12348
rect 40124 12068 40180 12078
rect 40124 11508 40180 12012
rect 40124 11452 40292 11508
rect 40012 11342 40014 11394
rect 40066 11342 40068 11394
rect 40012 11330 40068 11342
rect 39676 11284 39732 11294
rect 39564 11282 39732 11284
rect 39564 11230 39678 11282
rect 39730 11230 39732 11282
rect 39564 11228 39732 11230
rect 39228 10610 39284 10622
rect 39228 10558 39230 10610
rect 39282 10558 39284 10610
rect 39228 10500 39284 10558
rect 39228 10434 39284 10444
rect 39116 10210 39172 10220
rect 38556 9774 38558 9826
rect 38610 9774 38612 9826
rect 38556 9762 38612 9774
rect 38892 9828 38948 9838
rect 39452 9828 39508 9838
rect 38892 9826 39508 9828
rect 38892 9774 38894 9826
rect 38946 9774 39454 9826
rect 39506 9774 39508 9826
rect 38892 9772 39508 9774
rect 38892 9762 38948 9772
rect 39452 9762 39508 9772
rect 37884 9492 37940 9502
rect 37324 9324 37492 9380
rect 37268 9212 37380 9268
rect 37212 9202 37268 9212
rect 37324 9154 37380 9212
rect 37324 9102 37326 9154
rect 37378 9102 37380 9154
rect 37324 9090 37380 9102
rect 37212 9044 37268 9054
rect 36988 9042 37268 9044
rect 36988 8990 37214 9042
rect 37266 8990 37268 9042
rect 36988 8988 37268 8990
rect 36876 8082 36932 8092
rect 36428 7746 36484 7756
rect 36540 7588 36596 7598
rect 36204 7586 36596 7588
rect 36204 7534 36542 7586
rect 36594 7534 36596 7586
rect 36204 7532 36596 7534
rect 35196 7298 35252 7308
rect 36316 7364 36372 7374
rect 36316 7270 36372 7308
rect 35532 6916 35588 6926
rect 35196 6914 35588 6916
rect 35196 6862 35534 6914
rect 35586 6862 35588 6914
rect 35196 6860 35588 6862
rect 34972 6692 35028 6702
rect 34972 6598 35028 6636
rect 34860 6580 34916 6590
rect 34860 6486 34916 6524
rect 34188 6468 34244 6478
rect 33852 5794 33908 5806
rect 33852 5742 33854 5794
rect 33906 5742 33908 5794
rect 32844 4450 33348 4452
rect 32844 4398 32846 4450
rect 32898 4398 33348 4450
rect 32844 4396 33348 4398
rect 33516 5122 33572 5134
rect 33516 5070 33518 5122
rect 33570 5070 33572 5122
rect 32844 4386 32900 4396
rect 32732 4246 32788 4284
rect 33516 3780 33572 5070
rect 33852 4452 33908 5742
rect 34188 5348 34244 6412
rect 35084 6468 35140 6478
rect 35084 6374 35140 6412
rect 35084 6020 35140 6030
rect 35084 5906 35140 5964
rect 35084 5854 35086 5906
rect 35138 5854 35140 5906
rect 35084 5842 35140 5854
rect 34188 5282 34244 5292
rect 34412 5794 34468 5806
rect 34412 5742 34414 5794
rect 34466 5742 34468 5794
rect 34076 5236 34132 5246
rect 34076 5142 34132 5180
rect 34412 5124 34468 5742
rect 34412 5058 34468 5068
rect 34860 5794 34916 5806
rect 34860 5742 34862 5794
rect 34914 5742 34916 5794
rect 34860 5124 34916 5742
rect 34860 5010 34916 5068
rect 35196 5348 35252 6860
rect 35532 6850 35588 6860
rect 35308 6690 35364 6702
rect 35308 6638 35310 6690
rect 35362 6638 35364 6690
rect 35308 6132 35364 6638
rect 36092 6580 36148 6590
rect 35980 6578 36148 6580
rect 35980 6526 36094 6578
rect 36146 6526 36148 6578
rect 35980 6524 36148 6526
rect 35980 6468 36036 6524
rect 36092 6514 36148 6524
rect 36428 6580 36484 7532
rect 36540 7522 36596 7532
rect 37212 7252 37268 8988
rect 37212 7186 37268 7196
rect 37324 8484 37380 8494
rect 36428 6486 36484 6524
rect 35420 6132 35476 6142
rect 35308 6130 35476 6132
rect 35308 6078 35422 6130
rect 35474 6078 35476 6130
rect 35308 6076 35476 6078
rect 35420 6066 35476 6076
rect 35196 5122 35252 5292
rect 35196 5070 35198 5122
rect 35250 5070 35252 5122
rect 35196 5058 35252 5070
rect 35532 5796 35588 5806
rect 35532 5236 35588 5740
rect 35980 5684 36036 6412
rect 36204 6466 36260 6478
rect 36204 6414 36206 6466
rect 36258 6414 36260 6466
rect 36204 6244 36260 6414
rect 36764 6466 36820 6478
rect 36764 6414 36766 6466
rect 36818 6414 36820 6466
rect 36764 6244 36820 6414
rect 36204 6188 36820 6244
rect 36204 6132 36260 6188
rect 35980 5618 36036 5628
rect 36092 6076 36260 6132
rect 36988 6132 37044 6142
rect 34860 4958 34862 5010
rect 34914 4958 34916 5010
rect 34860 4946 34916 4958
rect 33628 4340 33684 4350
rect 33628 4246 33684 4284
rect 33516 3714 33572 3724
rect 32172 3602 32228 3612
rect 32508 3556 32564 3566
rect 30940 3390 30942 3442
rect 30994 3390 30996 3442
rect 30940 3378 30996 3390
rect 31612 3444 31668 3482
rect 32508 3462 32564 3500
rect 31612 3378 31668 3388
rect 32396 3444 32452 3454
rect 32396 2324 32452 3388
rect 33180 3444 33236 3482
rect 33180 3378 33236 3388
rect 33516 3332 33572 3342
rect 33852 3332 33908 4396
rect 34076 4564 34132 4574
rect 34076 4338 34132 4508
rect 35532 4562 35588 5180
rect 35532 4510 35534 4562
rect 35586 4510 35588 4562
rect 35532 4498 35588 4510
rect 35644 4452 35700 4462
rect 35644 4358 35700 4396
rect 35308 4340 35364 4350
rect 34076 4286 34078 4338
rect 34130 4286 34132 4338
rect 34076 3444 34132 4286
rect 35084 4338 35364 4340
rect 35084 4286 35310 4338
rect 35362 4286 35364 4338
rect 35084 4284 35364 4286
rect 34412 4228 34468 4238
rect 34188 3780 34244 3790
rect 34188 3686 34244 3724
rect 34300 3556 34356 3566
rect 34412 3556 34468 4172
rect 34300 3554 34468 3556
rect 34300 3502 34302 3554
rect 34354 3502 34468 3554
rect 34300 3500 34468 3502
rect 34860 3556 34916 3566
rect 34300 3490 34356 3500
rect 34188 3444 34244 3454
rect 34076 3442 34244 3444
rect 34076 3390 34190 3442
rect 34242 3390 34244 3442
rect 34076 3388 34244 3390
rect 34188 3378 34244 3388
rect 33516 3330 33908 3332
rect 33516 3278 33518 3330
rect 33570 3278 33908 3330
rect 33516 3276 33908 3278
rect 33516 3266 33572 3276
rect 32396 2268 32564 2324
rect 28812 1250 28868 1260
rect 30380 2156 30660 2212
rect 30380 800 30436 2156
rect 32508 800 32564 2268
rect 34860 2212 34916 3500
rect 34636 2156 34916 2212
rect 34636 800 34692 2156
rect 35084 1652 35140 4284
rect 35308 4274 35364 4284
rect 35980 3556 36036 3566
rect 35980 3462 36036 3500
rect 35196 3332 35252 3342
rect 35196 3330 35364 3332
rect 35196 3278 35198 3330
rect 35250 3278 35364 3330
rect 35196 3276 35364 3278
rect 35196 3266 35252 3276
rect 35084 1586 35140 1596
rect 35308 2772 35364 3276
rect 35308 1428 35364 2716
rect 36092 2212 36148 6076
rect 36316 6018 36372 6030
rect 36316 5966 36318 6018
rect 36370 5966 36372 6018
rect 36204 5906 36260 5918
rect 36204 5854 36206 5906
rect 36258 5854 36260 5906
rect 36204 5684 36260 5854
rect 36316 5796 36372 5966
rect 36316 5730 36372 5740
rect 36540 6020 36596 6030
rect 36204 5618 36260 5628
rect 36540 5010 36596 5964
rect 36876 5796 36932 5806
rect 36876 5702 36932 5740
rect 36540 4958 36542 5010
rect 36594 4958 36596 5010
rect 36540 4946 36596 4958
rect 36764 5012 36820 5022
rect 36764 4338 36820 4956
rect 36988 4452 37044 6076
rect 37324 6130 37380 8428
rect 37436 7140 37492 9324
rect 37884 9266 37940 9436
rect 37884 9214 37886 9266
rect 37938 9214 37940 9266
rect 37548 9042 37604 9054
rect 37548 8990 37550 9042
rect 37602 8990 37604 9042
rect 37548 8932 37604 8990
rect 37548 8866 37604 8876
rect 37884 8484 37940 9214
rect 37884 8418 37940 8428
rect 38108 8372 38164 8382
rect 38220 8372 38276 9548
rect 38668 9604 38724 9614
rect 39564 9604 39620 11228
rect 39676 11218 39732 11228
rect 39788 11172 39844 11210
rect 39788 11106 39844 11116
rect 39852 11004 40116 11014
rect 39908 10948 39956 11004
rect 40012 10948 40060 11004
rect 39852 10938 40116 10948
rect 40124 10612 40180 10622
rect 40124 10518 40180 10556
rect 40012 10500 40068 10510
rect 39900 10164 39956 10174
rect 39900 9826 39956 10108
rect 39900 9774 39902 9826
rect 39954 9774 39956 9826
rect 39900 9762 39956 9774
rect 40012 9828 40068 10444
rect 40124 9828 40180 9838
rect 40012 9826 40180 9828
rect 40012 9774 40126 9826
rect 40178 9774 40180 9826
rect 40012 9772 40180 9774
rect 40124 9762 40180 9772
rect 38668 9510 38724 9548
rect 39452 9548 39620 9604
rect 40012 9604 40068 9642
rect 38108 8370 38276 8372
rect 38108 8318 38110 8370
rect 38162 8318 38276 8370
rect 38108 8316 38276 8318
rect 38332 8930 38388 8942
rect 38332 8878 38334 8930
rect 38386 8878 38388 8930
rect 38108 8306 38164 8316
rect 37548 8258 37604 8270
rect 37548 8206 37550 8258
rect 37602 8206 37604 8258
rect 37548 7364 37604 8206
rect 37772 8260 37828 8270
rect 37772 8166 37828 8204
rect 38220 8148 38276 8158
rect 38220 8054 38276 8092
rect 37996 8034 38052 8046
rect 37996 7982 37998 8034
rect 38050 7982 38052 8034
rect 37772 7812 37828 7822
rect 37772 7474 37828 7756
rect 37772 7422 37774 7474
rect 37826 7422 37828 7474
rect 37772 7410 37828 7422
rect 37548 7298 37604 7308
rect 37660 7252 37716 7262
rect 37436 7084 37604 7140
rect 37436 6468 37492 6478
rect 37436 6374 37492 6412
rect 37324 6078 37326 6130
rect 37378 6078 37380 6130
rect 37324 5684 37380 6078
rect 37324 5618 37380 5628
rect 36988 4386 37044 4396
rect 36764 4286 36766 4338
rect 36818 4286 36820 4338
rect 36764 4274 36820 4286
rect 36204 4228 36260 4238
rect 36204 4134 36260 4172
rect 37100 4228 37156 4238
rect 37100 4134 37156 4172
rect 36764 3556 36820 3566
rect 36428 3444 36484 3482
rect 36428 3378 36484 3388
rect 36092 2146 36148 2156
rect 35308 1362 35364 1372
rect 36764 800 36820 3500
rect 37100 3556 37156 3566
rect 37100 3462 37156 3500
rect 37436 3330 37492 3342
rect 37436 3278 37438 3330
rect 37490 3278 37492 3330
rect 37436 2772 37492 3278
rect 37436 2324 37492 2716
rect 37436 2258 37492 2268
rect 37548 868 37604 7084
rect 37660 6468 37716 7196
rect 37884 6468 37940 6478
rect 37660 6402 37716 6412
rect 37772 6466 37940 6468
rect 37772 6414 37886 6466
rect 37938 6414 37940 6466
rect 37772 6412 37940 6414
rect 37772 5796 37828 6412
rect 37884 6402 37940 6412
rect 37996 6020 38052 7982
rect 38332 7252 38388 8878
rect 39452 8428 39508 9548
rect 40012 9538 40068 9548
rect 39852 9436 40116 9446
rect 39908 9380 39956 9436
rect 40012 9380 40060 9436
rect 39852 9370 40116 9380
rect 39228 8372 39508 8428
rect 39564 9268 39620 9278
rect 38444 7364 38500 7374
rect 38444 7270 38500 7308
rect 38332 7186 38388 7196
rect 37996 5954 38052 5964
rect 38892 7028 38948 7038
rect 38668 5908 38724 5918
rect 38668 5814 38724 5852
rect 37660 5794 37828 5796
rect 37660 5742 37774 5794
rect 37826 5742 37828 5794
rect 37660 5740 37828 5742
rect 37660 5348 37716 5740
rect 37772 5730 37828 5740
rect 37660 1652 37716 5292
rect 38108 5124 38164 5134
rect 38556 5124 38612 5134
rect 37996 5068 38108 5124
rect 37772 4898 37828 4910
rect 37772 4846 37774 4898
rect 37826 4846 37828 4898
rect 37772 4564 37828 4846
rect 37772 4498 37828 4508
rect 37884 4900 37940 4910
rect 37884 4562 37940 4844
rect 37884 4510 37886 4562
rect 37938 4510 37940 4562
rect 37884 4498 37940 4510
rect 37772 4340 37828 4350
rect 37996 4340 38052 5068
rect 38108 5030 38164 5068
rect 38220 5122 38612 5124
rect 38220 5070 38558 5122
rect 38610 5070 38612 5122
rect 38220 5068 38612 5070
rect 38108 4564 38164 4574
rect 38220 4564 38276 5068
rect 38556 5058 38612 5068
rect 38892 5124 38948 6972
rect 39116 6020 39172 6030
rect 39228 6020 39284 8372
rect 39116 6018 39284 6020
rect 39116 5966 39118 6018
rect 39170 5966 39284 6018
rect 39116 5964 39284 5966
rect 39340 7362 39396 7374
rect 39340 7310 39342 7362
rect 39394 7310 39396 7362
rect 39340 6580 39396 7310
rect 39564 7140 39620 9212
rect 40012 9156 40068 9166
rect 40012 9062 40068 9100
rect 39852 7868 40116 7878
rect 39908 7812 39956 7868
rect 40012 7812 40060 7868
rect 39852 7802 40116 7812
rect 40012 7700 40068 7710
rect 40236 7700 40292 11452
rect 40348 9604 40404 12460
rect 40460 12292 40516 16380
rect 40908 16212 40964 16222
rect 41020 16212 41076 17612
rect 41580 16322 41636 18396
rect 41804 18340 41860 18350
rect 41692 17780 41748 17790
rect 41692 17686 41748 17724
rect 41804 17554 41860 18284
rect 41804 17502 41806 17554
rect 41858 17502 41860 17554
rect 41804 17108 41860 17502
rect 41804 17042 41860 17052
rect 41580 16270 41582 16322
rect 41634 16270 41636 16322
rect 41580 16258 41636 16270
rect 41804 16884 41860 16894
rect 40908 16210 41524 16212
rect 40908 16158 40910 16210
rect 40962 16158 41524 16210
rect 40908 16156 41524 16158
rect 40908 16146 40964 16156
rect 41468 15988 41524 16156
rect 41580 15988 41636 15998
rect 41468 15986 41636 15988
rect 41468 15934 41582 15986
rect 41634 15934 41636 15986
rect 41468 15932 41636 15934
rect 41580 15922 41636 15932
rect 41692 15986 41748 15998
rect 41692 15934 41694 15986
rect 41746 15934 41748 15986
rect 41692 15876 41748 15934
rect 41692 15810 41748 15820
rect 40572 15204 40628 15214
rect 40572 14418 40628 15148
rect 41804 15148 41860 16828
rect 41916 16324 41972 18732
rect 42364 18564 42420 19070
rect 42588 19012 42644 19022
rect 42588 18918 42644 18956
rect 42252 18452 42308 18462
rect 42252 18358 42308 18396
rect 42364 18226 42420 18508
rect 42588 18340 42644 18350
rect 42588 18246 42644 18284
rect 42364 18174 42366 18226
rect 42418 18174 42420 18226
rect 42364 18162 42420 18174
rect 42588 18116 42644 18126
rect 42028 17554 42084 17566
rect 42028 17502 42030 17554
rect 42082 17502 42084 17554
rect 42028 17444 42084 17502
rect 42028 16996 42084 17388
rect 42028 16930 42084 16940
rect 42476 16996 42532 17006
rect 42476 16902 42532 16940
rect 41916 16258 41972 16268
rect 42028 16772 42084 16782
rect 42028 16548 42084 16716
rect 42028 16212 42084 16492
rect 42140 16212 42196 16222
rect 42028 16210 42196 16212
rect 42028 16158 42142 16210
rect 42194 16158 42196 16210
rect 42028 16156 42196 16158
rect 42140 16146 42196 16156
rect 42476 15316 42532 15326
rect 42476 15148 42532 15260
rect 41804 15092 41972 15148
rect 41916 14756 41972 15092
rect 41916 14690 41972 14700
rect 42028 15092 42084 15102
rect 40684 14532 40740 14542
rect 40684 14438 40740 14476
rect 40572 14366 40574 14418
rect 40626 14366 40628 14418
rect 40572 14354 40628 14366
rect 41580 14308 41636 14318
rect 40684 14196 40740 14206
rect 40684 13970 40740 14140
rect 40684 13918 40686 13970
rect 40738 13918 40740 13970
rect 40684 13906 40740 13918
rect 40572 13748 40628 13758
rect 40572 13654 40628 13692
rect 40796 13746 40852 13758
rect 40796 13694 40798 13746
rect 40850 13694 40852 13746
rect 40796 13636 40852 13694
rect 40796 13570 40852 13580
rect 41580 13524 41636 14252
rect 41580 13458 41636 13468
rect 42028 13076 42084 15036
rect 42364 15092 42532 15148
rect 42252 14644 42308 14654
rect 42364 14644 42420 15092
rect 42252 14642 42420 14644
rect 42252 14590 42254 14642
rect 42306 14590 42420 14642
rect 42252 14588 42420 14590
rect 42476 14644 42532 14654
rect 42252 14308 42308 14588
rect 42476 14418 42532 14588
rect 42476 14366 42478 14418
rect 42530 14366 42532 14418
rect 42476 14354 42532 14366
rect 42252 14242 42308 14252
rect 42588 13186 42644 18060
rect 42700 15876 42756 15886
rect 42700 15782 42756 15820
rect 43036 15316 43092 15326
rect 43036 15222 43092 15260
rect 43148 15202 43204 15214
rect 43148 15150 43150 15202
rect 43202 15150 43204 15202
rect 43148 13970 43204 15150
rect 43260 15148 43316 26684
rect 43932 26516 43988 26526
rect 43372 26404 43428 26414
rect 43372 25618 43428 26348
rect 43820 26404 43876 26414
rect 43820 26310 43876 26348
rect 43932 26402 43988 26460
rect 43932 26350 43934 26402
rect 43986 26350 43988 26402
rect 43932 26338 43988 26350
rect 44044 26292 44100 27022
rect 44604 27074 44660 27086
rect 44604 27022 44606 27074
rect 44658 27022 44660 27074
rect 44604 26908 44660 27022
rect 45052 27076 45108 27086
rect 44604 26852 44772 26908
rect 44044 26226 44100 26236
rect 44380 26404 44436 26414
rect 43372 25566 43374 25618
rect 43426 25566 43428 25618
rect 43372 25554 43428 25566
rect 43820 26066 43876 26078
rect 43820 26014 43822 26066
rect 43874 26014 43876 26066
rect 43484 25506 43540 25518
rect 43484 25454 43486 25506
rect 43538 25454 43540 25506
rect 43484 24836 43540 25454
rect 43820 25506 43876 26014
rect 43820 25454 43822 25506
rect 43874 25454 43876 25506
rect 43820 25442 43876 25454
rect 44380 25508 44436 26348
rect 44492 26292 44548 26302
rect 44492 26198 44548 26236
rect 44380 24948 44436 25452
rect 44716 26066 44772 26852
rect 45052 26514 45108 27020
rect 45500 27074 45556 27132
rect 45500 27022 45502 27074
rect 45554 27022 45556 27074
rect 45500 27010 45556 27022
rect 45724 27074 45780 27916
rect 46284 27972 46340 27982
rect 46284 27878 46340 27916
rect 46060 27858 46116 27870
rect 46060 27806 46062 27858
rect 46114 27806 46116 27858
rect 45948 27636 46004 27646
rect 45948 27298 46004 27580
rect 45948 27246 45950 27298
rect 46002 27246 46004 27298
rect 45948 27234 46004 27246
rect 45724 27022 45726 27074
rect 45778 27022 45780 27074
rect 45724 26908 45780 27022
rect 46060 27076 46116 27806
rect 46620 27860 46676 27870
rect 46620 27766 46676 27804
rect 46508 27748 46564 27758
rect 46508 27654 46564 27692
rect 46844 27636 46900 27646
rect 46060 26982 46116 27020
rect 46284 27076 46340 27086
rect 45724 26852 45892 26908
rect 45052 26462 45054 26514
rect 45106 26462 45108 26514
rect 45052 26450 45108 26462
rect 45500 26516 45556 26526
rect 45500 26422 45556 26460
rect 44716 26014 44718 26066
rect 44770 26014 44772 26066
rect 44604 25396 44660 25406
rect 44492 24948 44548 24958
rect 44380 24946 44548 24948
rect 44380 24894 44494 24946
rect 44546 24894 44548 24946
rect 44380 24892 44548 24894
rect 44492 24882 44548 24892
rect 44604 24946 44660 25340
rect 44604 24894 44606 24946
rect 44658 24894 44660 24946
rect 44604 24882 44660 24894
rect 43484 24704 43540 24780
rect 44044 24836 44100 24846
rect 44044 24742 44100 24780
rect 44268 24722 44324 24734
rect 44268 24670 44270 24722
rect 44322 24670 44324 24722
rect 44268 24612 44324 24670
rect 44268 24546 44324 24556
rect 44716 24050 44772 26014
rect 44940 25508 44996 25518
rect 44940 24946 44996 25452
rect 45836 25506 45892 26852
rect 46284 26850 46340 27020
rect 46284 26798 46286 26850
rect 46338 26798 46340 26850
rect 46284 26786 46340 26798
rect 45836 25454 45838 25506
rect 45890 25454 45892 25506
rect 45836 25442 45892 25454
rect 45500 25396 45556 25406
rect 45500 25302 45556 25340
rect 45612 25284 45668 25294
rect 45612 25190 45668 25228
rect 44940 24894 44942 24946
rect 44994 24894 44996 24946
rect 44940 24882 44996 24894
rect 46844 24946 46900 27580
rect 47404 26852 47460 33180
rect 48412 33012 48468 33022
rect 48076 32788 48132 32798
rect 48076 32694 48132 32732
rect 47628 32562 47684 32574
rect 47628 32510 47630 32562
rect 47682 32510 47684 32562
rect 47628 31780 47684 32510
rect 47628 31648 47684 31724
rect 47516 31556 47572 31566
rect 47516 31462 47572 31500
rect 47852 31556 47908 31566
rect 47852 30324 47908 31500
rect 48076 31556 48132 31566
rect 48076 31462 48132 31500
rect 48412 31218 48468 32956
rect 48412 31166 48414 31218
rect 48466 31166 48468 31218
rect 48412 31154 48468 31166
rect 48748 30994 48804 31006
rect 48748 30942 48750 30994
rect 48802 30942 48804 30994
rect 48300 30324 48356 30334
rect 47852 30322 48356 30324
rect 47852 30270 47854 30322
rect 47906 30270 48302 30322
rect 48354 30270 48356 30322
rect 47852 30268 48356 30270
rect 47852 30258 47908 30268
rect 48300 30258 48356 30268
rect 48748 30324 48804 30942
rect 48748 30258 48804 30268
rect 47740 30100 47796 30110
rect 47740 30006 47796 30044
rect 48188 29314 48244 29326
rect 48188 29262 48190 29314
rect 48242 29262 48244 29314
rect 48188 28756 48244 29262
rect 48412 29204 48468 29214
rect 48188 28690 48244 28700
rect 48300 29202 48468 29204
rect 48300 29150 48414 29202
rect 48466 29150 48468 29202
rect 48300 29148 48468 29150
rect 48076 28644 48132 28654
rect 48076 27298 48132 28588
rect 48300 28644 48356 29148
rect 48412 29138 48468 29148
rect 48748 29204 48804 29214
rect 48748 29110 48804 29148
rect 48300 28550 48356 28588
rect 48412 28756 48468 28766
rect 48412 28530 48468 28700
rect 48636 28644 48692 28654
rect 48636 28550 48692 28588
rect 48412 28478 48414 28530
rect 48466 28478 48468 28530
rect 48076 27246 48078 27298
rect 48130 27246 48132 27298
rect 48076 27234 48132 27246
rect 48300 27300 48356 27310
rect 48412 27300 48468 28478
rect 48300 27298 48468 27300
rect 48300 27246 48302 27298
rect 48354 27246 48468 27298
rect 48300 27244 48468 27246
rect 48748 27748 48804 27758
rect 48748 27298 48804 27692
rect 48748 27246 48750 27298
rect 48802 27246 48804 27298
rect 48300 27234 48356 27244
rect 48748 27234 48804 27246
rect 48524 27076 48580 27086
rect 48524 26982 48580 27020
rect 48972 27074 49028 27086
rect 48972 27022 48974 27074
rect 49026 27022 49028 27074
rect 48972 26908 49028 27022
rect 47404 25732 47460 26796
rect 48860 26852 49028 26908
rect 48748 26516 48804 26526
rect 48860 26516 48916 26852
rect 48748 26514 48916 26516
rect 48748 26462 48750 26514
rect 48802 26462 48916 26514
rect 48748 26460 48916 26462
rect 49196 26740 49252 34638
rect 49512 33740 49776 33750
rect 49568 33684 49616 33740
rect 49672 33684 49720 33740
rect 49512 33674 49776 33684
rect 49308 33458 49364 33470
rect 49308 33406 49310 33458
rect 49362 33406 49364 33458
rect 49308 31780 49364 33406
rect 49644 33348 49700 33358
rect 49644 33254 49700 33292
rect 49868 33346 49924 35422
rect 49868 33294 49870 33346
rect 49922 33294 49924 33346
rect 49868 33282 49924 33294
rect 49980 34914 50036 34926
rect 49980 34862 49982 34914
rect 50034 34862 50036 34914
rect 49980 34692 50036 34862
rect 49980 33124 50036 34636
rect 50316 34692 50372 34702
rect 50316 34598 50372 34636
rect 50316 34020 50372 34030
rect 50316 34018 50484 34020
rect 50316 33966 50318 34018
rect 50370 33966 50484 34018
rect 50316 33964 50484 33966
rect 50316 33954 50372 33964
rect 50428 33572 50484 33964
rect 50540 33908 50596 35532
rect 50876 34916 50932 34926
rect 50876 34822 50932 34860
rect 51772 34804 51828 34814
rect 51660 34802 51828 34804
rect 51660 34750 51774 34802
rect 51826 34750 51828 34802
rect 51660 34748 51828 34750
rect 51212 34690 51268 34702
rect 51212 34638 51214 34690
rect 51266 34638 51268 34690
rect 51212 34468 51268 34638
rect 51212 34402 51268 34412
rect 51548 34244 51604 34254
rect 50988 34242 51604 34244
rect 50988 34190 51550 34242
rect 51602 34190 51604 34242
rect 50988 34188 51604 34190
rect 50652 34132 50708 34142
rect 50988 34132 51044 34188
rect 51548 34178 51604 34188
rect 50652 34130 51044 34132
rect 50652 34078 50654 34130
rect 50706 34078 51044 34130
rect 50652 34076 51044 34078
rect 50652 34066 50708 34076
rect 51100 34020 51156 34030
rect 51660 34020 51716 34748
rect 51772 34738 51828 34748
rect 51884 34356 51940 35532
rect 51996 35698 52052 35710
rect 51996 35646 51998 35698
rect 52050 35646 52052 35698
rect 51996 34692 52052 35646
rect 52108 34804 52164 34814
rect 52220 34804 52276 35868
rect 52780 36370 52836 36382
rect 52780 36318 52782 36370
rect 52834 36318 52836 36370
rect 52780 35812 52836 36318
rect 52780 35746 52836 35756
rect 53116 36258 53172 36270
rect 53116 36206 53118 36258
rect 53170 36206 53172 36258
rect 53116 35924 53172 36206
rect 53116 35700 53172 35868
rect 53116 35634 53172 35644
rect 53340 35924 53396 35934
rect 53564 35924 53620 36428
rect 53676 36418 53732 36428
rect 57708 36484 57764 37436
rect 58380 36596 58436 39200
rect 60844 39060 60900 39200
rect 61180 39060 61236 39228
rect 60844 39004 61236 39060
rect 58380 36530 58436 36540
rect 58828 36596 58884 36606
rect 58828 36502 58884 36540
rect 61740 36594 61796 39228
rect 63280 39200 63392 40000
rect 65744 39200 65856 40000
rect 66108 39228 66500 39284
rect 61740 36542 61742 36594
rect 61794 36542 61796 36594
rect 61740 36530 61796 36542
rect 63196 37604 63252 37614
rect 57708 36482 58212 36484
rect 57708 36430 57710 36482
rect 57762 36430 58212 36482
rect 57708 36428 58212 36430
rect 57708 36418 57764 36428
rect 53340 35922 53620 35924
rect 53340 35870 53342 35922
rect 53394 35870 53620 35922
rect 53340 35868 53620 35870
rect 52556 35588 52612 35598
rect 52556 35494 52612 35532
rect 52108 34802 52276 34804
rect 52108 34750 52110 34802
rect 52162 34750 52276 34802
rect 52108 34748 52276 34750
rect 52108 34738 52164 34748
rect 51996 34580 52052 34636
rect 51996 34524 52276 34580
rect 51884 34300 52052 34356
rect 51100 34018 51716 34020
rect 51100 33966 51102 34018
rect 51154 33966 51716 34018
rect 51100 33964 51716 33966
rect 51772 34242 51828 34254
rect 51772 34190 51774 34242
rect 51826 34190 51828 34242
rect 51100 33954 51156 33964
rect 50540 33852 50932 33908
rect 50428 33516 50596 33572
rect 49756 33068 50036 33124
rect 50092 33348 50148 33358
rect 49756 32674 49812 33068
rect 49756 32622 49758 32674
rect 49810 32622 49812 32674
rect 49756 32610 49812 32622
rect 49868 32786 49924 32798
rect 49868 32734 49870 32786
rect 49922 32734 49924 32786
rect 49532 32564 49588 32574
rect 49532 32470 49588 32508
rect 49512 32172 49776 32182
rect 49568 32116 49616 32172
rect 49672 32116 49720 32172
rect 49512 32106 49776 32116
rect 49308 31714 49364 31724
rect 49756 31780 49812 31790
rect 49868 31780 49924 32734
rect 50092 32674 50148 33292
rect 50428 33348 50484 33358
rect 50540 33348 50596 33516
rect 50764 33348 50820 33358
rect 50540 33346 50820 33348
rect 50540 33294 50766 33346
rect 50818 33294 50820 33346
rect 50540 33292 50820 33294
rect 50876 33348 50932 33852
rect 51772 33460 51828 34190
rect 51884 34132 51940 34142
rect 51884 34038 51940 34076
rect 51548 33404 51828 33460
rect 50988 33348 51044 33358
rect 50876 33292 50988 33348
rect 50428 33254 50484 33292
rect 50652 33124 50708 33134
rect 50652 32786 50708 33068
rect 50652 32734 50654 32786
rect 50706 32734 50708 32786
rect 50652 32722 50708 32734
rect 50764 32788 50820 33292
rect 50988 33124 51044 33292
rect 51548 33236 51604 33404
rect 51548 33170 51604 33180
rect 51772 33236 51828 33246
rect 51772 33142 51828 33180
rect 50988 33058 51044 33068
rect 51436 33122 51492 33134
rect 51436 33070 51438 33122
rect 51490 33070 51492 33122
rect 50764 32722 50820 32732
rect 50092 32622 50094 32674
rect 50146 32622 50148 32674
rect 50092 32610 50148 32622
rect 51436 32450 51492 33070
rect 51660 33124 51716 33134
rect 51660 33030 51716 33068
rect 51436 32398 51438 32450
rect 51490 32398 51492 32450
rect 51436 32386 51492 32398
rect 51548 32562 51604 32574
rect 51548 32510 51550 32562
rect 51602 32510 51604 32562
rect 51548 31948 51604 32510
rect 51996 31948 52052 34300
rect 52220 34244 52276 34524
rect 52444 34244 52500 34254
rect 52220 34242 52500 34244
rect 52220 34190 52446 34242
rect 52498 34190 52500 34242
rect 52220 34188 52500 34190
rect 52444 34178 52500 34188
rect 52556 34242 52612 34254
rect 52556 34190 52558 34242
rect 52610 34190 52612 34242
rect 52556 33348 52612 34190
rect 52780 34132 52836 34142
rect 52780 34038 52836 34076
rect 52556 33282 52612 33292
rect 53116 34018 53172 34030
rect 53116 33966 53118 34018
rect 53170 33966 53172 34018
rect 53116 33348 53172 33966
rect 53116 33282 53172 33292
rect 52332 33236 52388 33246
rect 52332 33122 52388 33180
rect 52332 33070 52334 33122
rect 52386 33070 52388 33122
rect 52220 32676 52276 32686
rect 52220 32582 52276 32620
rect 52332 32340 52388 33070
rect 52332 32274 52388 32284
rect 52780 33124 52836 33134
rect 51436 31892 51604 31948
rect 51660 31892 52052 31948
rect 49756 31778 49924 31780
rect 49756 31726 49758 31778
rect 49810 31726 49924 31778
rect 49756 31724 49924 31726
rect 49980 31780 50036 31790
rect 50036 31724 50260 31780
rect 49756 31108 49812 31724
rect 49980 31686 50036 31724
rect 49756 31042 49812 31052
rect 50204 30996 50260 31724
rect 51100 31668 51156 31678
rect 51100 31574 51156 31612
rect 50316 31556 50372 31566
rect 51212 31556 51268 31566
rect 50316 31554 50596 31556
rect 50316 31502 50318 31554
rect 50370 31502 50596 31554
rect 50316 31500 50596 31502
rect 50316 31490 50372 31500
rect 50428 31108 50484 31118
rect 50428 31014 50484 31052
rect 50316 30996 50372 31006
rect 50204 30994 50372 30996
rect 50204 30942 50318 30994
rect 50370 30942 50372 30994
rect 50204 30940 50372 30942
rect 50316 30930 50372 30940
rect 49512 30604 49776 30614
rect 49568 30548 49616 30604
rect 49672 30548 49720 30604
rect 49512 30538 49776 30548
rect 49756 30324 49812 30334
rect 49756 30230 49812 30268
rect 50540 30322 50596 31500
rect 50988 30882 51044 30894
rect 50988 30830 50990 30882
rect 51042 30830 51044 30882
rect 50988 30660 51044 30830
rect 50988 30594 51044 30604
rect 50540 30270 50542 30322
rect 50594 30270 50596 30322
rect 50428 30210 50484 30222
rect 50428 30158 50430 30210
rect 50482 30158 50484 30210
rect 50428 29652 50484 30158
rect 50316 29596 50428 29652
rect 49644 29428 49700 29438
rect 49644 29334 49700 29372
rect 50204 29426 50260 29438
rect 50204 29374 50206 29426
rect 50258 29374 50260 29426
rect 49868 29204 49924 29214
rect 49512 29036 49776 29046
rect 49568 28980 49616 29036
rect 49672 28980 49720 29036
rect 49512 28970 49776 28980
rect 49868 28642 49924 29148
rect 49868 28590 49870 28642
rect 49922 28590 49924 28642
rect 49868 28578 49924 28590
rect 49868 27858 49924 27870
rect 49868 27806 49870 27858
rect 49922 27806 49924 27858
rect 49756 27746 49812 27758
rect 49756 27694 49758 27746
rect 49810 27694 49812 27746
rect 49756 27636 49812 27694
rect 49868 27748 49924 27806
rect 49868 27682 49924 27692
rect 50204 27748 50260 29374
rect 50316 28642 50372 29596
rect 50428 29586 50484 29596
rect 50316 28590 50318 28642
rect 50370 28590 50372 28642
rect 50316 28578 50372 28590
rect 50428 29314 50484 29326
rect 50428 29262 50430 29314
rect 50482 29262 50484 29314
rect 50428 28530 50484 29262
rect 50428 28478 50430 28530
rect 50482 28478 50484 28530
rect 50428 28466 50484 28478
rect 50540 28756 50596 30270
rect 51100 29652 51156 29662
rect 51100 29558 51156 29596
rect 50540 28530 50596 28700
rect 50540 28478 50542 28530
rect 50594 28478 50596 28530
rect 50540 28466 50596 28478
rect 49756 27570 49812 27580
rect 50204 27634 50260 27692
rect 50204 27582 50206 27634
rect 50258 27582 50260 27634
rect 50204 27570 50260 27582
rect 49512 27468 49776 27478
rect 49568 27412 49616 27468
rect 49672 27412 49720 27468
rect 49512 27402 49776 27412
rect 49420 27076 49476 27086
rect 49420 27074 49700 27076
rect 49420 27022 49422 27074
rect 49474 27022 49700 27074
rect 49420 27020 49700 27022
rect 49420 27010 49476 27020
rect 49308 26964 49364 26974
rect 49308 26852 49364 26908
rect 49420 26852 49476 26862
rect 49308 26850 49476 26852
rect 49308 26798 49422 26850
rect 49474 26798 49476 26850
rect 49308 26796 49476 26798
rect 49420 26786 49476 26796
rect 48748 26450 48804 26460
rect 48188 26404 48244 26414
rect 48188 26180 48244 26348
rect 49196 26292 49252 26684
rect 49644 26514 49700 27020
rect 49644 26462 49646 26514
rect 49698 26462 49700 26514
rect 49644 26450 49700 26462
rect 49756 26404 49812 26414
rect 49756 26310 49812 26348
rect 50428 26402 50484 26414
rect 50428 26350 50430 26402
rect 50482 26350 50484 26402
rect 49196 26226 49252 26236
rect 50428 26292 50484 26350
rect 50428 26226 50484 26236
rect 50764 26292 50820 26302
rect 50764 26198 50820 26236
rect 47404 25666 47460 25676
rect 48076 26178 48244 26180
rect 48076 26126 48190 26178
rect 48242 26126 48244 26178
rect 48076 26124 48244 26126
rect 46844 24894 46846 24946
rect 46898 24894 46900 24946
rect 46844 24882 46900 24894
rect 48076 24834 48132 26124
rect 48188 26114 48244 26124
rect 48076 24782 48078 24834
rect 48130 24782 48132 24834
rect 46956 24722 47012 24734
rect 47852 24724 47908 24734
rect 46956 24670 46958 24722
rect 47010 24670 47012 24722
rect 45388 24612 45444 24622
rect 45388 24518 45444 24556
rect 44716 23998 44718 24050
rect 44770 23998 44772 24050
rect 44716 23986 44772 23998
rect 44268 23938 44324 23950
rect 44268 23886 44270 23938
rect 44322 23886 44324 23938
rect 44268 23156 44324 23886
rect 44268 23090 44324 23100
rect 44492 23938 44548 23950
rect 44492 23886 44494 23938
rect 44546 23886 44548 23938
rect 44492 23044 44548 23886
rect 46956 23828 47012 24670
rect 47740 24722 47908 24724
rect 47740 24670 47854 24722
rect 47906 24670 47908 24722
rect 47740 24668 47908 24670
rect 46172 23268 46228 23278
rect 46172 23174 46228 23212
rect 44716 23156 44772 23166
rect 44492 22594 44548 22988
rect 44492 22542 44494 22594
rect 44546 22542 44548 22594
rect 44492 22530 44548 22542
rect 44604 23154 44772 23156
rect 44604 23102 44718 23154
rect 44770 23102 44772 23154
rect 44604 23100 44772 23102
rect 43820 22482 43876 22494
rect 43820 22430 43822 22482
rect 43874 22430 43876 22482
rect 43820 22260 43876 22430
rect 43820 21588 43876 22204
rect 44268 22370 44324 22382
rect 44268 22318 44270 22370
rect 44322 22318 44324 22370
rect 44268 21700 44324 22318
rect 44492 21812 44548 21822
rect 44604 21812 44660 23100
rect 44716 23090 44772 23100
rect 45500 23156 45556 23166
rect 45500 22370 45556 23100
rect 45612 23044 45668 23054
rect 45612 22950 45668 22988
rect 46956 22930 47012 23772
rect 47516 23938 47572 23950
rect 47516 23886 47518 23938
rect 47570 23886 47572 23938
rect 47516 23828 47572 23886
rect 47516 23762 47572 23772
rect 47740 23938 47796 24668
rect 47852 24658 47908 24668
rect 47740 23886 47742 23938
rect 47794 23886 47796 23938
rect 47180 23268 47236 23278
rect 47180 23174 47236 23212
rect 47740 23268 47796 23886
rect 48076 23378 48132 24782
rect 48412 26068 48468 26078
rect 48412 24050 48468 26012
rect 49532 26068 49588 26106
rect 49532 26002 49588 26012
rect 49512 25900 49776 25910
rect 49568 25844 49616 25900
rect 49672 25844 49720 25900
rect 49512 25834 49776 25844
rect 49308 24948 49364 24958
rect 48412 23998 48414 24050
rect 48466 23998 48468 24050
rect 48412 23986 48468 23998
rect 48748 24164 48804 24174
rect 48076 23326 48078 23378
rect 48130 23326 48132 23378
rect 48076 23314 48132 23326
rect 46956 22878 46958 22930
rect 47010 22878 47012 22930
rect 45500 22318 45502 22370
rect 45554 22318 45556 22370
rect 45500 22306 45556 22318
rect 45724 22372 45780 22382
rect 45724 22278 45780 22316
rect 45948 22370 46004 22382
rect 45948 22318 45950 22370
rect 46002 22318 46004 22370
rect 44492 21810 44660 21812
rect 44492 21758 44494 21810
rect 44546 21758 44660 21810
rect 44492 21756 44660 21758
rect 44828 22260 44884 22270
rect 44828 21810 44884 22204
rect 44828 21758 44830 21810
rect 44882 21758 44884 21810
rect 44492 21746 44548 21756
rect 44828 21746 44884 21758
rect 45388 22148 45444 22158
rect 45388 21810 45444 22092
rect 45948 22148 46004 22318
rect 45948 22082 46004 22092
rect 45388 21758 45390 21810
rect 45442 21758 45444 21810
rect 45388 21746 45444 21758
rect 44268 21606 44324 21644
rect 44156 21588 44212 21598
rect 43820 21586 44212 21588
rect 43820 21534 44158 21586
rect 44210 21534 44212 21586
rect 43820 21532 44212 21534
rect 43372 19908 43428 19918
rect 43372 18676 43428 19852
rect 43596 19348 43652 19358
rect 43596 19254 43652 19292
rect 43820 19236 43876 21532
rect 44156 21522 44212 21532
rect 46508 21588 46564 21598
rect 45836 21476 45892 21486
rect 45836 21474 46004 21476
rect 45836 21422 45838 21474
rect 45890 21422 46004 21474
rect 45836 21420 46004 21422
rect 45836 21410 45892 21420
rect 45948 20916 46004 21420
rect 46060 20916 46116 20926
rect 45948 20914 46116 20916
rect 45948 20862 46062 20914
rect 46114 20862 46116 20914
rect 45948 20860 46116 20862
rect 45836 20804 45892 20814
rect 45388 20802 45892 20804
rect 45388 20750 45838 20802
rect 45890 20750 45892 20802
rect 45388 20748 45892 20750
rect 44604 20692 44660 20702
rect 44492 20636 44604 20692
rect 44380 20580 44436 20590
rect 44380 20486 44436 20524
rect 44492 20242 44548 20636
rect 44604 20598 44660 20636
rect 44716 20690 44772 20702
rect 44716 20638 44718 20690
rect 44770 20638 44772 20690
rect 44492 20190 44494 20242
rect 44546 20190 44548 20242
rect 44492 20178 44548 20190
rect 44716 20132 44772 20638
rect 45388 20580 45444 20748
rect 45836 20738 45892 20748
rect 45388 20242 45444 20524
rect 45388 20190 45390 20242
rect 45442 20190 45444 20242
rect 45388 20178 45444 20190
rect 44716 20066 44772 20076
rect 44156 20020 44212 20030
rect 44044 19964 44156 20020
rect 43932 19908 43988 19918
rect 43932 19814 43988 19852
rect 43932 19460 43988 19470
rect 44044 19460 44100 19964
rect 44156 19926 44212 19964
rect 44940 20018 44996 20030
rect 44940 19966 44942 20018
rect 44994 19966 44996 20018
rect 43932 19458 44100 19460
rect 43932 19406 43934 19458
rect 43986 19406 44100 19458
rect 43932 19404 44100 19406
rect 43932 19394 43988 19404
rect 43820 19180 43988 19236
rect 43372 18610 43428 18620
rect 43820 19010 43876 19022
rect 43820 18958 43822 19010
rect 43874 18958 43876 19010
rect 43596 18564 43652 18574
rect 43484 18340 43540 18350
rect 43484 18246 43540 18284
rect 43596 17892 43652 18508
rect 43708 18562 43764 18574
rect 43708 18510 43710 18562
rect 43762 18510 43764 18562
rect 43708 18452 43764 18510
rect 43708 18386 43764 18396
rect 43820 18338 43876 18958
rect 43820 18286 43822 18338
rect 43874 18286 43876 18338
rect 43820 18274 43876 18286
rect 43596 17826 43652 17836
rect 43820 16994 43876 17006
rect 43820 16942 43822 16994
rect 43874 16942 43876 16994
rect 43820 16884 43876 16942
rect 43820 16818 43876 16828
rect 43932 16436 43988 19180
rect 44492 19012 44548 19022
rect 44940 19012 44996 19966
rect 45612 20020 45668 20030
rect 46060 20020 46116 20860
rect 46508 20914 46564 21532
rect 46956 21588 47012 22878
rect 47292 22932 47348 22942
rect 47292 22838 47348 22876
rect 47404 22596 47460 22606
rect 47292 22148 47348 22158
rect 47292 22054 47348 22092
rect 46956 21522 47012 21532
rect 46508 20862 46510 20914
rect 46562 20862 46564 20914
rect 46508 20850 46564 20862
rect 46284 20130 46340 20142
rect 46284 20078 46286 20130
rect 46338 20078 46340 20130
rect 45612 20018 46116 20020
rect 45612 19966 45614 20018
rect 45666 19966 46116 20018
rect 45612 19964 46116 19966
rect 46172 20020 46228 20030
rect 45500 19908 45556 19918
rect 45500 19814 45556 19852
rect 44492 19010 44996 19012
rect 44492 18958 44494 19010
rect 44546 18958 44996 19010
rect 44492 18956 44996 18958
rect 45276 19572 45332 19582
rect 44492 18116 44548 18956
rect 44492 18050 44548 18060
rect 44940 18452 44996 18462
rect 44940 18338 44996 18396
rect 44940 18286 44942 18338
rect 44994 18286 44996 18338
rect 44716 17444 44772 17454
rect 44940 17444 44996 18286
rect 44716 17442 44996 17444
rect 44716 17390 44718 17442
rect 44770 17390 44996 17442
rect 44716 17388 44996 17390
rect 44044 16772 44100 16782
rect 44268 16772 44324 16782
rect 44044 16770 44212 16772
rect 44044 16718 44046 16770
rect 44098 16718 44212 16770
rect 44044 16716 44212 16718
rect 44044 16706 44100 16716
rect 43932 16370 43988 16380
rect 43372 15428 43428 15438
rect 43372 15334 43428 15372
rect 44044 15426 44100 15438
rect 44044 15374 44046 15426
rect 44098 15374 44100 15426
rect 43820 15314 43876 15326
rect 43820 15262 43822 15314
rect 43874 15262 43876 15314
rect 43260 15092 43652 15148
rect 43596 14868 43652 15092
rect 43596 14802 43652 14812
rect 43372 14644 43428 14654
rect 43148 13918 43150 13970
rect 43202 13918 43204 13970
rect 43148 13906 43204 13918
rect 43260 14084 43316 14094
rect 43260 13970 43316 14028
rect 43260 13918 43262 13970
rect 43314 13918 43316 13970
rect 43260 13906 43316 13918
rect 43372 13970 43428 14588
rect 43372 13918 43374 13970
rect 43426 13918 43428 13970
rect 43372 13906 43428 13918
rect 43820 13746 43876 15262
rect 44044 15316 44100 15374
rect 44044 15250 44100 15260
rect 44156 15428 44212 16716
rect 44156 14418 44212 15372
rect 44156 14366 44158 14418
rect 44210 14366 44212 14418
rect 44156 14354 44212 14366
rect 43820 13694 43822 13746
rect 43874 13694 43876 13746
rect 43820 13682 43876 13694
rect 42588 13134 42590 13186
rect 42642 13134 42644 13186
rect 42588 13122 42644 13134
rect 44268 13186 44324 16716
rect 44604 15316 44660 15326
rect 44604 15222 44660 15260
rect 44716 14980 44772 17388
rect 45276 17108 45332 19516
rect 45276 17042 45332 17052
rect 45388 19012 45444 19022
rect 45612 19012 45668 19964
rect 46172 19926 46228 19964
rect 46284 19796 46340 20078
rect 46508 20132 46564 20142
rect 46508 20038 46564 20076
rect 46284 19730 46340 19740
rect 46844 19906 46900 19918
rect 46844 19854 46846 19906
rect 46898 19854 46900 19906
rect 46844 19796 46900 19854
rect 46844 19730 46900 19740
rect 45388 19010 45668 19012
rect 45388 18958 45390 19010
rect 45442 18958 45668 19010
rect 45388 18956 45668 18958
rect 47068 19684 47124 19694
rect 45388 16772 45444 18956
rect 45836 18676 45892 18686
rect 45836 18582 45892 18620
rect 45612 18562 45668 18574
rect 45612 18510 45614 18562
rect 45666 18510 45668 18562
rect 45500 18452 45556 18462
rect 45500 18358 45556 18396
rect 45612 17780 45668 18510
rect 45836 18452 45892 18462
rect 45724 17780 45780 17790
rect 45612 17724 45724 17780
rect 45724 17666 45780 17724
rect 45836 17778 45892 18396
rect 45836 17726 45838 17778
rect 45890 17726 45892 17778
rect 45836 17714 45892 17726
rect 46956 18450 47012 18462
rect 46956 18398 46958 18450
rect 47010 18398 47012 18450
rect 45724 17614 45726 17666
rect 45778 17614 45780 17666
rect 45724 17602 45780 17614
rect 46620 17668 46676 17678
rect 46956 17668 47012 18398
rect 47068 18452 47124 19628
rect 47068 18386 47124 18396
rect 46620 17666 46956 17668
rect 46620 17614 46622 17666
rect 46674 17614 46956 17666
rect 46620 17612 46956 17614
rect 46620 17602 46676 17612
rect 46956 17536 47012 17612
rect 47180 18338 47236 18350
rect 47180 18286 47182 18338
rect 47234 18286 47236 18338
rect 47180 17444 47236 18286
rect 46172 17164 46676 17220
rect 46172 16994 46228 17164
rect 46172 16942 46174 16994
rect 46226 16942 46228 16994
rect 46172 16930 46228 16942
rect 46284 16994 46340 17006
rect 46284 16942 46286 16994
rect 46338 16942 46340 16994
rect 45388 16706 45444 16716
rect 45612 16770 45668 16782
rect 45612 16718 45614 16770
rect 45666 16718 45668 16770
rect 45612 16548 45668 16718
rect 45500 15540 45556 15550
rect 45612 15540 45668 16492
rect 46284 16548 46340 16942
rect 46284 16482 46340 16492
rect 46396 16996 46452 17006
rect 46284 16100 46340 16110
rect 45500 15538 45668 15540
rect 45500 15486 45502 15538
rect 45554 15486 45668 15538
rect 45500 15484 45668 15486
rect 45500 15474 45556 15484
rect 45612 15316 45668 15484
rect 46060 16098 46340 16100
rect 46060 16046 46286 16098
rect 46338 16046 46340 16098
rect 46060 16044 46340 16046
rect 45948 15316 46004 15326
rect 45612 15314 46004 15316
rect 45612 15262 45950 15314
rect 46002 15262 46004 15314
rect 45612 15260 46004 15262
rect 45948 15250 46004 15260
rect 44716 14914 44772 14924
rect 45948 14530 46004 14542
rect 45948 14478 45950 14530
rect 46002 14478 46004 14530
rect 44380 14418 44436 14430
rect 44380 14366 44382 14418
rect 44434 14366 44436 14418
rect 44380 13860 44436 14366
rect 45948 14196 46004 14478
rect 46060 14532 46116 16044
rect 46284 16034 46340 16044
rect 46396 16098 46452 16940
rect 46396 16046 46398 16098
rect 46450 16046 46452 16098
rect 46396 16034 46452 16046
rect 46508 16882 46564 16894
rect 46508 16830 46510 16882
rect 46562 16830 46564 16882
rect 46508 15988 46564 16830
rect 46620 16884 46676 17164
rect 46956 16884 47012 16894
rect 46620 16882 47012 16884
rect 46620 16830 46958 16882
rect 47010 16830 47012 16882
rect 46620 16828 47012 16830
rect 46620 15988 46676 15998
rect 46508 15986 46676 15988
rect 46508 15934 46622 15986
rect 46674 15934 46676 15986
rect 46508 15932 46676 15934
rect 46620 15922 46676 15932
rect 46172 15874 46228 15886
rect 46172 15822 46174 15874
rect 46226 15822 46228 15874
rect 46172 15538 46228 15822
rect 46172 15486 46174 15538
rect 46226 15486 46228 15538
rect 46172 15474 46228 15486
rect 46508 15764 46564 15774
rect 46396 15428 46452 15438
rect 46284 15426 46452 15428
rect 46284 15374 46398 15426
rect 46450 15374 46452 15426
rect 46284 15372 46452 15374
rect 46284 15314 46340 15372
rect 46396 15362 46452 15372
rect 46284 15262 46286 15314
rect 46338 15262 46340 15314
rect 46284 15250 46340 15262
rect 46060 14466 46116 14476
rect 46172 14642 46228 14654
rect 46172 14590 46174 14642
rect 46226 14590 46228 14642
rect 45948 14130 46004 14140
rect 45388 13860 45444 13870
rect 44380 13804 44660 13860
rect 44604 13748 44660 13804
rect 45388 13766 45444 13804
rect 46172 13860 46228 14590
rect 46284 14196 46340 14206
rect 46284 13970 46340 14140
rect 46284 13918 46286 13970
rect 46338 13918 46340 13970
rect 46284 13906 46340 13918
rect 46508 13970 46564 15708
rect 46732 15426 46788 16828
rect 46956 16818 47012 16828
rect 47068 16772 47124 16782
rect 47068 16678 47124 16716
rect 47180 16548 47236 17388
rect 46732 15374 46734 15426
rect 46786 15374 46788 15426
rect 46732 15362 46788 15374
rect 46956 16492 47236 16548
rect 47292 17442 47348 17454
rect 47292 17390 47294 17442
rect 47346 17390 47348 17442
rect 46844 15316 46900 15354
rect 46844 15250 46900 15260
rect 46956 15148 47012 16492
rect 47292 15764 47348 17390
rect 47404 16996 47460 22540
rect 47740 21812 47796 23212
rect 47852 23154 47908 23166
rect 47852 23102 47854 23154
rect 47906 23102 47908 23154
rect 47852 23044 47908 23102
rect 47852 22258 47908 22988
rect 48636 23044 48692 23054
rect 48636 22950 48692 22988
rect 48076 22932 48132 22942
rect 48076 22594 48132 22876
rect 48076 22542 48078 22594
rect 48130 22542 48132 22594
rect 48076 22530 48132 22542
rect 48188 22930 48244 22942
rect 48188 22878 48190 22930
rect 48242 22878 48244 22930
rect 48188 22482 48244 22878
rect 48188 22430 48190 22482
rect 48242 22430 48244 22482
rect 47852 22206 47854 22258
rect 47906 22206 47908 22258
rect 47852 22148 47908 22206
rect 47852 22082 47908 22092
rect 48076 22372 48132 22382
rect 47852 21812 47908 21822
rect 47740 21810 47908 21812
rect 47740 21758 47854 21810
rect 47906 21758 47908 21810
rect 47740 21756 47908 21758
rect 47852 21746 47908 21756
rect 48076 21810 48132 22316
rect 48188 22260 48244 22430
rect 48188 22194 48244 22204
rect 48076 21758 48078 21810
rect 48130 21758 48132 21810
rect 48076 21746 48132 21758
rect 48636 21698 48692 21710
rect 48636 21646 48638 21698
rect 48690 21646 48692 21698
rect 47740 21588 47796 21598
rect 47740 21494 47796 21532
rect 48300 21588 48356 21598
rect 48524 21588 48580 21598
rect 48300 20802 48356 21532
rect 48300 20750 48302 20802
rect 48354 20750 48356 20802
rect 48300 20692 48356 20750
rect 48300 20626 48356 20636
rect 48412 21586 48580 21588
rect 48412 21534 48526 21586
rect 48578 21534 48580 21586
rect 48412 21532 48580 21534
rect 48412 20804 48468 21532
rect 48524 21522 48580 21532
rect 47628 20244 47684 20254
rect 47628 18562 47684 20188
rect 48412 20244 48468 20748
rect 48636 20914 48692 21646
rect 48636 20862 48638 20914
rect 48690 20862 48692 20914
rect 48412 20130 48468 20188
rect 48412 20078 48414 20130
rect 48466 20078 48468 20130
rect 48412 20066 48468 20078
rect 48524 20356 48580 20366
rect 48524 20130 48580 20300
rect 48524 20078 48526 20130
rect 48578 20078 48580 20130
rect 48524 20066 48580 20078
rect 48636 20130 48692 20862
rect 48636 20078 48638 20130
rect 48690 20078 48692 20130
rect 48076 20020 48132 20030
rect 48076 19348 48132 19964
rect 48636 19908 48692 20078
rect 48636 19842 48692 19852
rect 47628 18510 47630 18562
rect 47682 18510 47684 18562
rect 47628 18498 47684 18510
rect 47740 19346 48132 19348
rect 47740 19294 48078 19346
rect 48130 19294 48132 19346
rect 47740 19292 48132 19294
rect 47628 17780 47684 17790
rect 47740 17780 47796 19292
rect 48076 19282 48132 19292
rect 48188 19234 48244 19246
rect 48188 19182 48190 19234
rect 48242 19182 48244 19234
rect 48188 18676 48244 19182
rect 48188 18610 48244 18620
rect 47628 17778 47796 17780
rect 47628 17726 47630 17778
rect 47682 17726 47796 17778
rect 47628 17724 47796 17726
rect 47852 18452 47908 18462
rect 47628 17714 47684 17724
rect 47516 17668 47572 17678
rect 47516 17574 47572 17612
rect 47740 17444 47796 17454
rect 47740 17350 47796 17388
rect 47628 17108 47684 17118
rect 47684 17052 47796 17108
rect 47628 17014 47684 17052
rect 47404 16930 47460 16940
rect 47628 16324 47684 16334
rect 47628 16098 47684 16268
rect 47628 16046 47630 16098
rect 47682 16046 47684 16098
rect 47628 16034 47684 16046
rect 47292 15698 47348 15708
rect 47740 15986 47796 17052
rect 47740 15934 47742 15986
rect 47794 15934 47796 15986
rect 47740 15652 47796 15934
rect 47404 15596 47796 15652
rect 47292 15540 47348 15550
rect 47404 15540 47460 15596
rect 47292 15538 47460 15540
rect 47292 15486 47294 15538
rect 47346 15486 47460 15538
rect 47292 15484 47460 15486
rect 47292 15474 47348 15484
rect 47852 15316 47908 18396
rect 48636 17108 48692 17118
rect 48636 17014 48692 17052
rect 48188 16996 48244 17006
rect 48188 16882 48244 16940
rect 48188 16830 48190 16882
rect 48242 16830 48244 16882
rect 48188 16818 48244 16830
rect 48748 16212 48804 24108
rect 49308 24052 49364 24892
rect 49512 24332 49776 24342
rect 49568 24276 49616 24332
rect 49672 24276 49720 24332
rect 49512 24266 49776 24276
rect 49308 23920 49364 23996
rect 49756 24164 49812 24174
rect 49756 24050 49812 24108
rect 50316 24164 50372 24174
rect 49756 23998 49758 24050
rect 49810 23998 49812 24050
rect 49756 23986 49812 23998
rect 49868 24052 49924 24062
rect 49868 23266 49924 23996
rect 49868 23214 49870 23266
rect 49922 23214 49924 23266
rect 49868 23202 49924 23214
rect 49980 23716 50036 23726
rect 49512 22764 49776 22774
rect 49568 22708 49616 22764
rect 49672 22708 49720 22764
rect 49512 22698 49776 22708
rect 49532 22596 49588 22606
rect 49532 22502 49588 22540
rect 49420 22372 49476 22382
rect 49980 22372 50036 23660
rect 50092 23492 50148 23502
rect 50092 23378 50148 23436
rect 50092 23326 50094 23378
rect 50146 23326 50148 23378
rect 50092 23314 50148 23326
rect 50316 23378 50372 24108
rect 50988 23714 51044 23726
rect 50988 23662 50990 23714
rect 51042 23662 51044 23714
rect 50988 23492 51044 23662
rect 50988 23426 51044 23436
rect 50316 23326 50318 23378
rect 50370 23326 50372 23378
rect 50316 23314 50372 23326
rect 50540 23156 50596 23166
rect 50988 23156 51044 23166
rect 50540 23154 51044 23156
rect 50540 23102 50542 23154
rect 50594 23102 50990 23154
rect 51042 23102 51044 23154
rect 50540 23100 51044 23102
rect 50540 23090 50596 23100
rect 49420 22278 49476 22316
rect 49756 22316 50036 22372
rect 50204 23042 50260 23054
rect 50204 22990 50206 23042
rect 50258 22990 50260 23042
rect 48860 21588 48916 21598
rect 49420 21588 49476 21598
rect 48860 21586 49476 21588
rect 48860 21534 48862 21586
rect 48914 21534 49422 21586
rect 49474 21534 49476 21586
rect 48860 21532 49476 21534
rect 48860 21522 48916 21532
rect 49420 21522 49476 21532
rect 49756 21364 49812 22316
rect 49980 22148 50036 22158
rect 49980 21810 50036 22092
rect 50204 21924 50260 22990
rect 50988 22708 51044 23100
rect 50988 22642 51044 22652
rect 50204 21858 50260 21868
rect 49980 21758 49982 21810
rect 50034 21758 50036 21810
rect 49980 21746 50036 21758
rect 50316 21700 50372 21710
rect 49868 21588 49924 21598
rect 49868 21494 49924 21532
rect 50092 21586 50148 21598
rect 50092 21534 50094 21586
rect 50146 21534 50148 21586
rect 49756 21308 49924 21364
rect 49512 21196 49776 21206
rect 49568 21140 49616 21196
rect 49672 21140 49720 21196
rect 49512 21130 49776 21140
rect 49868 21026 49924 21308
rect 49868 20974 49870 21026
rect 49922 20974 49924 21026
rect 49868 20962 49924 20974
rect 49644 20804 49700 20814
rect 49644 20710 49700 20748
rect 50092 20356 50148 21534
rect 50092 20290 50148 20300
rect 49532 20020 49588 20058
rect 49532 19954 49588 19964
rect 49532 19796 49588 19806
rect 49308 19794 49588 19796
rect 49308 19742 49534 19794
rect 49586 19742 49588 19794
rect 49308 19740 49588 19742
rect 49308 19012 49364 19740
rect 49532 19730 49588 19740
rect 49868 19794 49924 19806
rect 49868 19742 49870 19794
rect 49922 19742 49924 19794
rect 49512 19628 49776 19638
rect 49568 19572 49616 19628
rect 49672 19572 49720 19628
rect 49512 19562 49776 19572
rect 49644 19460 49700 19470
rect 49308 18956 49588 19012
rect 49308 18788 49364 18798
rect 48972 17442 49028 17454
rect 48972 17390 48974 17442
rect 49026 17390 49028 17442
rect 48972 16772 49028 17390
rect 48972 16706 49028 16716
rect 48860 16212 48916 16222
rect 48748 16210 48916 16212
rect 48748 16158 48862 16210
rect 48914 16158 48916 16210
rect 48748 16156 48916 16158
rect 48860 16146 48916 16156
rect 48524 16100 48580 16110
rect 48300 16044 48524 16100
rect 47964 15876 48020 15886
rect 47964 15874 48132 15876
rect 47964 15822 47966 15874
rect 48018 15822 48132 15874
rect 47964 15820 48132 15822
rect 47964 15810 48020 15820
rect 47964 15316 48020 15326
rect 47852 15314 48020 15316
rect 47852 15262 47966 15314
rect 48018 15262 48020 15314
rect 47852 15260 48020 15262
rect 47964 15250 48020 15260
rect 46732 15092 47012 15148
rect 46732 14754 46788 15092
rect 46732 14702 46734 14754
rect 46786 14702 46788 14754
rect 46732 14690 46788 14702
rect 48076 14644 48132 15820
rect 48076 14578 48132 14588
rect 46508 13918 46510 13970
rect 46562 13918 46564 13970
rect 46508 13906 46564 13918
rect 44940 13748 44996 13758
rect 44604 13746 44996 13748
rect 44604 13694 44942 13746
rect 44994 13694 44996 13746
rect 46172 13728 46228 13804
rect 44604 13692 44996 13694
rect 44268 13134 44270 13186
rect 44322 13134 44324 13186
rect 44268 13122 44324 13134
rect 44492 13634 44548 13646
rect 44492 13582 44494 13634
rect 44546 13582 44548 13634
rect 42028 13010 42084 13020
rect 43596 13074 43652 13086
rect 43596 13022 43598 13074
rect 43650 13022 43652 13074
rect 40796 12964 40852 12974
rect 40796 12870 40852 12908
rect 42476 12964 42532 12974
rect 43484 12964 43540 12974
rect 42476 12870 42532 12908
rect 42924 12962 43540 12964
rect 42924 12910 43486 12962
rect 43538 12910 43540 12962
rect 42924 12908 43540 12910
rect 40460 12226 40516 12236
rect 41916 12740 41972 12750
rect 42588 12740 42644 12750
rect 41916 12738 42644 12740
rect 41916 12686 41918 12738
rect 41970 12686 42590 12738
rect 42642 12686 42644 12738
rect 41916 12684 42644 12686
rect 41916 11508 41972 12684
rect 42588 12404 42644 12684
rect 42924 12404 42980 12908
rect 43484 12898 43540 12908
rect 43596 12964 43652 13022
rect 43596 12898 43652 12908
rect 44492 12852 44548 13582
rect 44940 12964 44996 13692
rect 45948 13636 46004 13646
rect 45948 13074 46004 13580
rect 45948 13022 45950 13074
rect 46002 13022 46004 13074
rect 45948 13010 46004 13022
rect 46844 13412 46900 13422
rect 44940 12898 44996 12908
rect 45836 12964 45892 12974
rect 45836 12870 45892 12908
rect 42588 12402 42980 12404
rect 42588 12350 42926 12402
rect 42978 12350 42980 12402
rect 42588 12348 42980 12350
rect 42924 12338 42980 12348
rect 44268 12740 44324 12750
rect 43820 12180 43876 12190
rect 43596 12178 43876 12180
rect 43596 12126 43822 12178
rect 43874 12126 43876 12178
rect 43596 12124 43876 12126
rect 42588 12068 42644 12078
rect 42588 11974 42644 12012
rect 43596 12068 43652 12124
rect 43820 12114 43876 12124
rect 43932 12180 43988 12190
rect 41916 11442 41972 11452
rect 43596 11506 43652 12012
rect 43932 11620 43988 12124
rect 43932 11554 43988 11564
rect 44156 12066 44212 12078
rect 44156 12014 44158 12066
rect 44210 12014 44212 12066
rect 43596 11454 43598 11506
rect 43650 11454 43652 11506
rect 40572 11282 40628 11294
rect 40572 11230 40574 11282
rect 40626 11230 40628 11282
rect 40460 11170 40516 11182
rect 40460 11118 40462 11170
rect 40514 11118 40516 11170
rect 40460 10164 40516 11118
rect 40572 11172 40628 11230
rect 41020 11172 41076 11182
rect 40572 11170 41076 11172
rect 40572 11118 41022 11170
rect 41074 11118 41076 11170
rect 40572 11116 41076 11118
rect 40572 10612 40628 11116
rect 41020 11106 41076 11116
rect 43596 11172 43652 11454
rect 43596 11106 43652 11116
rect 44156 11394 44212 12014
rect 44268 11618 44324 12684
rect 44492 11954 44548 12796
rect 46060 12852 46116 12862
rect 46060 12758 46116 12796
rect 45612 12740 45668 12750
rect 45612 12646 45668 12684
rect 44492 11902 44494 11954
rect 44546 11902 44548 11954
rect 44492 11890 44548 11902
rect 45388 12292 45444 12302
rect 44268 11566 44270 11618
rect 44322 11566 44324 11618
rect 44268 11554 44324 11566
rect 44156 11342 44158 11394
rect 44210 11342 44212 11394
rect 42252 10724 42308 10734
rect 44156 10724 44212 11342
rect 44268 11172 44324 11182
rect 44268 11078 44324 11116
rect 45388 10834 45444 12236
rect 45388 10782 45390 10834
rect 45442 10782 45444 10834
rect 45388 10770 45444 10782
rect 44380 10724 44436 10734
rect 44156 10722 44436 10724
rect 44156 10670 44382 10722
rect 44434 10670 44436 10722
rect 44156 10668 44436 10670
rect 40572 10546 40628 10556
rect 40796 10612 40852 10622
rect 40796 10518 40852 10556
rect 41468 10500 41524 10510
rect 41468 10406 41524 10444
rect 40460 10098 40516 10108
rect 40572 9828 40628 9838
rect 40572 9604 40628 9772
rect 40348 9538 40404 9548
rect 40460 9602 40628 9604
rect 40460 9550 40574 9602
rect 40626 9550 40628 9602
rect 40460 9548 40628 9550
rect 40460 8820 40516 9548
rect 40572 9538 40628 9548
rect 41132 9826 41188 9838
rect 41132 9774 41134 9826
rect 41186 9774 41188 9826
rect 40684 9268 40740 9278
rect 40684 9174 40740 9212
rect 40460 8428 40516 8764
rect 40572 9156 40628 9166
rect 40572 8596 40628 9100
rect 40908 9044 40964 9054
rect 40908 8950 40964 8988
rect 40572 8530 40628 8540
rect 41132 8428 41188 9774
rect 41356 9828 41412 9838
rect 41356 9734 41412 9772
rect 41692 9602 41748 9614
rect 41692 9550 41694 9602
rect 41746 9550 41748 9602
rect 41580 9044 41636 9054
rect 40460 8372 40740 8428
rect 40684 8034 40740 8372
rect 40796 8372 41188 8428
rect 41468 8988 41580 9044
rect 41692 9044 41748 9550
rect 42140 9604 42196 9614
rect 42140 9510 42196 9548
rect 42140 9268 42196 9278
rect 42252 9268 42308 10668
rect 44380 10658 44436 10668
rect 42812 10612 42868 10622
rect 43820 10612 43876 10622
rect 44828 10612 44884 10622
rect 42812 10610 43204 10612
rect 42812 10558 42814 10610
rect 42866 10558 43204 10610
rect 42812 10556 43204 10558
rect 42812 10546 42868 10556
rect 42476 10388 42532 10398
rect 42476 10294 42532 10332
rect 42812 10388 42868 10398
rect 42812 10294 42868 10332
rect 43148 10050 43204 10556
rect 43820 10518 43876 10556
rect 44604 10610 44884 10612
rect 44604 10558 44830 10610
rect 44882 10558 44884 10610
rect 44604 10556 44884 10558
rect 44044 10500 44100 10510
rect 44044 10406 44100 10444
rect 43148 9998 43150 10050
rect 43202 9998 43204 10050
rect 43148 9986 43204 9998
rect 44604 10050 44660 10556
rect 44828 10546 44884 10556
rect 45276 10612 45332 10622
rect 45276 10518 45332 10556
rect 45500 10610 45556 10622
rect 45500 10558 45502 10610
rect 45554 10558 45556 10610
rect 44604 9998 44606 10050
rect 44658 9998 44660 10050
rect 44604 9986 44660 9998
rect 45500 10500 45556 10558
rect 44716 9828 44772 9838
rect 44716 9734 44772 9772
rect 45500 9826 45556 10444
rect 45500 9774 45502 9826
rect 45554 9774 45556 9826
rect 45500 9762 45556 9774
rect 45724 9828 45780 9838
rect 43484 9714 43540 9726
rect 43484 9662 43486 9714
rect 43538 9662 43540 9714
rect 42140 9266 42308 9268
rect 42140 9214 42142 9266
rect 42194 9214 42308 9266
rect 42140 9212 42308 9214
rect 42364 9604 42420 9614
rect 42140 9202 42196 9212
rect 42364 9156 42420 9548
rect 41804 9044 41860 9054
rect 41692 9042 41860 9044
rect 41692 8990 41806 9042
rect 41858 8990 41860 9042
rect 41692 8988 41860 8990
rect 40796 8306 40852 8316
rect 41468 8370 41524 8988
rect 41580 8950 41636 8988
rect 41804 8978 41860 8988
rect 42028 9042 42084 9054
rect 42028 8990 42030 9042
rect 42082 8990 42084 9042
rect 41692 8820 41748 8830
rect 41692 8596 41748 8764
rect 41468 8318 41470 8370
rect 41522 8318 41524 8370
rect 41468 8306 41524 8318
rect 41580 8372 41636 8382
rect 41580 8146 41636 8316
rect 41580 8094 41582 8146
rect 41634 8094 41636 8146
rect 41580 8082 41636 8094
rect 40684 7982 40686 8034
rect 40738 7982 40740 8034
rect 40684 7924 40740 7982
rect 40684 7858 40740 7868
rect 40012 7698 40292 7700
rect 40012 7646 40014 7698
rect 40066 7646 40292 7698
rect 40012 7644 40292 7646
rect 40012 7634 40068 7644
rect 39564 7074 39620 7084
rect 39900 7474 39956 7486
rect 39900 7422 39902 7474
rect 39954 7422 39956 7474
rect 39900 6916 39956 7422
rect 39116 5954 39172 5964
rect 39340 5908 39396 6524
rect 39340 5842 39396 5852
rect 39452 6914 39956 6916
rect 39452 6862 39902 6914
rect 39954 6862 39956 6914
rect 39452 6860 39956 6862
rect 39452 5794 39508 6860
rect 39900 6850 39956 6860
rect 40124 7474 40180 7486
rect 40124 7422 40126 7474
rect 40178 7422 40180 7474
rect 39676 6692 39732 6702
rect 39676 6598 39732 6636
rect 40124 6580 40180 7422
rect 40572 7476 40628 7486
rect 40572 7474 41076 7476
rect 40572 7422 40574 7474
rect 40626 7422 41076 7474
rect 40572 7420 41076 7422
rect 40572 7410 40628 7420
rect 40124 6514 40180 6524
rect 40348 6690 40404 6702
rect 40348 6638 40350 6690
rect 40402 6638 40404 6690
rect 40348 6468 40404 6638
rect 41020 6690 41076 7420
rect 41020 6638 41022 6690
rect 41074 6638 41076 6690
rect 41020 6626 41076 6638
rect 41356 6692 41412 6702
rect 41356 6598 41412 6636
rect 39676 6356 39732 6366
rect 39564 5908 39620 5918
rect 39564 5814 39620 5852
rect 39452 5742 39454 5794
rect 39506 5742 39508 5794
rect 39452 5730 39508 5742
rect 39676 5348 39732 6300
rect 39852 6300 40116 6310
rect 39908 6244 39956 6300
rect 40012 6244 40060 6300
rect 39852 6234 40116 6244
rect 39788 5348 39844 5358
rect 39676 5346 39844 5348
rect 39676 5294 39790 5346
rect 39842 5294 39844 5346
rect 39676 5292 39844 5294
rect 39116 5236 39172 5246
rect 39116 5142 39172 5180
rect 38108 4562 38276 4564
rect 38108 4510 38110 4562
rect 38162 4510 38276 4562
rect 38108 4508 38276 4510
rect 38108 4498 38164 4508
rect 37772 4338 38052 4340
rect 37772 4286 37774 4338
rect 37826 4286 38052 4338
rect 37772 4284 38052 4286
rect 37772 4274 37828 4284
rect 38668 4228 38724 4238
rect 38892 4228 38948 5068
rect 39004 5012 39060 5022
rect 39004 4918 39060 4956
rect 39228 4898 39284 4910
rect 39228 4846 39230 4898
rect 39282 4846 39284 4898
rect 38668 4134 38724 4172
rect 38780 4226 38948 4228
rect 38780 4174 38894 4226
rect 38946 4174 38948 4226
rect 38780 4172 38948 4174
rect 38668 3668 38724 3678
rect 38780 3668 38836 4172
rect 38892 4162 38948 4172
rect 39116 4564 39172 4574
rect 38668 3666 38836 3668
rect 38668 3614 38670 3666
rect 38722 3614 38836 3666
rect 38668 3612 38836 3614
rect 38668 3602 38724 3612
rect 38220 3556 38276 3566
rect 39116 3556 39172 4508
rect 39228 4228 39284 4846
rect 39452 4900 39508 4910
rect 39452 4338 39508 4844
rect 39452 4286 39454 4338
rect 39506 4286 39508 4338
rect 39452 4274 39508 4286
rect 39228 4162 39284 4172
rect 38220 3462 38276 3500
rect 38892 3554 39172 3556
rect 38892 3502 39118 3554
rect 39170 3502 39172 3554
rect 38892 3500 39172 3502
rect 39676 3556 39732 5292
rect 39788 5124 39844 5292
rect 40348 5236 40404 6412
rect 41244 6468 41300 6478
rect 41244 6374 41300 6412
rect 40796 5908 40852 5918
rect 40796 5814 40852 5852
rect 41692 5794 41748 8540
rect 42028 7700 42084 8990
rect 42252 9044 42308 9054
rect 42364 9044 42420 9100
rect 42252 9042 42420 9044
rect 42252 8990 42254 9042
rect 42306 8990 42420 9042
rect 42252 8988 42420 8990
rect 42700 9604 42756 9614
rect 42252 8932 42308 8988
rect 42252 8866 42308 8876
rect 42700 8708 42756 9548
rect 43260 9604 43316 9614
rect 43260 9510 43316 9548
rect 43484 9492 43540 9662
rect 44604 9716 44660 9726
rect 43484 9426 43540 9436
rect 43932 9602 43988 9614
rect 43932 9550 43934 9602
rect 43986 9550 43988 9602
rect 43932 9492 43988 9550
rect 43932 9426 43988 9436
rect 42700 8642 42756 8652
rect 42924 9380 42980 9390
rect 42924 9042 42980 9324
rect 43036 9268 43092 9278
rect 43596 9268 43652 9278
rect 43092 9266 43652 9268
rect 43092 9214 43598 9266
rect 43650 9214 43652 9266
rect 43092 9212 43652 9214
rect 43036 9136 43092 9212
rect 43596 9202 43652 9212
rect 44044 9268 44100 9278
rect 44044 9174 44100 9212
rect 42924 8990 42926 9042
rect 42978 8990 42980 9042
rect 42924 8484 42980 8990
rect 43260 9042 43316 9054
rect 43260 8990 43262 9042
rect 43314 8990 43316 9042
rect 43260 8708 43316 8990
rect 43260 8642 43316 8652
rect 44604 8428 44660 9660
rect 45388 9604 45444 9614
rect 45276 9268 45332 9278
rect 45276 8820 45332 9212
rect 45276 8754 45332 8764
rect 42924 8418 42980 8428
rect 44380 8372 44660 8428
rect 43484 8260 43540 8270
rect 43484 8166 43540 8204
rect 43260 8146 43316 8158
rect 43260 8094 43262 8146
rect 43314 8094 43316 8146
rect 43260 7924 43316 8094
rect 43260 7858 43316 7868
rect 42028 7634 42084 7644
rect 44380 7698 44436 8372
rect 45388 8148 45444 9548
rect 45724 8372 45780 9772
rect 45948 9826 46004 9838
rect 45948 9774 45950 9826
rect 46002 9774 46004 9826
rect 45948 9716 46004 9774
rect 45948 9650 46004 9660
rect 45836 8372 45892 8382
rect 45724 8370 45892 8372
rect 45724 8318 45838 8370
rect 45890 8318 45892 8370
rect 45724 8316 45892 8318
rect 45836 8306 45892 8316
rect 46284 8260 46340 8270
rect 46732 8260 46788 8270
rect 46284 8166 46340 8204
rect 46620 8204 46732 8260
rect 45388 8082 45444 8092
rect 44380 7646 44382 7698
rect 44434 7646 44436 7698
rect 44380 7634 44436 7646
rect 42924 7476 42980 7486
rect 42812 7252 42868 7262
rect 42588 6692 42644 6702
rect 42588 6598 42644 6636
rect 42140 6468 42196 6478
rect 41692 5742 41694 5794
rect 41746 5742 41748 5794
rect 41692 5730 41748 5742
rect 42028 6466 42196 6468
rect 42028 6414 42142 6466
rect 42194 6414 42196 6466
rect 42028 6412 42196 6414
rect 40348 5170 40404 5180
rect 40460 5348 40516 5358
rect 39788 5058 39844 5068
rect 40124 5122 40180 5134
rect 40124 5070 40126 5122
rect 40178 5070 40180 5122
rect 40124 5012 40180 5070
rect 40124 4946 40180 4956
rect 40460 5010 40516 5292
rect 41020 5124 41076 5134
rect 41020 5030 41076 5068
rect 41468 5122 41524 5134
rect 41468 5070 41470 5122
rect 41522 5070 41524 5122
rect 40460 4958 40462 5010
rect 40514 4958 40516 5010
rect 40460 4946 40516 4958
rect 40236 4898 40292 4910
rect 40236 4846 40238 4898
rect 40290 4846 40292 4898
rect 40236 4788 40292 4846
rect 40348 4900 40404 4910
rect 40348 4806 40404 4844
rect 39852 4732 40116 4742
rect 39908 4676 39956 4732
rect 40012 4676 40060 4732
rect 39852 4666 40116 4676
rect 40236 4228 40292 4732
rect 41468 4788 41524 5070
rect 41468 4722 41524 4732
rect 41804 5012 41860 5022
rect 41356 4676 41412 4686
rect 40460 4564 40516 4574
rect 40348 4452 40404 4462
rect 40348 4358 40404 4396
rect 40460 4450 40516 4508
rect 40460 4398 40462 4450
rect 40514 4398 40516 4450
rect 40460 4386 40516 4398
rect 41356 4340 41412 4620
rect 41356 4274 41412 4284
rect 41580 4676 41636 4686
rect 40236 4172 40404 4228
rect 40348 4114 40404 4172
rect 40348 4062 40350 4114
rect 40402 4062 40404 4114
rect 40236 4004 40292 4014
rect 39900 3556 39956 3566
rect 39676 3554 39956 3556
rect 39676 3502 39902 3554
rect 39954 3502 39956 3554
rect 39676 3500 39956 3502
rect 37660 1586 37716 1596
rect 37548 802 37604 812
rect 38892 800 38948 3500
rect 39116 3490 39172 3500
rect 39900 3490 39956 3500
rect 40124 3556 40180 3566
rect 39452 3444 39508 3454
rect 39452 3350 39508 3388
rect 40124 3330 40180 3500
rect 40236 3554 40292 3948
rect 40236 3502 40238 3554
rect 40290 3502 40292 3554
rect 40236 3444 40292 3502
rect 40236 3378 40292 3388
rect 40124 3278 40126 3330
rect 40178 3278 40180 3330
rect 40124 3266 40180 3278
rect 40348 3220 40404 4062
rect 41580 3668 41636 4620
rect 41692 4564 41748 4574
rect 41804 4564 41860 4956
rect 41916 4900 41972 4910
rect 41916 4806 41972 4844
rect 42028 4676 42084 6412
rect 42140 6402 42196 6412
rect 42140 5908 42196 5918
rect 42588 5908 42644 5918
rect 42140 5814 42196 5852
rect 42252 5906 42644 5908
rect 42252 5854 42590 5906
rect 42642 5854 42644 5906
rect 42252 5852 42644 5854
rect 42028 4610 42084 4620
rect 42140 5460 42196 5470
rect 41916 4564 41972 4574
rect 41804 4562 41972 4564
rect 41804 4510 41918 4562
rect 41970 4510 41972 4562
rect 41804 4508 41972 4510
rect 41692 4470 41748 4508
rect 41916 4498 41972 4508
rect 42028 4452 42084 4462
rect 42140 4452 42196 5404
rect 42028 4450 42196 4452
rect 42028 4398 42030 4450
rect 42082 4398 42196 4450
rect 42028 4396 42196 4398
rect 42252 4900 42308 5852
rect 42588 5842 42644 5852
rect 42476 5684 42532 5694
rect 42476 5236 42532 5628
rect 42476 5234 42756 5236
rect 42476 5182 42478 5234
rect 42530 5182 42756 5234
rect 42476 5180 42756 5182
rect 42476 5170 42532 5180
rect 42252 4452 42308 4844
rect 42028 4386 42084 4396
rect 42252 4358 42308 4396
rect 42364 4788 42420 4798
rect 41804 4340 41860 4350
rect 41804 4246 41860 4284
rect 42364 4340 42420 4732
rect 42700 4564 42756 5180
rect 42812 4676 42868 7196
rect 42924 6468 42980 7420
rect 43932 7476 43988 7486
rect 44268 7476 44324 7486
rect 43036 7364 43092 7374
rect 43036 6690 43092 7308
rect 43484 6804 43540 6814
rect 43484 6710 43540 6748
rect 43036 6638 43038 6690
rect 43090 6638 43092 6690
rect 43036 6626 43092 6638
rect 42924 6412 43092 6468
rect 42924 6244 42980 6254
rect 42924 5460 42980 6188
rect 42924 5234 42980 5404
rect 42924 5182 42926 5234
rect 42978 5182 42980 5234
rect 42924 5170 42980 5182
rect 42812 4620 42980 4676
rect 42700 4432 42756 4508
rect 42364 4274 42420 4284
rect 42924 3780 42980 4620
rect 42924 3686 42980 3724
rect 41244 3444 41300 3454
rect 39852 3164 40116 3174
rect 39908 3108 39956 3164
rect 40012 3108 40060 3164
rect 39852 3098 40116 3108
rect 40236 3164 40404 3220
rect 41020 3388 41244 3444
rect 40236 2100 40292 3164
rect 40236 2034 40292 2044
rect 41020 800 41076 3388
rect 41244 3312 41300 3388
rect 41580 3330 41636 3612
rect 42812 3668 42868 3678
rect 42812 3554 42868 3612
rect 42812 3502 42814 3554
rect 42866 3502 42868 3554
rect 42812 3490 42868 3502
rect 42028 3444 42084 3454
rect 42028 3350 42084 3388
rect 41580 3278 41582 3330
rect 41634 3278 41636 3330
rect 41580 3266 41636 3278
rect 42924 3330 42980 3342
rect 42924 3278 42926 3330
rect 42978 3278 42980 3330
rect 42924 3220 42980 3278
rect 42924 3154 42980 3164
rect 43036 980 43092 6412
rect 43036 914 43092 924
rect 43148 5794 43204 5806
rect 43148 5742 43150 5794
rect 43202 5742 43204 5794
rect 43148 4452 43204 5742
rect 43484 5796 43540 5806
rect 43484 5794 43652 5796
rect 43484 5742 43486 5794
rect 43538 5742 43652 5794
rect 43484 5740 43652 5742
rect 43484 5730 43540 5740
rect 43372 5122 43428 5134
rect 43372 5070 43374 5122
rect 43426 5070 43428 5122
rect 43372 4788 43428 5070
rect 43372 4722 43428 4732
rect 43596 4900 43652 5740
rect 43484 4452 43540 4462
rect 43148 4450 43540 4452
rect 43148 4398 43486 4450
rect 43538 4398 43540 4450
rect 43148 4396 43540 4398
rect 43148 800 43204 4396
rect 43484 4386 43540 4396
rect 43596 3554 43652 4844
rect 43596 3502 43598 3554
rect 43650 3502 43652 3554
rect 43596 2884 43652 3502
rect 43596 2818 43652 2828
rect 43708 4788 43764 4798
rect 43708 1540 43764 4732
rect 43708 1474 43764 1484
rect 43932 1540 43988 7420
rect 44156 7474 44324 7476
rect 44156 7422 44270 7474
rect 44322 7422 44324 7474
rect 44156 7420 44324 7422
rect 44156 6804 44212 7420
rect 44268 7410 44324 7420
rect 44492 7474 44548 7486
rect 44492 7422 44494 7474
rect 44546 7422 44548 7474
rect 44492 7364 44548 7422
rect 44940 7476 44996 7486
rect 44940 7474 45332 7476
rect 44940 7422 44942 7474
rect 44994 7422 45332 7474
rect 44940 7420 45332 7422
rect 44940 7410 44996 7420
rect 44492 7298 44548 7308
rect 44156 5794 44212 6748
rect 44156 5742 44158 5794
rect 44210 5742 44212 5794
rect 44156 5730 44212 5742
rect 44380 6466 44436 6478
rect 44716 6468 44772 6478
rect 44380 6414 44382 6466
rect 44434 6414 44436 6466
rect 44380 5124 44436 6414
rect 44604 6466 44772 6468
rect 44604 6414 44718 6466
rect 44770 6414 44772 6466
rect 44604 6412 44772 6414
rect 44604 6356 44660 6412
rect 44716 6402 44772 6412
rect 44044 5068 44436 5124
rect 44492 5124 44548 5134
rect 44604 5124 44660 6300
rect 44940 5906 44996 5918
rect 44940 5854 44942 5906
rect 44994 5854 44996 5906
rect 44828 5794 44884 5806
rect 44828 5742 44830 5794
rect 44882 5742 44884 5794
rect 44828 5236 44884 5742
rect 44828 5170 44884 5180
rect 44492 5122 44660 5124
rect 44492 5070 44494 5122
rect 44546 5070 44660 5122
rect 44492 5068 44660 5070
rect 44044 4340 44100 5068
rect 44492 5058 44548 5068
rect 44716 5010 44772 5022
rect 44716 4958 44718 5010
rect 44770 4958 44772 5010
rect 44156 4898 44212 4910
rect 44156 4846 44158 4898
rect 44210 4846 44212 4898
rect 44156 4788 44212 4846
rect 44268 4900 44324 4910
rect 44268 4806 44324 4844
rect 44380 4898 44436 4910
rect 44380 4846 44382 4898
rect 44434 4846 44436 4898
rect 44156 4564 44212 4732
rect 44156 4498 44212 4508
rect 44380 4340 44436 4846
rect 44716 4788 44772 4958
rect 44940 5012 44996 5854
rect 45276 5124 45332 7420
rect 45388 7362 45444 7374
rect 45388 7310 45390 7362
rect 45442 7310 45444 7362
rect 45388 7252 45444 7310
rect 46620 7362 46676 8204
rect 46732 8166 46788 8204
rect 46620 7310 46622 7362
rect 46674 7310 46676 7362
rect 46620 7298 46676 7310
rect 46844 7812 46900 13356
rect 48300 13412 48356 16044
rect 48524 16006 48580 16044
rect 48412 15316 48468 15326
rect 48412 15222 48468 15260
rect 49308 14756 49364 18732
rect 49532 18674 49588 18956
rect 49532 18622 49534 18674
rect 49586 18622 49588 18674
rect 49532 18610 49588 18622
rect 49644 18674 49700 19404
rect 49868 19348 49924 19742
rect 49868 19234 49924 19292
rect 50316 19346 50372 21644
rect 50316 19294 50318 19346
rect 50370 19294 50372 19346
rect 50316 19282 50372 19294
rect 50988 20020 51044 20030
rect 49868 19182 49870 19234
rect 49922 19182 49924 19234
rect 49868 18788 49924 19182
rect 50988 19122 51044 19964
rect 51100 19348 51156 19358
rect 51100 19234 51156 19292
rect 51100 19182 51102 19234
rect 51154 19182 51156 19234
rect 51100 19170 51156 19182
rect 50988 19070 50990 19122
rect 51042 19070 51044 19122
rect 50988 19058 51044 19070
rect 49868 18722 49924 18732
rect 50204 19012 50260 19022
rect 49644 18622 49646 18674
rect 49698 18622 49700 18674
rect 49644 18610 49700 18622
rect 49756 18676 49812 18686
rect 49756 18582 49812 18620
rect 50204 18450 50260 18956
rect 50764 19012 50820 19022
rect 50764 18918 50820 18956
rect 50204 18398 50206 18450
rect 50258 18398 50260 18450
rect 50204 18386 50260 18398
rect 50316 18900 50372 18910
rect 49512 18060 49776 18070
rect 49568 18004 49616 18060
rect 49672 18004 49720 18060
rect 49512 17994 49776 18004
rect 49980 17892 50036 17902
rect 49420 17442 49476 17454
rect 49420 17390 49422 17442
rect 49474 17390 49476 17442
rect 49420 16996 49476 17390
rect 49420 16884 49476 16940
rect 49980 16996 50036 17836
rect 50316 17668 50372 18844
rect 50876 18788 50932 18798
rect 50652 18452 50708 18462
rect 50652 18358 50708 18396
rect 50316 17442 50372 17612
rect 50764 17556 50820 17566
rect 50764 17462 50820 17500
rect 50316 17390 50318 17442
rect 50370 17390 50372 17442
rect 49980 16994 50148 16996
rect 49980 16942 49982 16994
rect 50034 16942 50148 16994
rect 49980 16940 50148 16942
rect 49980 16930 50036 16940
rect 49532 16884 49588 16894
rect 49420 16882 49588 16884
rect 49420 16830 49534 16882
rect 49586 16830 49588 16882
rect 49420 16828 49588 16830
rect 49532 16818 49588 16828
rect 49756 16882 49812 16894
rect 49756 16830 49758 16882
rect 49810 16830 49812 16882
rect 49756 16772 49812 16830
rect 49756 16660 49812 16716
rect 50092 16772 50148 16940
rect 50316 16884 50372 17390
rect 50540 17444 50596 17454
rect 50540 17106 50596 17388
rect 50540 17054 50542 17106
rect 50594 17054 50596 17106
rect 50540 17042 50596 17054
rect 50316 16882 50596 16884
rect 50316 16830 50318 16882
rect 50370 16830 50596 16882
rect 50316 16828 50596 16830
rect 50316 16818 50372 16828
rect 50092 16706 50148 16716
rect 49756 16604 50036 16660
rect 49512 16492 49776 16502
rect 49568 16436 49616 16492
rect 49672 16436 49720 16492
rect 49512 16426 49776 16436
rect 49868 16324 49924 16334
rect 49868 16210 49924 16268
rect 49868 16158 49870 16210
rect 49922 16158 49924 16210
rect 49868 16146 49924 16158
rect 49420 16100 49476 16110
rect 49420 16006 49476 16044
rect 49980 15316 50036 16604
rect 49980 15250 50036 15260
rect 50428 15876 50484 15886
rect 49512 14924 49776 14934
rect 49568 14868 49616 14924
rect 49672 14868 49720 14924
rect 49512 14858 49776 14868
rect 49308 14700 49476 14756
rect 49420 14642 49476 14700
rect 49420 14590 49422 14642
rect 49474 14590 49476 14642
rect 49420 14578 49476 14590
rect 48748 14530 48804 14542
rect 48748 14478 48750 14530
rect 48802 14478 48804 14530
rect 48412 14308 48468 14318
rect 48412 13970 48468 14252
rect 48748 14084 48804 14478
rect 48748 14018 48804 14028
rect 49308 14530 49364 14542
rect 49308 14478 49310 14530
rect 49362 14478 49364 14530
rect 48412 13918 48414 13970
rect 48466 13918 48468 13970
rect 48412 13906 48468 13918
rect 48636 13858 48692 13870
rect 48636 13806 48638 13858
rect 48690 13806 48692 13858
rect 48636 13636 48692 13806
rect 49308 13860 49364 14478
rect 49980 14420 50036 14430
rect 49868 14418 50036 14420
rect 49868 14366 49982 14418
rect 50034 14366 50036 14418
rect 49868 14364 50036 14366
rect 49532 13860 49588 13870
rect 49868 13860 49924 14364
rect 49980 14354 50036 14364
rect 50316 14420 50372 14430
rect 50316 14326 50372 14364
rect 50092 14306 50148 14318
rect 50092 14254 50094 14306
rect 50146 14254 50148 14306
rect 50092 14084 50148 14254
rect 50092 14018 50148 14028
rect 49308 13858 49924 13860
rect 49308 13806 49534 13858
rect 49586 13806 49924 13858
rect 49308 13804 49924 13806
rect 50428 13860 50484 15820
rect 50540 15426 50596 16828
rect 50652 16772 50708 16782
rect 50652 16212 50708 16716
rect 50876 16772 50932 18732
rect 51100 18452 51156 18462
rect 50988 16884 51044 16894
rect 50988 16790 51044 16828
rect 50876 16706 50932 16716
rect 50652 16210 50820 16212
rect 50652 16158 50654 16210
rect 50706 16158 50820 16210
rect 50652 16156 50820 16158
rect 50652 16146 50708 16156
rect 50540 15374 50542 15426
rect 50594 15374 50596 15426
rect 50540 15316 50596 15374
rect 50652 15428 50708 15438
rect 50652 15334 50708 15372
rect 50540 15250 50596 15260
rect 50764 15204 50820 16156
rect 50876 15876 50932 15886
rect 50876 15538 50932 15820
rect 50876 15486 50878 15538
rect 50930 15486 50932 15538
rect 50876 15474 50932 15486
rect 50764 15138 50820 15148
rect 51100 14530 51156 18396
rect 51212 18228 51268 31500
rect 51436 31554 51492 31892
rect 51436 31502 51438 31554
rect 51490 31502 51492 31554
rect 51436 30996 51492 31502
rect 51436 30930 51492 30940
rect 51548 30994 51604 31006
rect 51548 30942 51550 30994
rect 51602 30942 51604 30994
rect 51548 30884 51604 30942
rect 51548 30818 51604 30828
rect 51324 29538 51380 29550
rect 51324 29486 51326 29538
rect 51378 29486 51380 29538
rect 51324 29204 51380 29486
rect 51324 29138 51380 29148
rect 51436 29426 51492 29438
rect 51436 29374 51438 29426
rect 51490 29374 51492 29426
rect 51436 28644 51492 29374
rect 51436 28578 51492 28588
rect 51660 26908 51716 31892
rect 52220 31668 52276 31678
rect 52220 31574 52276 31612
rect 51772 31556 51828 31566
rect 51772 31462 51828 31500
rect 52780 31556 52836 33068
rect 53340 31948 53396 35868
rect 55356 35700 55412 35710
rect 55356 35606 55412 35644
rect 55916 35700 55972 35710
rect 55692 35026 55748 35038
rect 55692 34974 55694 35026
rect 55746 34974 55748 35026
rect 55244 34914 55300 34926
rect 55244 34862 55246 34914
rect 55298 34862 55300 34914
rect 53900 34244 53956 34254
rect 55132 34244 55188 34254
rect 53900 34242 54068 34244
rect 53900 34190 53902 34242
rect 53954 34190 54068 34242
rect 53900 34188 54068 34190
rect 53900 34178 53956 34188
rect 53788 34130 53844 34142
rect 53788 34078 53790 34130
rect 53842 34078 53844 34130
rect 53788 33458 53844 34078
rect 53788 33406 53790 33458
rect 53842 33406 53844 33458
rect 53788 32676 53844 33406
rect 53900 33906 53956 33918
rect 53900 33854 53902 33906
rect 53954 33854 53956 33906
rect 53900 33236 53956 33854
rect 54012 33348 54068 34188
rect 55132 34150 55188 34188
rect 55244 34018 55300 34862
rect 55244 33966 55246 34018
rect 55298 33966 55300 34018
rect 55244 33954 55300 33966
rect 55692 34020 55748 34974
rect 55916 34804 55972 35644
rect 56028 35698 56084 35710
rect 56028 35646 56030 35698
rect 56082 35646 56084 35698
rect 56028 35252 56084 35646
rect 56028 35186 56084 35196
rect 56140 35698 56196 35710
rect 56140 35646 56142 35698
rect 56194 35646 56196 35698
rect 56028 34916 56084 34926
rect 56140 34916 56196 35646
rect 58044 35700 58100 35710
rect 56588 35588 56644 35598
rect 56588 35494 56644 35532
rect 57484 35588 57540 35598
rect 57484 35494 57540 35532
rect 58044 35586 58100 35644
rect 58044 35534 58046 35586
rect 58098 35534 58100 35586
rect 58044 35522 58100 35534
rect 57036 35476 57092 35486
rect 57036 35026 57092 35420
rect 57708 35476 57764 35486
rect 57708 35382 57764 35420
rect 57036 34974 57038 35026
rect 57090 34974 57092 35026
rect 57036 34962 57092 34974
rect 57260 35252 57316 35262
rect 56588 34916 56644 34926
rect 56028 34914 56644 34916
rect 56028 34862 56030 34914
rect 56082 34862 56590 34914
rect 56642 34862 56644 34914
rect 56028 34860 56644 34862
rect 56028 34850 56084 34860
rect 56588 34850 56644 34860
rect 57260 34914 57316 35196
rect 57260 34862 57262 34914
rect 57314 34862 57316 34914
rect 57260 34850 57316 34862
rect 57372 35138 57428 35150
rect 57372 35086 57374 35138
rect 57426 35086 57428 35138
rect 55916 34738 55972 34748
rect 56812 34804 56868 34814
rect 56812 34710 56868 34748
rect 54908 33908 54964 33918
rect 54124 33348 54180 33358
rect 54572 33348 54628 33358
rect 54908 33348 54964 33852
rect 55692 33458 55748 33964
rect 55692 33406 55694 33458
rect 55746 33406 55748 33458
rect 55692 33394 55748 33406
rect 54012 33346 54292 33348
rect 54012 33294 54126 33346
rect 54178 33294 54292 33346
rect 54012 33292 54292 33294
rect 54124 33282 54180 33292
rect 53900 33170 53956 33180
rect 53788 32610 53844 32620
rect 52780 31490 52836 31500
rect 52892 31892 53396 31948
rect 53788 32452 53844 32462
rect 51884 30994 51940 31006
rect 51884 30942 51886 30994
rect 51938 30942 51940 30994
rect 51884 29204 51940 30942
rect 52444 30884 52500 30894
rect 52444 29652 52500 30828
rect 52444 29586 52500 29596
rect 52892 29428 52948 31892
rect 53788 31666 53844 32396
rect 54124 32004 54180 32014
rect 54124 31778 54180 31948
rect 54124 31726 54126 31778
rect 54178 31726 54180 31778
rect 54124 31714 54180 31726
rect 53788 31614 53790 31666
rect 53842 31614 53844 31666
rect 53788 31444 53844 31614
rect 54012 31668 54068 31678
rect 53788 31378 53844 31388
rect 53900 31556 53956 31566
rect 53564 30884 53620 30894
rect 53900 30884 53956 31500
rect 53564 30882 53956 30884
rect 53564 30830 53566 30882
rect 53618 30830 53956 30882
rect 53564 30828 53956 30830
rect 54012 31108 54068 31612
rect 54236 31220 54292 33292
rect 54572 33346 54964 33348
rect 54572 33294 54574 33346
rect 54626 33294 54964 33346
rect 54572 33292 54964 33294
rect 56140 33346 56196 33358
rect 56140 33294 56142 33346
rect 56194 33294 56196 33346
rect 54572 33282 54628 33292
rect 56028 32788 56084 32798
rect 56140 32788 56196 33294
rect 56588 33348 56644 33358
rect 56588 33254 56644 33292
rect 57148 33346 57204 33358
rect 57148 33294 57150 33346
rect 57202 33294 57204 33346
rect 57148 33236 57204 33294
rect 57148 33170 57204 33180
rect 56028 32786 56196 32788
rect 56028 32734 56030 32786
rect 56082 32734 56196 32786
rect 56028 32732 56196 32734
rect 56028 32722 56084 32732
rect 55916 32674 55972 32686
rect 55916 32622 55918 32674
rect 55970 32622 55972 32674
rect 55356 32562 55412 32574
rect 55356 32510 55358 32562
rect 55410 32510 55412 32562
rect 54348 32450 54404 32462
rect 54348 32398 54350 32450
rect 54402 32398 54404 32450
rect 54348 31948 54404 32398
rect 54572 32338 54628 32350
rect 54572 32286 54574 32338
rect 54626 32286 54628 32338
rect 54572 32004 54628 32286
rect 54348 31892 54516 31948
rect 54572 31938 54628 31948
rect 54908 32338 54964 32350
rect 54908 32286 54910 32338
rect 54962 32286 54964 32338
rect 54908 31948 54964 32286
rect 55356 32004 55412 32510
rect 55692 32564 55748 32574
rect 55692 32470 55748 32508
rect 54908 31892 55076 31948
rect 54460 31668 54516 31892
rect 54908 31668 54964 31678
rect 54460 31666 54964 31668
rect 54460 31614 54910 31666
rect 54962 31614 54964 31666
rect 54460 31612 54964 31614
rect 54348 31220 54404 31230
rect 54236 31218 54404 31220
rect 54236 31166 54350 31218
rect 54402 31166 54404 31218
rect 54236 31164 54404 31166
rect 54348 31154 54404 31164
rect 53564 30324 53620 30828
rect 53564 30258 53620 30268
rect 53900 30212 53956 30222
rect 54012 30212 54068 31052
rect 54236 30996 54292 31006
rect 54236 30902 54292 30940
rect 54460 30994 54516 31006
rect 54460 30942 54462 30994
rect 54514 30942 54516 30994
rect 53900 30210 54068 30212
rect 53900 30158 53902 30210
rect 53954 30158 54068 30210
rect 53900 30156 54068 30158
rect 54236 30772 54292 30782
rect 54236 30210 54292 30716
rect 54460 30660 54516 30942
rect 54684 30884 54740 30894
rect 54684 30790 54740 30828
rect 54796 30772 54852 31612
rect 54908 31602 54964 31612
rect 54908 30996 54964 31006
rect 55020 30996 55076 31892
rect 55356 31778 55412 31948
rect 55356 31726 55358 31778
rect 55410 31726 55412 31778
rect 55356 31714 55412 31726
rect 55580 31780 55636 31790
rect 54908 30994 55076 30996
rect 54908 30942 54910 30994
rect 54962 30942 55076 30994
rect 54908 30940 55076 30942
rect 55356 31108 55412 31118
rect 54908 30930 54964 30940
rect 54796 30706 54852 30716
rect 54460 30604 54740 30660
rect 54684 30548 54740 30604
rect 55356 30548 55412 31052
rect 54684 30492 54852 30548
rect 54236 30158 54238 30210
rect 54290 30158 54292 30210
rect 53900 30146 53956 30156
rect 54236 30146 54292 30158
rect 54796 30434 54852 30492
rect 55356 30482 55412 30492
rect 55580 30884 55636 31724
rect 55916 31556 55972 32622
rect 56364 32564 56420 32574
rect 56364 31948 56420 32508
rect 56252 31892 56420 31948
rect 56140 31780 56196 31790
rect 56140 31686 56196 31724
rect 55804 30884 55860 30894
rect 54796 30382 54798 30434
rect 54850 30382 54852 30434
rect 54796 30212 54852 30382
rect 55580 30434 55636 30828
rect 55580 30382 55582 30434
rect 55634 30382 55636 30434
rect 55580 30370 55636 30382
rect 55692 30882 55860 30884
rect 55692 30830 55806 30882
rect 55858 30830 55860 30882
rect 55692 30828 55860 30830
rect 55692 30324 55748 30828
rect 55804 30818 55860 30828
rect 55916 30772 55972 31500
rect 55916 30660 55972 30716
rect 55692 30258 55748 30268
rect 55804 30604 55972 30660
rect 56252 30882 56308 31892
rect 56812 31668 56868 31678
rect 56812 31574 56868 31612
rect 57260 31556 57316 31566
rect 57260 31462 57316 31500
rect 56252 30830 56254 30882
rect 56306 30830 56308 30882
rect 54796 30146 54852 30156
rect 54684 30100 54740 30110
rect 54684 30006 54740 30044
rect 55692 30100 55748 30110
rect 55692 30006 55748 30044
rect 53452 29986 53508 29998
rect 53452 29934 53454 29986
rect 53506 29934 53508 29986
rect 53452 29876 53508 29934
rect 53452 29810 53508 29820
rect 54012 29986 54068 29998
rect 54012 29934 54014 29986
rect 54066 29934 54068 29986
rect 54012 29876 54068 29934
rect 54012 29810 54068 29820
rect 54796 29986 54852 29998
rect 54796 29934 54798 29986
rect 54850 29934 54852 29986
rect 54796 29876 54852 29934
rect 55580 29988 55636 29998
rect 55580 29894 55636 29932
rect 54796 29810 54852 29820
rect 51884 29138 51940 29148
rect 52220 29372 52948 29428
rect 53004 29538 53060 29550
rect 53004 29486 53006 29538
rect 53058 29486 53060 29538
rect 52220 26908 52276 29372
rect 52668 29204 52724 29214
rect 52780 29204 52836 29214
rect 52724 29202 52836 29204
rect 52724 29150 52782 29202
rect 52834 29150 52836 29202
rect 52724 29148 52836 29150
rect 52332 28756 52388 28766
rect 52332 28662 52388 28700
rect 52444 28418 52500 28430
rect 52444 28366 52446 28418
rect 52498 28366 52500 28418
rect 52444 27972 52500 28366
rect 52444 27906 52500 27916
rect 52556 27858 52612 27870
rect 52556 27806 52558 27858
rect 52610 27806 52612 27858
rect 52556 27188 52612 27806
rect 52668 27634 52724 29148
rect 52780 29138 52836 29148
rect 53004 28756 53060 29486
rect 54908 29540 54964 29550
rect 54908 29446 54964 29484
rect 54572 29428 54628 29438
rect 54572 29334 54628 29372
rect 54684 29426 54740 29438
rect 54684 29374 54686 29426
rect 54738 29374 54740 29426
rect 53004 28690 53060 28700
rect 53116 29202 53172 29214
rect 53116 29150 53118 29202
rect 53170 29150 53172 29202
rect 53116 28532 53172 29150
rect 54684 28756 54740 29374
rect 55132 29428 55188 29438
rect 55132 29426 55412 29428
rect 55132 29374 55134 29426
rect 55186 29374 55412 29426
rect 55132 29372 55412 29374
rect 55132 29362 55188 29372
rect 54460 28700 54740 28756
rect 54012 28642 54068 28654
rect 54012 28590 54014 28642
rect 54066 28590 54068 28642
rect 53116 28466 53172 28476
rect 53452 28530 53508 28542
rect 53452 28478 53454 28530
rect 53506 28478 53508 28530
rect 52892 27858 52948 27870
rect 52892 27806 52894 27858
rect 52946 27806 52948 27858
rect 52892 27748 52948 27806
rect 52892 27682 52948 27692
rect 52668 27582 52670 27634
rect 52722 27582 52724 27634
rect 52668 27570 52724 27582
rect 53452 27188 53508 28478
rect 53676 28418 53732 28430
rect 53900 28420 53956 28430
rect 53676 28366 53678 28418
rect 53730 28366 53732 28418
rect 53564 28196 53620 28206
rect 53564 27858 53620 28140
rect 53564 27806 53566 27858
rect 53618 27806 53620 27858
rect 53564 27794 53620 27806
rect 53676 27412 53732 28366
rect 52556 27132 53508 27188
rect 53564 27356 53732 27412
rect 53788 28418 53956 28420
rect 53788 28366 53902 28418
rect 53954 28366 53956 28418
rect 53788 28364 53956 28366
rect 53788 27970 53844 28364
rect 53900 28354 53956 28364
rect 54012 28420 54068 28590
rect 54012 28354 54068 28364
rect 54460 28420 54516 28700
rect 55356 28644 55412 29372
rect 55356 28588 55636 28644
rect 54572 28532 54628 28542
rect 54572 28438 54628 28476
rect 54796 28532 54852 28542
rect 55244 28532 55300 28542
rect 54796 28530 55300 28532
rect 54796 28478 54798 28530
rect 54850 28478 55246 28530
rect 55298 28478 55300 28530
rect 54796 28476 55300 28478
rect 54796 28466 54852 28476
rect 55244 28466 55300 28476
rect 55580 28530 55636 28588
rect 55580 28478 55582 28530
rect 55634 28478 55636 28530
rect 54460 28354 54516 28364
rect 54684 28418 54740 28430
rect 54684 28366 54686 28418
rect 54738 28366 54740 28418
rect 53788 27918 53790 27970
rect 53842 27918 53844 27970
rect 51436 26852 51716 26908
rect 52108 26852 52276 26908
rect 52668 26962 52724 26974
rect 52668 26910 52670 26962
rect 52722 26910 52724 26962
rect 52332 26852 52388 26862
rect 51436 22484 51492 26852
rect 51436 22258 51492 22428
rect 51436 22206 51438 22258
rect 51490 22206 51492 22258
rect 51436 22194 51492 22206
rect 51772 22260 51828 22270
rect 52108 22260 52164 26852
rect 52332 26758 52388 26796
rect 52668 26516 52724 26910
rect 52780 26908 52836 27132
rect 53564 27076 53620 27356
rect 53788 27300 53844 27918
rect 54348 28196 54404 28206
rect 54348 27858 54404 28140
rect 54684 28084 54740 28366
rect 55468 28420 55524 28430
rect 55468 28326 55524 28364
rect 54684 28028 54852 28084
rect 54572 27972 54628 27982
rect 54572 27878 54628 27916
rect 54348 27806 54350 27858
rect 54402 27806 54404 27858
rect 54348 27794 54404 27806
rect 54684 27858 54740 27870
rect 54684 27806 54686 27858
rect 54738 27806 54740 27858
rect 54684 27748 54740 27806
rect 54684 27682 54740 27692
rect 53788 27234 53844 27244
rect 54012 27356 54628 27412
rect 53900 27076 53956 27086
rect 53564 27010 53620 27020
rect 53676 27074 53956 27076
rect 53676 27022 53902 27074
rect 53954 27022 53956 27074
rect 53676 27020 53956 27022
rect 52780 26852 52948 26908
rect 52668 26450 52724 26460
rect 52780 26628 52836 26638
rect 52668 26292 52724 26302
rect 52668 26198 52724 26236
rect 52556 24722 52612 24734
rect 52556 24670 52558 24722
rect 52610 24670 52612 24722
rect 52444 24610 52500 24622
rect 52444 24558 52446 24610
rect 52498 24558 52500 24610
rect 52444 23828 52500 24558
rect 52220 23826 52500 23828
rect 52220 23774 52446 23826
rect 52498 23774 52500 23826
rect 52220 23772 52500 23774
rect 52220 22596 52276 23772
rect 52444 23762 52500 23772
rect 52556 23716 52612 24670
rect 52780 23938 52836 26572
rect 52780 23886 52782 23938
rect 52834 23886 52836 23938
rect 52780 23874 52836 23886
rect 52892 26292 52948 26852
rect 53564 26850 53620 26862
rect 53564 26798 53566 26850
rect 53618 26798 53620 26850
rect 53564 26628 53620 26798
rect 53564 26562 53620 26572
rect 53452 26516 53508 26526
rect 53116 26292 53172 26302
rect 52892 26290 53172 26292
rect 52892 26238 53118 26290
rect 53170 26238 53172 26290
rect 52892 26236 53172 26238
rect 52556 23622 52612 23660
rect 52556 23380 52612 23390
rect 52220 22530 52276 22540
rect 52332 23324 52556 23380
rect 52108 22204 52276 22260
rect 51772 22166 51828 22204
rect 51884 21924 51940 21934
rect 51940 21868 52052 21924
rect 51884 21858 51940 21868
rect 51548 19012 51604 19022
rect 51548 19010 51940 19012
rect 51548 18958 51550 19010
rect 51602 18958 51940 19010
rect 51548 18956 51940 18958
rect 51548 18946 51604 18956
rect 51324 18788 51380 18798
rect 51324 18674 51380 18732
rect 51324 18622 51326 18674
rect 51378 18622 51380 18674
rect 51324 18610 51380 18622
rect 51660 18676 51716 18686
rect 51660 18582 51716 18620
rect 51884 18562 51940 18956
rect 51884 18510 51886 18562
rect 51938 18510 51940 18562
rect 51436 18450 51492 18462
rect 51436 18398 51438 18450
rect 51490 18398 51492 18450
rect 51436 18340 51492 18398
rect 51436 18274 51492 18284
rect 51548 18338 51604 18350
rect 51548 18286 51550 18338
rect 51602 18286 51604 18338
rect 51212 17780 51268 18172
rect 51212 17668 51268 17724
rect 51324 17668 51380 17678
rect 51212 17666 51380 17668
rect 51212 17614 51326 17666
rect 51378 17614 51380 17666
rect 51212 17612 51380 17614
rect 51324 17602 51380 17612
rect 51436 17556 51492 17566
rect 51436 17462 51492 17500
rect 51324 17332 51380 17342
rect 51324 16210 51380 17276
rect 51548 16322 51604 18286
rect 51660 17442 51716 17454
rect 51660 17390 51662 17442
rect 51714 17390 51716 17442
rect 51660 17108 51716 17390
rect 51660 16882 51716 17052
rect 51884 16996 51940 18510
rect 51884 16930 51940 16940
rect 51660 16830 51662 16882
rect 51714 16830 51716 16882
rect 51660 16818 51716 16830
rect 51548 16270 51550 16322
rect 51602 16270 51604 16322
rect 51548 16258 51604 16270
rect 51884 16772 51940 16782
rect 51884 16322 51940 16716
rect 51884 16270 51886 16322
rect 51938 16270 51940 16322
rect 51884 16258 51940 16270
rect 51324 16158 51326 16210
rect 51378 16158 51380 16210
rect 51324 16146 51380 16158
rect 51212 15428 51268 15438
rect 51212 15334 51268 15372
rect 51660 15316 51716 15326
rect 51660 15222 51716 15260
rect 51996 15148 52052 21868
rect 51100 14478 51102 14530
rect 51154 14478 51156 14530
rect 51100 14466 51156 14478
rect 51772 15092 52052 15148
rect 52108 21812 52164 21822
rect 50764 14420 50820 14430
rect 50764 14326 50820 14364
rect 50876 14308 50932 14318
rect 50876 14214 50932 14252
rect 49532 13794 49588 13804
rect 50428 13794 50484 13804
rect 48748 13746 48804 13758
rect 48748 13694 48750 13746
rect 48802 13694 48804 13746
rect 48748 13636 48804 13694
rect 49980 13746 50036 13758
rect 49980 13694 49982 13746
rect 50034 13694 50036 13746
rect 49868 13636 49924 13646
rect 48748 13634 49924 13636
rect 48748 13582 49870 13634
rect 49922 13582 49924 13634
rect 48748 13580 49924 13582
rect 48636 13570 48692 13580
rect 48300 13346 48356 13356
rect 48972 13074 49028 13580
rect 49868 13570 49924 13580
rect 49980 13636 50036 13694
rect 49980 13570 50036 13580
rect 49512 13356 49776 13366
rect 49568 13300 49616 13356
rect 49672 13300 49720 13356
rect 49512 13290 49776 13300
rect 48972 13022 48974 13074
rect 49026 13022 49028 13074
rect 48972 13010 49028 13022
rect 50988 13076 51044 13086
rect 50988 12982 51044 13020
rect 49644 12964 49700 12974
rect 49644 12870 49700 12908
rect 49868 12964 49924 12974
rect 50876 12964 50932 12974
rect 49868 12962 50148 12964
rect 49868 12910 49870 12962
rect 49922 12910 50148 12962
rect 49868 12908 50148 12910
rect 49868 12898 49924 12908
rect 50092 12852 50148 12908
rect 48860 12740 48916 12750
rect 48860 12402 48916 12684
rect 48860 12350 48862 12402
rect 48914 12350 48916 12402
rect 48860 12338 48916 12350
rect 48636 12292 48692 12302
rect 48636 12198 48692 12236
rect 49756 12292 49812 12302
rect 48524 12180 48580 12190
rect 48412 12178 48580 12180
rect 48412 12126 48526 12178
rect 48578 12126 48580 12178
rect 48412 12124 48580 12126
rect 48412 12068 48468 12124
rect 48524 12114 48580 12124
rect 49756 12178 49812 12236
rect 49756 12126 49758 12178
rect 49810 12126 49812 12178
rect 49756 12114 49812 12126
rect 48188 11844 48244 11854
rect 46956 11396 47012 11406
rect 46956 10610 47012 11340
rect 46956 10558 46958 10610
rect 47010 10558 47012 10610
rect 46956 10546 47012 10558
rect 47292 10724 47348 10734
rect 47292 10610 47348 10668
rect 47292 10558 47294 10610
rect 47346 10558 47348 10610
rect 47292 10546 47348 10558
rect 47516 10724 47572 10734
rect 47516 8370 47572 10668
rect 47516 8318 47518 8370
rect 47570 8318 47572 8370
rect 47516 8306 47572 8318
rect 47404 8260 47460 8270
rect 47404 8166 47460 8204
rect 48076 8258 48132 8270
rect 48076 8206 48078 8258
rect 48130 8206 48132 8258
rect 47628 8148 47684 8158
rect 47628 8054 47684 8092
rect 45388 7186 45444 7196
rect 45948 6804 46004 6814
rect 45948 6690 46004 6748
rect 45948 6638 45950 6690
rect 46002 6638 46004 6690
rect 45948 6626 46004 6638
rect 46620 6804 46676 6814
rect 46844 6804 46900 7756
rect 48076 7698 48132 8206
rect 48076 7646 48078 7698
rect 48130 7646 48132 7698
rect 48076 7634 48132 7646
rect 48188 7700 48244 11788
rect 48300 10610 48356 10622
rect 48300 10558 48302 10610
rect 48354 10558 48356 10610
rect 48300 9714 48356 10558
rect 48412 10386 48468 12012
rect 49868 12068 49924 12078
rect 49868 11974 49924 12012
rect 50092 11954 50148 12796
rect 50652 12740 50708 12750
rect 50652 12646 50708 12684
rect 50876 12738 50932 12908
rect 51100 12852 51156 12862
rect 51100 12758 51156 12796
rect 51324 12852 51380 12862
rect 50876 12686 50878 12738
rect 50930 12686 50932 12738
rect 50876 12292 50932 12686
rect 50876 12226 50932 12236
rect 51324 12180 51380 12796
rect 51324 12114 51380 12124
rect 50092 11902 50094 11954
rect 50146 11902 50148 11954
rect 50092 11890 50148 11902
rect 49512 11788 49776 11798
rect 49568 11732 49616 11788
rect 49672 11732 49720 11788
rect 49512 11722 49776 11732
rect 48860 11396 48916 11406
rect 48860 11302 48916 11340
rect 49308 11394 49364 11406
rect 49308 11342 49310 11394
rect 49362 11342 49364 11394
rect 48748 11284 48804 11294
rect 48748 11190 48804 11228
rect 48636 11172 48692 11182
rect 48412 10334 48414 10386
rect 48466 10334 48468 10386
rect 48412 10322 48468 10334
rect 48524 11170 48692 11172
rect 48524 11118 48638 11170
rect 48690 11118 48692 11170
rect 48524 11116 48692 11118
rect 48524 9938 48580 11116
rect 48636 11106 48692 11116
rect 49308 10836 49364 11342
rect 51548 11396 51604 11406
rect 51548 11302 51604 11340
rect 50988 11172 51044 11182
rect 49420 10836 49476 10846
rect 49308 10834 49476 10836
rect 49308 10782 49422 10834
rect 49474 10782 49476 10834
rect 49308 10780 49476 10782
rect 49420 10770 49476 10780
rect 48524 9886 48526 9938
rect 48578 9886 48580 9938
rect 48524 9874 48580 9886
rect 48636 10724 48692 10734
rect 48636 9826 48692 10668
rect 49644 10724 49700 10734
rect 49644 10630 49700 10668
rect 49756 10612 49812 10622
rect 49756 10610 49924 10612
rect 49756 10558 49758 10610
rect 49810 10558 49924 10610
rect 49756 10556 49924 10558
rect 49756 10546 49812 10556
rect 49512 10220 49776 10230
rect 49568 10164 49616 10220
rect 49672 10164 49720 10220
rect 49512 10154 49776 10164
rect 48636 9774 48638 9826
rect 48690 9774 48692 9826
rect 48636 9762 48692 9774
rect 49756 9826 49812 9838
rect 49756 9774 49758 9826
rect 49810 9774 49812 9826
rect 48300 9662 48302 9714
rect 48354 9662 48356 9714
rect 48300 9380 48356 9662
rect 48300 9314 48356 9324
rect 49196 9602 49252 9614
rect 49196 9550 49198 9602
rect 49250 9550 49252 9602
rect 49196 9268 49252 9550
rect 48748 9156 48804 9166
rect 48748 9062 48804 9100
rect 49196 8708 49252 9212
rect 49420 9156 49476 9166
rect 49420 9062 49476 9100
rect 49756 9156 49812 9774
rect 49868 9380 49924 10556
rect 50316 10500 50372 10510
rect 50316 10406 50372 10444
rect 50764 10500 50820 10510
rect 50764 10276 50820 10444
rect 50988 10388 51044 11116
rect 50988 10322 51044 10332
rect 49868 9314 49924 9324
rect 49980 9826 50036 9838
rect 49980 9774 49982 9826
rect 50034 9774 50036 9826
rect 49980 9268 50036 9774
rect 50540 9716 50596 9726
rect 49980 9174 50036 9212
rect 50316 9602 50372 9614
rect 50316 9550 50318 9602
rect 50370 9550 50372 9602
rect 49756 9090 49812 9100
rect 49196 8642 49252 8652
rect 49512 8652 49776 8662
rect 49568 8596 49616 8652
rect 49672 8596 49720 8652
rect 49512 8586 49776 8596
rect 50316 8260 50372 9550
rect 50540 8370 50596 9660
rect 50764 9716 50820 10220
rect 50988 9828 51044 9838
rect 50876 9716 50932 9726
rect 50764 9714 50932 9716
rect 50764 9662 50878 9714
rect 50930 9662 50932 9714
rect 50764 9660 50932 9662
rect 50764 9044 50820 9660
rect 50876 9650 50932 9660
rect 50988 9714 51044 9772
rect 51548 9828 51604 9838
rect 51548 9734 51604 9772
rect 50988 9662 50990 9714
rect 51042 9662 51044 9714
rect 50988 9604 51044 9662
rect 50988 9538 51044 9548
rect 51212 9602 51268 9614
rect 51212 9550 51214 9602
rect 51266 9550 51268 9602
rect 50876 9156 50932 9166
rect 50876 9062 50932 9100
rect 50764 8978 50820 8988
rect 51212 9042 51268 9550
rect 51212 8990 51214 9042
rect 51266 8990 51268 9042
rect 51100 8484 51156 8494
rect 51212 8484 51268 8990
rect 51100 8482 51268 8484
rect 51100 8430 51102 8482
rect 51154 8430 51268 8482
rect 51100 8428 51268 8430
rect 51772 8428 51828 15092
rect 51996 14644 52052 14654
rect 51996 14550 52052 14588
rect 51996 11394 52052 11406
rect 51996 11342 51998 11394
rect 52050 11342 52052 11394
rect 51996 11172 52052 11342
rect 51996 11106 52052 11116
rect 52108 9828 52164 21756
rect 52220 20692 52276 22204
rect 52332 22258 52388 23324
rect 52444 23156 52500 23166
rect 52444 22708 52500 23100
rect 52556 23042 52612 23324
rect 52892 23266 52948 26236
rect 53116 26226 53172 26236
rect 53452 25618 53508 26460
rect 53564 26292 53620 26302
rect 53676 26292 53732 27020
rect 53900 27010 53956 27020
rect 53788 26852 53844 26862
rect 53788 26850 53956 26852
rect 53788 26798 53790 26850
rect 53842 26798 53956 26850
rect 53788 26796 53956 26798
rect 53788 26786 53844 26796
rect 53564 26290 53732 26292
rect 53564 26238 53566 26290
rect 53618 26238 53732 26290
rect 53564 26236 53732 26238
rect 53788 26628 53844 26638
rect 53564 26226 53620 26236
rect 53452 25566 53454 25618
rect 53506 25566 53508 25618
rect 53452 25554 53508 25566
rect 53340 25508 53396 25518
rect 53340 24834 53396 25452
rect 53340 24782 53342 24834
rect 53394 24782 53396 24834
rect 53340 24770 53396 24782
rect 53788 24836 53844 26572
rect 53900 25508 53956 26796
rect 54012 26850 54068 27356
rect 54572 27298 54628 27356
rect 54572 27246 54574 27298
rect 54626 27246 54628 27298
rect 54572 27234 54628 27246
rect 54012 26798 54014 26850
rect 54066 26798 54068 26850
rect 54012 25620 54068 26798
rect 54348 27188 54404 27198
rect 54236 25620 54292 25630
rect 54012 25618 54292 25620
rect 54012 25566 54238 25618
rect 54290 25566 54292 25618
rect 54012 25564 54292 25566
rect 54236 25554 54292 25564
rect 53900 25414 53956 25452
rect 54348 24948 54404 27132
rect 54684 26964 54740 26974
rect 54684 26870 54740 26908
rect 54124 24892 54404 24948
rect 53900 24836 53956 24846
rect 53788 24834 53956 24836
rect 53788 24782 53902 24834
rect 53954 24782 53956 24834
rect 53788 24780 53956 24782
rect 53900 24770 53956 24780
rect 54012 24722 54068 24734
rect 54012 24670 54014 24722
rect 54066 24670 54068 24722
rect 54012 24388 54068 24670
rect 53900 24332 54068 24388
rect 53452 23940 53508 23950
rect 53676 23940 53732 23950
rect 52892 23214 52894 23266
rect 52946 23214 52948 23266
rect 52892 23202 52948 23214
rect 53004 23938 53508 23940
rect 53004 23886 53454 23938
rect 53506 23886 53508 23938
rect 53004 23884 53508 23886
rect 52556 22990 52558 23042
rect 52610 22990 52612 23042
rect 52556 22978 52612 22990
rect 53004 22932 53060 23884
rect 53452 23874 53508 23884
rect 53564 23938 53732 23940
rect 53564 23886 53678 23938
rect 53730 23886 53732 23938
rect 53564 23884 53732 23886
rect 53452 23380 53508 23390
rect 53452 23286 53508 23324
rect 53564 23378 53620 23884
rect 53676 23874 53732 23884
rect 53564 23326 53566 23378
rect 53618 23326 53620 23378
rect 53564 23314 53620 23326
rect 53788 23716 53844 23726
rect 53676 23266 53732 23278
rect 53676 23214 53678 23266
rect 53730 23214 53732 23266
rect 53676 23156 53732 23214
rect 53788 23266 53844 23660
rect 53788 23214 53790 23266
rect 53842 23214 53844 23266
rect 53788 23202 53844 23214
rect 53900 23266 53956 24332
rect 54012 24164 54068 24174
rect 54124 24164 54180 24892
rect 54012 24162 54180 24164
rect 54012 24110 54014 24162
rect 54066 24110 54180 24162
rect 54012 24108 54180 24110
rect 54348 24722 54404 24734
rect 54348 24670 54350 24722
rect 54402 24670 54404 24722
rect 54012 24098 54068 24108
rect 54348 23716 54404 24670
rect 54348 23650 54404 23660
rect 53900 23214 53902 23266
rect 53954 23214 53956 23266
rect 53676 23090 53732 23100
rect 52668 22876 53060 22932
rect 52444 22652 52612 22708
rect 52332 22206 52334 22258
rect 52386 22206 52388 22258
rect 52332 21700 52388 22206
rect 52444 22148 52500 22186
rect 52556 22148 52612 22652
rect 52668 22370 52724 22876
rect 53900 22596 53956 23214
rect 53900 22530 53956 22540
rect 54348 22484 54404 22494
rect 54796 22484 54852 28028
rect 55132 27636 55188 27646
rect 54908 27634 55188 27636
rect 54908 27582 55134 27634
rect 55186 27582 55188 27634
rect 54908 27580 55188 27582
rect 54908 27298 54964 27580
rect 55132 27570 55188 27580
rect 54908 27246 54910 27298
rect 54962 27246 54964 27298
rect 54908 27234 54964 27246
rect 55356 27188 55412 27198
rect 55580 27188 55636 28478
rect 55804 27748 55860 30604
rect 55916 30212 55972 30222
rect 56252 30212 56308 30830
rect 55916 29314 55972 30156
rect 56140 30156 56308 30212
rect 56364 31444 56420 31454
rect 56364 30324 56420 31388
rect 56140 30100 56196 30156
rect 56140 30034 56196 30044
rect 56252 29986 56308 29998
rect 56252 29934 56254 29986
rect 56306 29934 56308 29986
rect 56252 29876 56308 29934
rect 56252 29810 56308 29820
rect 55916 29262 55918 29314
rect 55970 29262 55972 29314
rect 55916 29250 55972 29262
rect 56028 29428 56084 29438
rect 56028 28642 56084 29372
rect 56028 28590 56030 28642
rect 56082 28590 56084 28642
rect 55916 27748 55972 27758
rect 55804 27746 55972 27748
rect 55804 27694 55918 27746
rect 55970 27694 55972 27746
rect 55804 27692 55972 27694
rect 55412 27132 55636 27188
rect 55356 27122 55412 27132
rect 55916 26852 55972 27692
rect 55916 26786 55972 26796
rect 55580 23156 55636 23166
rect 55580 23062 55636 23100
rect 56028 22820 56084 28590
rect 56252 29428 56308 29438
rect 56140 27300 56196 27310
rect 56252 27300 56308 29372
rect 56140 27298 56308 27300
rect 56140 27246 56142 27298
rect 56194 27246 56308 27298
rect 56140 27244 56308 27246
rect 56140 27234 56196 27244
rect 56364 27188 56420 30268
rect 57148 30322 57204 30334
rect 57148 30270 57150 30322
rect 57202 30270 57204 30322
rect 57148 30212 57204 30270
rect 57372 30212 57428 35086
rect 58156 35138 58212 36428
rect 59836 36482 59892 36494
rect 59836 36430 59838 36482
rect 59890 36430 59892 36482
rect 59836 36260 59892 36430
rect 61292 36482 61348 36494
rect 61292 36430 61294 36482
rect 61346 36430 61348 36482
rect 59836 36194 59892 36204
rect 60060 36372 60116 36382
rect 59172 36092 59436 36102
rect 59228 36036 59276 36092
rect 59332 36036 59380 36092
rect 59172 36026 59436 36036
rect 60060 35922 60116 36316
rect 60060 35870 60062 35922
rect 60114 35870 60116 35922
rect 60060 35858 60116 35870
rect 60508 36260 60564 36270
rect 60508 35924 60564 36204
rect 60508 35868 60900 35924
rect 59164 35700 59220 35710
rect 60732 35700 60788 35710
rect 59164 35698 60228 35700
rect 59164 35646 59166 35698
rect 59218 35646 60228 35698
rect 59164 35644 60228 35646
rect 59164 35634 59220 35644
rect 58940 35588 58996 35598
rect 58940 35494 58996 35532
rect 58156 35086 58158 35138
rect 58210 35086 58212 35138
rect 58156 35026 58212 35086
rect 58156 34974 58158 35026
rect 58210 34974 58212 35026
rect 58156 34962 58212 34974
rect 58268 35476 58324 35486
rect 57708 34916 57764 34926
rect 57596 34804 57652 34814
rect 57596 34690 57652 34748
rect 57596 34638 57598 34690
rect 57650 34638 57652 34690
rect 57484 34020 57540 34030
rect 57484 33926 57540 33964
rect 57596 33796 57652 34638
rect 57708 34132 57764 34860
rect 58268 34354 58324 35420
rect 59388 35474 59444 35486
rect 59388 35422 59390 35474
rect 59442 35422 59444 35474
rect 59164 35252 59220 35262
rect 59164 35138 59220 35196
rect 59164 35086 59166 35138
rect 59218 35086 59220 35138
rect 59164 35074 59220 35086
rect 59052 34916 59108 34926
rect 59052 34822 59108 34860
rect 59388 34692 59444 35422
rect 59612 35476 59668 35486
rect 59612 35382 59668 35420
rect 59388 34626 59444 34636
rect 59724 34914 59780 34926
rect 59724 34862 59726 34914
rect 59778 34862 59780 34914
rect 59172 34524 59436 34534
rect 59228 34468 59276 34524
rect 59332 34468 59380 34524
rect 59172 34458 59436 34468
rect 58268 34302 58270 34354
rect 58322 34302 58324 34354
rect 58268 34290 58324 34302
rect 59724 34354 59780 34862
rect 59724 34302 59726 34354
rect 59778 34302 59780 34354
rect 59724 34290 59780 34302
rect 57932 34244 57988 34254
rect 57708 34130 57876 34132
rect 57708 34078 57710 34130
rect 57762 34078 57876 34130
rect 57708 34076 57876 34078
rect 57708 34066 57764 34076
rect 57596 33730 57652 33740
rect 57820 33908 57876 34076
rect 57932 34130 57988 34188
rect 59388 34244 59444 34254
rect 59388 34150 59444 34188
rect 59500 34242 59556 34254
rect 59500 34190 59502 34242
rect 59554 34190 59556 34242
rect 58156 34132 58212 34142
rect 57932 34078 57934 34130
rect 57986 34078 57988 34130
rect 57932 34066 57988 34078
rect 58044 34130 58212 34132
rect 58044 34078 58158 34130
rect 58210 34078 58212 34130
rect 58044 34076 58212 34078
rect 57484 33348 57540 33358
rect 57484 32674 57540 33292
rect 57708 33348 57764 33358
rect 57708 33254 57764 33292
rect 57820 33346 57876 33852
rect 57820 33294 57822 33346
rect 57874 33294 57876 33346
rect 57820 33282 57876 33294
rect 57484 32622 57486 32674
rect 57538 32622 57540 32674
rect 57484 32610 57540 32622
rect 57596 33122 57652 33134
rect 57596 33070 57598 33122
rect 57650 33070 57652 33122
rect 57596 32004 57652 33070
rect 57932 32788 57988 32798
rect 58044 32788 58100 34076
rect 58156 34066 58212 34076
rect 58380 34130 58436 34142
rect 58380 34078 58382 34130
rect 58434 34078 58436 34130
rect 57932 32786 58100 32788
rect 57932 32734 57934 32786
rect 57986 32734 58100 32786
rect 57932 32732 58100 32734
rect 58380 32788 58436 34078
rect 59164 33124 59220 33134
rect 58828 33122 59220 33124
rect 58828 33070 59166 33122
rect 59218 33070 59220 33122
rect 58828 33068 59220 33070
rect 58492 32788 58548 32798
rect 58380 32786 58548 32788
rect 58380 32734 58494 32786
rect 58546 32734 58548 32786
rect 58380 32732 58548 32734
rect 57932 32722 57988 32732
rect 58492 32722 58548 32732
rect 58156 32676 58212 32686
rect 58716 32676 58772 32686
rect 57596 31938 57652 31948
rect 57708 32562 57764 32574
rect 57708 32510 57710 32562
rect 57762 32510 57764 32562
rect 57708 31554 57764 32510
rect 58156 32562 58212 32620
rect 58156 32510 58158 32562
rect 58210 32510 58212 32562
rect 58156 32498 58212 32510
rect 58604 32674 58772 32676
rect 58604 32622 58718 32674
rect 58770 32622 58772 32674
rect 58604 32620 58772 32622
rect 58604 31948 58660 32620
rect 58716 32610 58772 32620
rect 58828 32674 58884 33068
rect 59164 33058 59220 33068
rect 59172 32956 59436 32966
rect 59228 32900 59276 32956
rect 59332 32900 59380 32956
rect 59172 32890 59436 32900
rect 58828 32622 58830 32674
rect 58882 32622 58884 32674
rect 58828 31948 58884 32622
rect 59276 32676 59332 32686
rect 59276 32582 59332 32620
rect 59164 32004 59220 32042
rect 58604 31892 58772 31948
rect 58828 31892 58996 31948
rect 59164 31938 59220 31948
rect 59500 32004 59556 34190
rect 60172 34242 60228 35644
rect 60508 35586 60564 35598
rect 60508 35534 60510 35586
rect 60562 35534 60564 35586
rect 60508 35476 60564 35534
rect 60284 35420 60564 35476
rect 60620 35474 60676 35486
rect 60620 35422 60622 35474
rect 60674 35422 60676 35474
rect 60284 35252 60340 35420
rect 60620 35364 60676 35422
rect 60284 35186 60340 35196
rect 60396 35308 60620 35364
rect 60172 34190 60174 34242
rect 60226 34190 60228 34242
rect 60172 34178 60228 34190
rect 60284 34132 60340 34142
rect 60396 34132 60452 35308
rect 60620 35232 60676 35308
rect 60732 34692 60788 35644
rect 60620 34636 60788 34692
rect 60284 34130 60452 34132
rect 60284 34078 60286 34130
rect 60338 34078 60452 34130
rect 60284 34076 60452 34078
rect 60508 34132 60564 34142
rect 60284 34066 60340 34076
rect 60508 34038 60564 34076
rect 60620 34130 60676 34636
rect 60620 34078 60622 34130
rect 60674 34078 60676 34130
rect 60620 34066 60676 34078
rect 60732 34468 60788 34478
rect 60508 33234 60564 33246
rect 60508 33182 60510 33234
rect 60562 33182 60564 33234
rect 59500 31938 59556 31948
rect 59836 32676 59892 32686
rect 58492 31780 58548 31790
rect 57708 31502 57710 31554
rect 57762 31502 57764 31554
rect 57708 31444 57764 31502
rect 58268 31556 58324 31566
rect 58268 31462 58324 31500
rect 57708 31378 57764 31388
rect 58492 31218 58548 31724
rect 58716 31556 58772 31892
rect 58716 31490 58772 31500
rect 58492 31166 58494 31218
rect 58546 31166 58548 31218
rect 58492 31154 58548 31166
rect 58604 31106 58660 31118
rect 58604 31054 58606 31106
rect 58658 31054 58660 31106
rect 58604 30996 58660 31054
rect 57484 30940 58660 30996
rect 57484 30434 57540 30940
rect 57484 30382 57486 30434
rect 57538 30382 57540 30434
rect 57484 30370 57540 30382
rect 58380 30770 58436 30782
rect 58380 30718 58382 30770
rect 58434 30718 58436 30770
rect 58380 30322 58436 30718
rect 58380 30270 58382 30322
rect 58434 30270 58436 30322
rect 58380 30258 58436 30270
rect 57148 30146 57204 30156
rect 57260 30156 57428 30212
rect 58492 30212 58548 30222
rect 58492 30210 58660 30212
rect 58492 30158 58494 30210
rect 58546 30158 58660 30210
rect 58492 30156 58660 30158
rect 56700 29988 56756 29998
rect 56588 29316 56644 29326
rect 56588 29222 56644 29260
rect 56700 28644 56756 29932
rect 56700 28578 56756 28588
rect 56812 29428 56868 29438
rect 56812 28082 56868 29372
rect 56812 28030 56814 28082
rect 56866 28030 56868 28082
rect 56812 28018 56868 28030
rect 56588 27972 56644 27982
rect 56588 27878 56644 27916
rect 57036 27972 57092 27982
rect 56476 27858 56532 27870
rect 56476 27806 56478 27858
rect 56530 27806 56532 27858
rect 56476 27748 56532 27806
rect 56476 27692 56756 27748
rect 56476 27300 56532 27310
rect 56476 27206 56532 27244
rect 56252 27132 56420 27188
rect 56252 26178 56308 27132
rect 56252 26126 56254 26178
rect 56306 26126 56308 26178
rect 56252 25396 56308 26126
rect 56364 26962 56420 26974
rect 56364 26910 56366 26962
rect 56418 26910 56420 26962
rect 56364 25732 56420 26910
rect 56364 25666 56420 25676
rect 56700 26852 56756 27692
rect 57036 27300 57092 27916
rect 57260 27300 57316 30156
rect 58492 30146 58548 30156
rect 58156 30098 58212 30110
rect 58156 30046 58158 30098
rect 58210 30046 58212 30098
rect 57372 29986 57428 29998
rect 57372 29934 57374 29986
rect 57426 29934 57428 29986
rect 57372 29428 57428 29934
rect 57372 29362 57428 29372
rect 58044 29876 58100 29886
rect 58044 28532 58100 29820
rect 58156 29316 58212 30046
rect 58604 29428 58660 30156
rect 58940 30100 58996 31892
rect 59500 31780 59556 31790
rect 59500 31686 59556 31724
rect 59724 31668 59780 31678
rect 59724 31574 59780 31612
rect 59172 31388 59436 31398
rect 59228 31332 59276 31388
rect 59332 31332 59380 31388
rect 59172 31322 59436 31332
rect 59724 30882 59780 30894
rect 59724 30830 59726 30882
rect 59778 30830 59780 30882
rect 59724 30660 59780 30830
rect 59724 30594 59780 30604
rect 58940 30034 58996 30044
rect 59172 29820 59436 29830
rect 59228 29764 59276 29820
rect 59332 29764 59380 29820
rect 59172 29754 59436 29764
rect 59836 29652 59892 32620
rect 60284 32674 60340 32686
rect 60284 32622 60286 32674
rect 60338 32622 60340 32674
rect 60060 32564 60116 32574
rect 60060 32470 60116 32508
rect 60284 32004 60340 32622
rect 60284 31938 60340 31948
rect 60396 32562 60452 32574
rect 60396 32510 60398 32562
rect 60450 32510 60452 32562
rect 60396 32002 60452 32510
rect 60508 32564 60564 33182
rect 60620 33124 60676 33134
rect 60620 33030 60676 33068
rect 60508 32498 60564 32508
rect 60396 31950 60398 32002
rect 60450 31950 60452 32002
rect 60396 31938 60452 31950
rect 60284 31780 60340 31790
rect 60284 31686 60340 31724
rect 60396 31668 60452 31678
rect 60396 31574 60452 31612
rect 60732 31106 60788 34412
rect 60844 31948 60900 35868
rect 61292 34690 61348 36430
rect 62860 36372 62916 36382
rect 62860 36278 62916 36316
rect 63196 36372 63252 37548
rect 63308 36596 63364 39200
rect 65772 39060 65828 39200
rect 66108 39060 66164 39228
rect 65772 39004 66164 39060
rect 63308 36530 63364 36540
rect 64652 36596 64708 36606
rect 64652 36502 64708 36540
rect 66444 36594 66500 39228
rect 68208 39200 68320 40000
rect 70672 39200 70784 40000
rect 73136 39200 73248 40000
rect 75600 39200 75712 40000
rect 75964 39228 77028 39284
rect 68236 38164 68292 39200
rect 68236 38108 68628 38164
rect 68460 37940 68516 37950
rect 66444 36542 66446 36594
rect 66498 36542 66500 36594
rect 66444 36530 66500 36542
rect 67452 37156 67508 37166
rect 65772 36484 65828 36494
rect 65772 36482 65940 36484
rect 65772 36430 65774 36482
rect 65826 36430 65940 36482
rect 65772 36428 65940 36430
rect 65772 36418 65828 36428
rect 63196 36240 63252 36316
rect 63868 36260 63924 36270
rect 65884 36260 65940 36428
rect 63868 36258 64484 36260
rect 63868 36206 63870 36258
rect 63922 36206 64484 36258
rect 63868 36204 64484 36206
rect 63868 36194 63924 36204
rect 62972 35810 63028 35822
rect 62972 35758 62974 35810
rect 63026 35758 63028 35810
rect 61404 35700 61460 35710
rect 61404 35606 61460 35644
rect 61852 35698 61908 35710
rect 61852 35646 61854 35698
rect 61906 35646 61908 35698
rect 61852 35588 61908 35646
rect 61852 35522 61908 35532
rect 62300 35586 62356 35598
rect 62300 35534 62302 35586
rect 62354 35534 62356 35586
rect 62300 35252 62356 35534
rect 62860 35588 62916 35598
rect 62860 35494 62916 35532
rect 62300 35186 62356 35196
rect 62524 35364 62580 35374
rect 62524 34914 62580 35308
rect 62972 35364 63028 35758
rect 64204 35698 64260 35710
rect 64204 35646 64206 35698
rect 64258 35646 64260 35698
rect 63196 35476 63252 35486
rect 62972 35298 63028 35308
rect 63084 35474 63252 35476
rect 63084 35422 63198 35474
rect 63250 35422 63252 35474
rect 63084 35420 63252 35422
rect 62524 34862 62526 34914
rect 62578 34862 62580 34914
rect 62524 34850 62580 34862
rect 62748 35026 62804 35038
rect 62748 34974 62750 35026
rect 62802 34974 62804 35026
rect 61292 34638 61294 34690
rect 61346 34638 61348 34690
rect 61292 34468 61348 34638
rect 61292 34402 61348 34412
rect 62748 34354 62804 34974
rect 62748 34302 62750 34354
rect 62802 34302 62804 34354
rect 62748 34290 62804 34302
rect 61516 34244 61572 34254
rect 61516 33570 61572 34188
rect 62972 34242 63028 34254
rect 62972 34190 62974 34242
rect 63026 34190 63028 34242
rect 61516 33518 61518 33570
rect 61570 33518 61572 33570
rect 61516 33506 61572 33518
rect 62524 33796 62580 33806
rect 61628 33236 61684 33246
rect 62524 33236 62580 33740
rect 62972 33572 63028 34190
rect 63084 34132 63140 35420
rect 63196 35410 63252 35420
rect 64204 34916 64260 35646
rect 64204 34850 64260 34860
rect 64428 35698 64484 36204
rect 64428 35646 64430 35698
rect 64482 35646 64484 35698
rect 63196 34804 63252 34814
rect 63196 34710 63252 34748
rect 63980 34804 64036 34814
rect 63980 34710 64036 34748
rect 64428 34804 64484 35646
rect 64764 35700 64820 35710
rect 64764 35606 64820 35644
rect 65548 35700 65604 35710
rect 64540 35588 64596 35598
rect 64540 35494 64596 35532
rect 64988 35252 65044 35262
rect 64988 35138 65044 35196
rect 64988 35086 64990 35138
rect 65042 35086 65044 35138
rect 64988 35074 65044 35086
rect 64428 34738 64484 34748
rect 64988 34916 65044 34926
rect 64092 34692 64148 34702
rect 64092 34598 64148 34636
rect 64764 34690 64820 34702
rect 64764 34638 64766 34690
rect 64818 34638 64820 34690
rect 64764 34580 64820 34638
rect 64764 34514 64820 34524
rect 64092 34356 64148 34366
rect 63084 34038 63140 34076
rect 63868 34244 63924 34254
rect 63196 33572 63252 33582
rect 62972 33570 63252 33572
rect 62972 33518 63198 33570
rect 63250 33518 63252 33570
rect 62972 33516 63252 33518
rect 63084 33236 63140 33246
rect 61628 33234 61796 33236
rect 61628 33182 61630 33234
rect 61682 33182 61796 33234
rect 61628 33180 61796 33182
rect 61628 33170 61684 33180
rect 61516 33124 61572 33134
rect 61516 33030 61572 33068
rect 61740 32788 61796 33180
rect 62524 33234 63140 33236
rect 62524 33182 62526 33234
rect 62578 33182 63086 33234
rect 63138 33182 63140 33234
rect 62524 33180 63140 33182
rect 62524 33170 62580 33180
rect 61404 32732 61796 32788
rect 63084 32788 63140 33180
rect 63196 33236 63252 33516
rect 63868 33460 63924 34188
rect 63868 33394 63924 33404
rect 64092 33460 64148 34300
rect 64988 34356 65044 34860
rect 65324 34916 65380 34926
rect 65324 34822 65380 34860
rect 65548 34914 65604 35644
rect 65660 35698 65716 35710
rect 65660 35646 65662 35698
rect 65714 35646 65716 35698
rect 65660 35252 65716 35646
rect 65772 35588 65828 35598
rect 65772 35494 65828 35532
rect 65660 35186 65716 35196
rect 65548 34862 65550 34914
rect 65602 34862 65604 34914
rect 65548 34850 65604 34862
rect 64988 34290 65044 34300
rect 65660 34692 65716 34702
rect 65660 34242 65716 34636
rect 65772 34356 65828 34366
rect 65772 34262 65828 34300
rect 65660 34190 65662 34242
rect 65714 34190 65716 34242
rect 65660 34178 65716 34190
rect 65100 34132 65156 34142
rect 65100 33570 65156 34076
rect 65100 33518 65102 33570
rect 65154 33518 65156 33570
rect 65100 33506 65156 33518
rect 64092 33394 64148 33404
rect 64204 33348 64260 33358
rect 64204 33254 64260 33292
rect 65436 33348 65492 33358
rect 65436 33254 65492 33292
rect 63196 33170 63252 33180
rect 63868 33234 63924 33246
rect 63868 33182 63870 33234
rect 63922 33182 63924 33234
rect 63532 32788 63588 32798
rect 63084 32786 63588 32788
rect 63084 32734 63534 32786
rect 63586 32734 63588 32786
rect 63084 32732 63588 32734
rect 60844 31892 61124 31948
rect 61068 31220 61124 31892
rect 60732 31054 60734 31106
rect 60786 31054 60788 31106
rect 60172 30882 60228 30894
rect 60172 30830 60174 30882
rect 60226 30830 60228 30882
rect 60172 30660 60228 30830
rect 60172 30594 60228 30604
rect 60732 30548 60788 31054
rect 60732 30482 60788 30492
rect 60956 31164 61124 31220
rect 60844 30100 60900 30110
rect 59724 29538 59780 29550
rect 59724 29486 59726 29538
rect 59778 29486 59780 29538
rect 58604 29334 58660 29372
rect 59500 29428 59556 29438
rect 59500 29334 59556 29372
rect 58156 29222 58212 29260
rect 59724 29316 59780 29486
rect 59836 29538 59892 29596
rect 59836 29486 59838 29538
rect 59890 29486 59892 29538
rect 59836 29474 59892 29486
rect 60620 29986 60676 29998
rect 60620 29934 60622 29986
rect 60674 29934 60676 29986
rect 60620 29540 60676 29934
rect 60620 29474 60676 29484
rect 60732 29652 60788 29662
rect 59724 29250 59780 29260
rect 60284 29316 60340 29326
rect 58940 29202 58996 29214
rect 58940 29150 58942 29202
rect 58994 29150 58996 29202
rect 58268 28644 58324 28654
rect 58156 28532 58212 28542
rect 58044 28530 58212 28532
rect 58044 28478 58158 28530
rect 58210 28478 58212 28530
rect 58044 28476 58212 28478
rect 57036 27186 57092 27244
rect 57036 27134 57038 27186
rect 57090 27134 57092 27186
rect 57036 27122 57092 27134
rect 57148 27244 57316 27300
rect 57372 27860 57428 27870
rect 57372 27746 57428 27804
rect 57372 27694 57374 27746
rect 57426 27694 57428 27746
rect 57372 27300 57428 27694
rect 58044 27748 58100 28476
rect 58156 28466 58212 28476
rect 58268 28418 58324 28588
rect 58828 28642 58884 28654
rect 58828 28590 58830 28642
rect 58882 28590 58884 28642
rect 58268 28366 58270 28418
rect 58322 28366 58324 28418
rect 58268 27860 58324 28366
rect 58268 27794 58324 27804
rect 58492 28418 58548 28430
rect 58492 28366 58494 28418
rect 58546 28366 58548 28418
rect 58492 27860 58548 28366
rect 58828 27860 58884 28590
rect 58940 28532 58996 29150
rect 58940 28466 58996 28476
rect 59724 28642 59780 28654
rect 59724 28590 59726 28642
rect 59778 28590 59780 28642
rect 59724 28532 59780 28590
rect 59724 28466 59780 28476
rect 60172 28642 60228 28654
rect 60172 28590 60174 28642
rect 60226 28590 60228 28642
rect 59500 28420 59556 28430
rect 59172 28252 59436 28262
rect 59228 28196 59276 28252
rect 59332 28196 59380 28252
rect 59172 28186 59436 28196
rect 59276 27972 59332 27982
rect 59276 27878 59332 27916
rect 58492 27858 58660 27860
rect 58492 27806 58494 27858
rect 58546 27806 58660 27858
rect 58492 27804 58660 27806
rect 58492 27794 58548 27804
rect 58044 27682 58100 27692
rect 58156 27634 58212 27646
rect 58156 27582 58158 27634
rect 58210 27582 58212 27634
rect 56700 26178 56756 26796
rect 56700 26126 56702 26178
rect 56754 26126 56756 26178
rect 56476 25396 56532 25406
rect 56252 25340 56476 25396
rect 56476 25282 56532 25340
rect 56476 25230 56478 25282
rect 56530 25230 56532 25282
rect 56140 23492 56196 23502
rect 56140 23154 56196 23436
rect 56140 23102 56142 23154
rect 56194 23102 56196 23154
rect 56140 23090 56196 23102
rect 56028 22764 56420 22820
rect 55916 22708 55972 22718
rect 54908 22484 54964 22494
rect 54348 22482 54964 22484
rect 54348 22430 54350 22482
rect 54402 22430 54910 22482
rect 54962 22430 54964 22482
rect 54348 22428 54964 22430
rect 52668 22318 52670 22370
rect 52722 22318 52724 22370
rect 52668 22306 52724 22318
rect 53900 22370 53956 22382
rect 53900 22318 53902 22370
rect 53954 22318 53956 22370
rect 53452 22260 53508 22270
rect 53452 22166 53508 22204
rect 52500 22092 52612 22148
rect 52444 22082 52500 22092
rect 52332 21634 52388 21644
rect 52444 21924 52500 21934
rect 52332 20692 52388 20702
rect 52220 20690 52388 20692
rect 52220 20638 52334 20690
rect 52386 20638 52388 20690
rect 52220 20636 52388 20638
rect 52332 20626 52388 20636
rect 52332 19796 52388 19806
rect 52332 19346 52388 19740
rect 52332 19294 52334 19346
rect 52386 19294 52388 19346
rect 52332 18676 52388 19294
rect 52332 18610 52388 18620
rect 52444 18788 52500 21868
rect 53564 21700 53620 21710
rect 53900 21700 53956 22318
rect 53564 21698 53956 21700
rect 53564 21646 53566 21698
rect 53618 21646 53956 21698
rect 53564 21644 53956 21646
rect 54236 21812 54292 21822
rect 54348 21812 54404 22428
rect 54908 22418 54964 22428
rect 55916 22482 55972 22652
rect 55916 22430 55918 22482
rect 55970 22430 55972 22482
rect 55916 22418 55972 22430
rect 55468 22148 55524 22158
rect 55468 22054 55524 22092
rect 54236 21810 54404 21812
rect 54236 21758 54238 21810
rect 54290 21758 54404 21810
rect 54236 21756 54404 21758
rect 56364 21810 56420 22764
rect 56476 22708 56532 25230
rect 56700 23492 56756 26126
rect 57148 25956 57204 27244
rect 57372 27234 57428 27244
rect 57596 27300 57652 27310
rect 58156 27300 58212 27582
rect 58492 27636 58548 27646
rect 58492 27542 58548 27580
rect 57596 27298 58324 27300
rect 57596 27246 57598 27298
rect 57650 27246 58324 27298
rect 57596 27244 58324 27246
rect 57596 27234 57652 27244
rect 58268 27186 58324 27244
rect 58268 27134 58270 27186
rect 58322 27134 58324 27186
rect 58268 27122 58324 27134
rect 57260 27074 57316 27086
rect 57260 27022 57262 27074
rect 57314 27022 57316 27074
rect 57260 26908 57316 27022
rect 57708 27076 57764 27086
rect 57260 26852 57652 26908
rect 57484 26290 57540 26302
rect 57484 26238 57486 26290
rect 57538 26238 57540 26290
rect 57148 25900 57428 25956
rect 57148 25732 57204 25742
rect 57148 25638 57204 25676
rect 57148 25508 57204 25518
rect 57036 25396 57092 25406
rect 57036 25302 57092 25340
rect 57148 25394 57204 25452
rect 57148 25342 57150 25394
rect 57202 25342 57204 25394
rect 57148 25330 57204 25342
rect 56700 23426 56756 23436
rect 56812 23940 56868 23950
rect 56700 23156 56756 23166
rect 56700 23062 56756 23100
rect 56476 22642 56532 22652
rect 56812 22484 56868 23884
rect 56924 22484 56980 22494
rect 57372 22484 57428 25900
rect 57484 25396 57540 26238
rect 57596 26178 57652 26852
rect 57708 26292 57764 27020
rect 58604 27074 58660 27804
rect 58828 27794 58884 27804
rect 59388 27748 59444 27758
rect 59500 27748 59556 28364
rect 60172 28420 60228 28590
rect 60172 28354 60228 28364
rect 60284 27972 60340 29260
rect 60284 27906 60340 27916
rect 60620 28530 60676 28542
rect 60620 28478 60622 28530
rect 60674 28478 60676 28530
rect 60620 27972 60676 28478
rect 60620 27906 60676 27916
rect 59388 27746 59556 27748
rect 59388 27694 59390 27746
rect 59442 27694 59556 27746
rect 59388 27692 59556 27694
rect 59724 27860 59780 27870
rect 59388 27682 59444 27692
rect 59052 27636 59108 27646
rect 59052 27542 59108 27580
rect 58604 27022 58606 27074
rect 58658 27022 58660 27074
rect 58604 27010 58660 27022
rect 59164 26964 59220 26974
rect 59164 26870 59220 26908
rect 57932 26852 57988 26862
rect 57932 26514 57988 26796
rect 59500 26852 59556 26862
rect 59172 26684 59436 26694
rect 59228 26628 59276 26684
rect 59332 26628 59380 26684
rect 59172 26618 59436 26628
rect 57932 26462 57934 26514
rect 57986 26462 57988 26514
rect 57932 26450 57988 26462
rect 57708 26198 57764 26236
rect 58156 26290 58212 26302
rect 58156 26238 58158 26290
rect 58210 26238 58212 26290
rect 57596 26126 57598 26178
rect 57650 26126 57652 26178
rect 57596 26114 57652 26126
rect 58156 26180 58212 26238
rect 59052 26292 59108 26302
rect 58604 26180 58660 26190
rect 58156 26178 58660 26180
rect 58156 26126 58606 26178
rect 58658 26126 58660 26178
rect 58156 26124 58660 26126
rect 57484 25330 57540 25340
rect 57708 25732 57764 25742
rect 57708 24722 57764 25676
rect 58380 25620 58436 25630
rect 58380 25526 58436 25564
rect 57708 24670 57710 24722
rect 57762 24670 57764 24722
rect 57708 24658 57764 24670
rect 57820 25506 57876 25518
rect 58044 25508 58100 25518
rect 57820 25454 57822 25506
rect 57874 25454 57876 25506
rect 57596 23940 57652 23950
rect 57596 23378 57652 23884
rect 57596 23326 57598 23378
rect 57650 23326 57652 23378
rect 57596 23314 57652 23326
rect 57820 23938 57876 25454
rect 57932 25506 58100 25508
rect 57932 25454 58046 25506
rect 58098 25454 58100 25506
rect 57932 25452 58100 25454
rect 57932 24498 57988 25452
rect 58044 25442 58100 25452
rect 58604 25508 58660 26124
rect 59052 26180 59108 26236
rect 59052 26178 59220 26180
rect 59052 26126 59054 26178
rect 59106 26126 59220 26178
rect 59052 26124 59220 26126
rect 59052 26114 59108 26124
rect 58604 25442 58660 25452
rect 59052 25508 59108 25518
rect 59052 25414 59108 25452
rect 58940 25396 58996 25406
rect 58268 25282 58324 25294
rect 58268 25230 58270 25282
rect 58322 25230 58324 25282
rect 57932 24446 57934 24498
rect 57986 24446 57988 24498
rect 57932 24050 57988 24446
rect 57932 23998 57934 24050
rect 57986 23998 57988 24050
rect 57932 23986 57988 23998
rect 58044 24722 58100 24734
rect 58044 24670 58046 24722
rect 58098 24670 58100 24722
rect 57820 23886 57822 23938
rect 57874 23886 57876 23938
rect 57484 23156 57540 23166
rect 57484 23062 57540 23100
rect 57596 22932 57652 22942
rect 57596 22838 57652 22876
rect 56812 22482 57204 22484
rect 56812 22430 56926 22482
rect 56978 22430 57204 22482
rect 56812 22428 57204 22430
rect 57372 22428 57764 22484
rect 56924 22418 56980 22428
rect 56476 22148 56532 22158
rect 56476 22054 56532 22092
rect 56364 21758 56366 21810
rect 56418 21758 56420 21810
rect 52668 20692 52724 20702
rect 53452 20692 53508 20702
rect 52668 20690 53508 20692
rect 52668 20638 52670 20690
rect 52722 20638 53454 20690
rect 53506 20638 53508 20690
rect 52668 20636 53508 20638
rect 52668 20626 52724 20636
rect 53452 20626 53508 20636
rect 53564 20580 53620 21644
rect 53564 20514 53620 20524
rect 53676 21474 53732 21486
rect 53676 21422 53678 21474
rect 53730 21422 53732 21474
rect 53676 20132 53732 21422
rect 53788 21476 53844 21486
rect 53788 21382 53844 21420
rect 54236 21476 54292 21756
rect 56364 21746 56420 21758
rect 55916 21588 55972 21598
rect 55916 21494 55972 21532
rect 54236 21410 54292 21420
rect 55020 21476 55076 21486
rect 55020 21028 55076 21420
rect 55020 20914 55076 20972
rect 55020 20862 55022 20914
rect 55074 20862 55076 20914
rect 55020 20850 55076 20862
rect 55468 21474 55524 21486
rect 55468 21422 55470 21474
rect 55522 21422 55524 21474
rect 54124 20802 54180 20814
rect 54124 20750 54126 20802
rect 54178 20750 54180 20802
rect 54124 20244 54180 20750
rect 54348 20804 54404 20814
rect 54348 20710 54404 20748
rect 54348 20580 54404 20590
rect 54236 20244 54292 20254
rect 54124 20242 54292 20244
rect 54124 20190 54238 20242
rect 54290 20190 54292 20242
rect 54124 20188 54292 20190
rect 54236 20178 54292 20188
rect 53676 20076 54180 20132
rect 53564 20020 53620 20030
rect 53564 19926 53620 19964
rect 54124 20018 54180 20076
rect 54124 19966 54126 20018
rect 54178 19966 54180 20018
rect 54124 19954 54180 19966
rect 53004 19908 53060 19918
rect 53004 19906 53172 19908
rect 53004 19854 53006 19906
rect 53058 19854 53172 19906
rect 53004 19852 53172 19854
rect 53004 19842 53060 19852
rect 53116 19348 53172 19852
rect 53228 19794 53284 19806
rect 53228 19742 53230 19794
rect 53282 19742 53284 19794
rect 53228 19572 53284 19742
rect 53228 19506 53284 19516
rect 53788 19460 53844 19470
rect 53116 19292 53732 19348
rect 52332 18452 52388 18462
rect 52444 18452 52500 18732
rect 53228 18562 53284 19292
rect 53676 19234 53732 19292
rect 53788 19346 53844 19404
rect 54348 19458 54404 20524
rect 55468 20580 55524 21422
rect 55692 21364 55748 21374
rect 55468 20514 55524 20524
rect 55580 21362 55748 21364
rect 55580 21310 55694 21362
rect 55746 21310 55748 21362
rect 55580 21308 55748 21310
rect 55580 20804 55636 21308
rect 55692 21298 55748 21308
rect 55804 21028 55860 21038
rect 55804 20934 55860 20972
rect 56140 20916 56196 20954
rect 56140 20850 56196 20860
rect 54460 20020 54516 20030
rect 54460 19926 54516 19964
rect 54348 19406 54350 19458
rect 54402 19406 54404 19458
rect 54348 19394 54404 19406
rect 53788 19294 53790 19346
rect 53842 19294 53844 19346
rect 53788 19282 53844 19294
rect 53676 19182 53678 19234
rect 53730 19182 53732 19234
rect 53676 19170 53732 19182
rect 55580 19236 55636 20748
rect 55916 20692 55972 20702
rect 55916 20242 55972 20636
rect 56140 20690 56196 20702
rect 56140 20638 56142 20690
rect 56194 20638 56196 20690
rect 56140 20580 56196 20638
rect 56364 20692 56420 20702
rect 56364 20598 56420 20636
rect 56140 20514 56196 20524
rect 55916 20190 55918 20242
rect 55970 20190 55972 20242
rect 55916 20178 55972 20190
rect 55804 20020 55860 20030
rect 55804 19926 55860 19964
rect 56028 20018 56084 20030
rect 56028 19966 56030 20018
rect 56082 19966 56084 20018
rect 55804 19236 55860 19246
rect 55580 19234 55860 19236
rect 55580 19182 55806 19234
rect 55858 19182 55860 19234
rect 55580 19180 55860 19182
rect 56028 19236 56084 19966
rect 56476 20020 56532 20030
rect 56476 20018 56644 20020
rect 56476 19966 56478 20018
rect 56530 19966 56644 20018
rect 56476 19964 56644 19966
rect 56476 19954 56532 19964
rect 56588 19348 56644 19964
rect 56588 19254 56644 19292
rect 56252 19236 56308 19246
rect 56028 19234 56308 19236
rect 56028 19182 56254 19234
rect 56306 19182 56308 19234
rect 56028 19180 56308 19182
rect 55804 19170 55860 19180
rect 55356 18676 55412 18686
rect 55356 18582 55412 18620
rect 56252 18676 56308 19180
rect 56252 18610 56308 18620
rect 53228 18510 53230 18562
rect 53282 18510 53284 18562
rect 53228 18498 53284 18510
rect 52332 18450 52500 18452
rect 52332 18398 52334 18450
rect 52386 18398 52500 18450
rect 52332 18396 52500 18398
rect 53788 18452 53844 18462
rect 52332 18386 52388 18396
rect 53788 18358 53844 18396
rect 54796 18452 54852 18462
rect 54796 18358 54852 18396
rect 54124 18340 54180 18350
rect 54124 18246 54180 18284
rect 55020 18340 55076 18350
rect 55020 18246 55076 18284
rect 55468 18340 55524 18350
rect 53340 17780 53396 17790
rect 53340 17686 53396 17724
rect 52444 17556 52500 17566
rect 53676 17556 53732 17566
rect 52444 17554 52836 17556
rect 52444 17502 52446 17554
rect 52498 17502 52836 17554
rect 52444 17500 52836 17502
rect 52444 17490 52500 17500
rect 52220 17444 52276 17454
rect 52220 17350 52276 17388
rect 52332 17442 52388 17454
rect 52332 17390 52334 17442
rect 52386 17390 52388 17442
rect 52332 16324 52388 17390
rect 52780 17106 52836 17500
rect 52780 17054 52782 17106
rect 52834 17054 52836 17106
rect 52780 17042 52836 17054
rect 52892 17108 52948 17118
rect 52892 17014 52948 17052
rect 53676 17106 53732 17500
rect 53676 17054 53678 17106
rect 53730 17054 53732 17106
rect 53676 16884 53732 17054
rect 54460 17220 54516 17230
rect 53676 16818 53732 16828
rect 54236 16884 54292 16894
rect 54236 16790 54292 16828
rect 52668 16772 52724 16782
rect 52668 16678 52724 16716
rect 54460 16770 54516 17164
rect 54460 16718 54462 16770
rect 54514 16718 54516 16770
rect 54460 16706 54516 16718
rect 55020 17220 55076 17230
rect 55020 16996 55076 17164
rect 54796 16658 54852 16670
rect 54796 16606 54798 16658
rect 54850 16606 54852 16658
rect 52332 16258 52388 16268
rect 54236 16324 54292 16334
rect 53116 16100 53172 16110
rect 52780 15876 52836 15886
rect 52444 15316 52500 15326
rect 52444 14644 52500 15260
rect 52780 15314 52836 15820
rect 52780 15262 52782 15314
rect 52834 15262 52836 15314
rect 52780 15250 52836 15262
rect 53116 15316 53172 16044
rect 53116 15184 53172 15260
rect 54124 15316 54180 15326
rect 54124 15222 54180 15260
rect 52444 14578 52500 14588
rect 54012 15090 54068 15102
rect 54012 15038 54014 15090
rect 54066 15038 54068 15090
rect 53116 14532 53172 14542
rect 54012 14532 54068 15038
rect 54236 14532 54292 16268
rect 54572 16100 54628 16110
rect 54572 16006 54628 16044
rect 54796 15988 54852 16606
rect 55020 16210 55076 16940
rect 55468 16994 55524 18284
rect 55468 16942 55470 16994
rect 55522 16942 55524 16994
rect 55468 16930 55524 16942
rect 55020 16158 55022 16210
rect 55074 16158 55076 16210
rect 55020 16146 55076 16158
rect 55132 16884 55188 16894
rect 54796 15316 54852 15932
rect 54796 15250 54852 15260
rect 53116 13524 53172 14476
rect 53788 14530 54068 14532
rect 53788 14478 54014 14530
rect 54066 14478 54068 14530
rect 53788 14476 54068 14478
rect 53788 13858 53844 14476
rect 54012 14466 54068 14476
rect 54124 14530 54292 14532
rect 54124 14478 54238 14530
rect 54290 14478 54292 14530
rect 54124 14476 54292 14478
rect 53788 13806 53790 13858
rect 53842 13806 53844 13858
rect 53788 13794 53844 13806
rect 54012 13748 54068 13758
rect 54124 13748 54180 14476
rect 54236 14466 54292 14476
rect 54908 14532 54964 14542
rect 54964 14476 55076 14532
rect 54908 14438 54964 14476
rect 54012 13746 54180 13748
rect 54012 13694 54014 13746
rect 54066 13694 54180 13746
rect 54012 13692 54180 13694
rect 54460 14418 54516 14430
rect 54460 14366 54462 14418
rect 54514 14366 54516 14418
rect 54012 13682 54068 13692
rect 52668 12738 52724 12750
rect 52668 12686 52670 12738
rect 52722 12686 52724 12738
rect 52668 12516 52724 12686
rect 52668 12450 52724 12460
rect 53116 12402 53172 13468
rect 54012 13524 54068 13534
rect 53788 12964 53844 12974
rect 53116 12350 53118 12402
rect 53170 12350 53172 12402
rect 53116 12338 53172 12350
rect 53676 12740 53732 12750
rect 53564 12292 53620 12302
rect 53564 12198 53620 12236
rect 52332 11506 52388 11518
rect 52332 11454 52334 11506
rect 52386 11454 52388 11506
rect 52220 11172 52276 11182
rect 52332 11172 52388 11454
rect 53452 11284 53508 11294
rect 53004 11282 53508 11284
rect 53004 11230 53454 11282
rect 53506 11230 53508 11282
rect 53004 11228 53508 11230
rect 53004 11172 53060 11228
rect 53452 11218 53508 11228
rect 52332 11116 53060 11172
rect 52220 10836 52276 11116
rect 52780 10948 52836 10958
rect 52444 10836 52500 10846
rect 52220 10834 52500 10836
rect 52220 10782 52446 10834
rect 52498 10782 52500 10834
rect 52220 10780 52500 10782
rect 52444 10724 52500 10780
rect 52444 10658 52500 10668
rect 52108 9762 52164 9772
rect 52780 9716 52836 10892
rect 53004 10834 53060 11116
rect 53676 11060 53732 12684
rect 53788 12516 53844 12908
rect 53788 12450 53844 12460
rect 54012 12178 54068 13468
rect 54348 13524 54404 13534
rect 54348 13430 54404 13468
rect 54460 13300 54516 14366
rect 54348 13244 54460 13300
rect 54348 13074 54404 13244
rect 54460 13234 54516 13244
rect 54908 13746 54964 13758
rect 54908 13694 54910 13746
rect 54962 13694 54964 13746
rect 54348 13022 54350 13074
rect 54402 13022 54404 13074
rect 54348 13010 54404 13022
rect 54460 13074 54516 13086
rect 54460 13022 54462 13074
rect 54514 13022 54516 13074
rect 54012 12126 54014 12178
rect 54066 12126 54068 12178
rect 54012 12114 54068 12126
rect 54460 12292 54516 13022
rect 54460 12178 54516 12236
rect 54460 12126 54462 12178
rect 54514 12126 54516 12178
rect 54460 12114 54516 12126
rect 54908 12068 54964 13694
rect 55020 13748 55076 14476
rect 55132 13970 55188 16828
rect 55916 16884 55972 16894
rect 55916 16790 55972 16828
rect 56364 16772 56420 16782
rect 56364 16678 56420 16716
rect 56700 16772 56756 16782
rect 55916 16156 56644 16212
rect 55580 16100 55636 16110
rect 55580 16006 55636 16044
rect 55916 16098 55972 16156
rect 55916 16046 55918 16098
rect 55970 16046 55972 16098
rect 55916 16034 55972 16046
rect 56588 16098 56644 16156
rect 56588 16046 56590 16098
rect 56642 16046 56644 16098
rect 56588 16034 56644 16046
rect 56364 15988 56420 15998
rect 56364 15894 56420 15932
rect 55692 15876 55748 15886
rect 55692 15782 55748 15820
rect 56588 15874 56644 15886
rect 56588 15822 56590 15874
rect 56642 15822 56644 15874
rect 56588 15428 56644 15822
rect 56588 15362 56644 15372
rect 56700 14754 56756 16716
rect 56924 16100 56980 16110
rect 56924 16006 56980 16044
rect 56700 14702 56702 14754
rect 56754 14702 56756 14754
rect 56700 14690 56756 14702
rect 57148 14756 57204 22428
rect 57484 22260 57540 22270
rect 57484 22166 57540 22204
rect 57596 22146 57652 22158
rect 57596 22094 57598 22146
rect 57650 22094 57652 22146
rect 57596 21924 57652 22094
rect 57596 21858 57652 21868
rect 57708 21812 57764 22428
rect 57820 22370 57876 23886
rect 58044 22932 58100 24670
rect 58268 23716 58324 25230
rect 58492 25282 58548 25294
rect 58492 25230 58494 25282
rect 58546 25230 58548 25282
rect 58492 24948 58548 25230
rect 58492 24882 58548 24892
rect 58380 23940 58436 23950
rect 58380 23846 58436 23884
rect 58940 23938 58996 25340
rect 59164 25284 59220 26124
rect 59164 25218 59220 25228
rect 59500 25282 59556 26796
rect 59500 25230 59502 25282
rect 59554 25230 59556 25282
rect 59172 25116 59436 25126
rect 59228 25060 59276 25116
rect 59332 25060 59380 25116
rect 59172 25050 59436 25060
rect 59052 24948 59108 24958
rect 59052 24854 59108 24892
rect 59276 24836 59332 24846
rect 59276 24742 59332 24780
rect 59388 24836 59444 24846
rect 59500 24836 59556 25230
rect 59388 24834 59556 24836
rect 59388 24782 59390 24834
rect 59442 24782 59556 24834
rect 59388 24780 59556 24782
rect 59388 24770 59444 24780
rect 58940 23886 58942 23938
rect 58994 23886 58996 23938
rect 58940 23874 58996 23886
rect 59052 23828 59108 23838
rect 59724 23828 59780 27804
rect 60396 27860 60452 27870
rect 60396 27766 60452 27804
rect 59836 27748 59892 27758
rect 59836 27654 59892 27692
rect 60620 27634 60676 27646
rect 60620 27582 60622 27634
rect 60674 27582 60676 27634
rect 60060 26404 60116 26414
rect 60060 26310 60116 26348
rect 60620 26178 60676 27582
rect 60620 26126 60622 26178
rect 60674 26126 60676 26178
rect 59948 25508 60004 25518
rect 59948 25284 60004 25452
rect 60396 25396 60452 25406
rect 59948 25282 60116 25284
rect 59948 25230 59950 25282
rect 60002 25230 60116 25282
rect 59948 25228 60116 25230
rect 59948 25218 60004 25228
rect 60060 24836 60116 25228
rect 59052 23734 59108 23772
rect 58268 23650 58324 23660
rect 59276 23716 59332 23792
rect 59724 23734 59780 23772
rect 59948 24610 60004 24622
rect 59948 24558 59950 24610
rect 60002 24558 60004 24610
rect 59836 23716 59892 23726
rect 59332 23660 59556 23716
rect 59276 23650 59332 23660
rect 59172 23548 59436 23558
rect 59228 23492 59276 23548
rect 59332 23492 59380 23548
rect 59172 23482 59436 23492
rect 58044 22866 58100 22876
rect 58156 23156 58212 23166
rect 58156 23042 58212 23100
rect 58156 22990 58158 23042
rect 58210 22990 58212 23042
rect 57820 22318 57822 22370
rect 57874 22318 57876 22370
rect 57820 22306 57876 22318
rect 58156 21924 58212 22990
rect 58716 23042 58772 23054
rect 58716 22990 58718 23042
rect 58770 22990 58772 23042
rect 58380 22484 58436 22494
rect 57820 21812 57876 21822
rect 57708 21810 57876 21812
rect 57708 21758 57822 21810
rect 57874 21758 57876 21810
rect 57708 21756 57876 21758
rect 57820 21746 57876 21756
rect 58044 21588 58100 21598
rect 57932 21586 58100 21588
rect 57932 21534 58046 21586
rect 58098 21534 58100 21586
rect 57932 21532 58100 21534
rect 57932 20914 57988 21532
rect 58044 21522 58100 21532
rect 57932 20862 57934 20914
rect 57986 20862 57988 20914
rect 57932 20850 57988 20862
rect 58156 20692 58212 21868
rect 58268 22258 58324 22270
rect 58268 22206 58270 22258
rect 58322 22206 58324 22258
rect 58268 22148 58324 22206
rect 58268 21476 58324 22092
rect 58380 22146 58436 22428
rect 58604 22260 58660 22270
rect 58604 22166 58660 22204
rect 58380 22094 58382 22146
rect 58434 22094 58436 22146
rect 58380 22036 58436 22094
rect 58716 22148 58772 22990
rect 58940 23044 58996 23054
rect 58940 22950 58996 22988
rect 59500 23044 59556 23660
rect 59836 23622 59892 23660
rect 59948 23492 60004 24558
rect 60060 24612 60116 24780
rect 60284 24612 60340 24622
rect 60060 24610 60340 24612
rect 60060 24558 60286 24610
rect 60338 24558 60340 24610
rect 60060 24556 60340 24558
rect 59500 22978 59556 22988
rect 59724 23436 60004 23492
rect 60060 23714 60116 23726
rect 60060 23662 60062 23714
rect 60114 23662 60116 23714
rect 59276 22930 59332 22942
rect 59276 22878 59278 22930
rect 59330 22878 59332 22930
rect 59276 22596 59332 22878
rect 59500 22596 59556 22606
rect 59276 22594 59556 22596
rect 59276 22542 59502 22594
rect 59554 22542 59556 22594
rect 59276 22540 59556 22542
rect 59500 22530 59556 22540
rect 59164 22484 59220 22494
rect 58716 22082 58772 22092
rect 59052 22258 59108 22270
rect 59052 22206 59054 22258
rect 59106 22206 59108 22258
rect 58380 21970 58436 21980
rect 59052 21812 59108 22206
rect 59164 22258 59220 22428
rect 59164 22206 59166 22258
rect 59218 22206 59220 22258
rect 59164 22194 59220 22206
rect 59388 22148 59444 22186
rect 59388 22082 59444 22092
rect 59724 22148 59780 23436
rect 60060 23380 60116 23662
rect 60284 23716 60340 24556
rect 60396 24050 60452 25340
rect 60620 25284 60676 26126
rect 60732 25732 60788 29596
rect 60844 27746 60900 30044
rect 60844 27694 60846 27746
rect 60898 27694 60900 27746
rect 60844 27634 60900 27694
rect 60844 27582 60846 27634
rect 60898 27582 60900 27634
rect 60844 27570 60900 27582
rect 60732 25666 60788 25676
rect 60844 25284 60900 25294
rect 60620 25228 60844 25284
rect 60396 23998 60398 24050
rect 60450 23998 60452 24050
rect 60396 23986 60452 23998
rect 60732 24610 60788 24622
rect 60732 24558 60734 24610
rect 60786 24558 60788 24610
rect 60284 23650 60340 23660
rect 60396 23828 60452 23838
rect 60060 23314 60116 23324
rect 59948 23154 60004 23166
rect 59948 23102 59950 23154
rect 60002 23102 60004 23154
rect 59948 22932 60004 23102
rect 60060 23156 60116 23166
rect 60060 23062 60116 23100
rect 60172 23154 60228 23166
rect 60172 23102 60174 23154
rect 60226 23102 60228 23154
rect 59948 22866 60004 22876
rect 59836 22484 59892 22494
rect 60172 22484 60228 23102
rect 60284 23154 60340 23166
rect 60284 23102 60286 23154
rect 60338 23102 60340 23154
rect 60284 22594 60340 23102
rect 60284 22542 60286 22594
rect 60338 22542 60340 22594
rect 60284 22530 60340 22542
rect 59836 22390 59892 22428
rect 59948 22428 60228 22484
rect 59724 22082 59780 22092
rect 59948 22260 60004 22428
rect 59172 21980 59436 21990
rect 59228 21924 59276 21980
rect 59332 21924 59380 21980
rect 59172 21914 59436 21924
rect 59052 21746 59108 21756
rect 59500 21812 59556 21822
rect 59500 21718 59556 21756
rect 59164 21700 59220 21710
rect 59052 21588 59108 21598
rect 59164 21588 59220 21644
rect 59052 21586 59220 21588
rect 59052 21534 59054 21586
rect 59106 21534 59220 21586
rect 59052 21532 59220 21534
rect 59052 21522 59108 21532
rect 58604 21476 58660 21486
rect 58268 21474 58660 21476
rect 58268 21422 58606 21474
rect 58658 21422 58660 21474
rect 58268 21420 58660 21422
rect 57932 20636 58212 20692
rect 57820 19348 57876 19358
rect 57820 19254 57876 19292
rect 57708 19122 57764 19134
rect 57708 19070 57710 19122
rect 57762 19070 57764 19122
rect 57596 18676 57652 18686
rect 57708 18676 57764 19070
rect 57596 18674 57764 18676
rect 57596 18622 57598 18674
rect 57650 18622 57764 18674
rect 57596 18620 57764 18622
rect 57596 18610 57652 18620
rect 57484 16884 57540 16894
rect 57484 16790 57540 16828
rect 57708 16772 57764 16782
rect 57708 16678 57764 16716
rect 57484 16210 57540 16222
rect 57484 16158 57486 16210
rect 57538 16158 57540 16210
rect 57484 16100 57540 16158
rect 57484 16034 57540 16044
rect 57372 15988 57428 15998
rect 57372 15538 57428 15932
rect 57820 15988 57876 15998
rect 57820 15894 57876 15932
rect 57596 15876 57652 15886
rect 57596 15782 57652 15820
rect 57372 15486 57374 15538
rect 57426 15486 57428 15538
rect 57372 15474 57428 15486
rect 57148 14700 57540 14756
rect 57036 14644 57092 14654
rect 57036 14550 57092 14588
rect 55132 13918 55134 13970
rect 55186 13918 55188 13970
rect 55132 13906 55188 13918
rect 57148 14530 57204 14542
rect 57148 14478 57150 14530
rect 57202 14478 57204 14530
rect 55132 13748 55188 13758
rect 55020 13746 55188 13748
rect 55020 13694 55134 13746
rect 55186 13694 55188 13746
rect 55020 13692 55188 13694
rect 55132 13682 55188 13692
rect 55468 13748 55524 13758
rect 55468 13746 55748 13748
rect 55468 13694 55470 13746
rect 55522 13694 55748 13746
rect 55468 13692 55748 13694
rect 55468 13682 55524 13692
rect 55356 13300 55412 13310
rect 55356 13186 55412 13244
rect 55356 13134 55358 13186
rect 55410 13134 55412 13186
rect 55356 13122 55412 13134
rect 55692 13186 55748 13692
rect 56924 13412 56980 13422
rect 55692 13134 55694 13186
rect 55746 13134 55748 13186
rect 55692 13122 55748 13134
rect 55916 13188 55972 13198
rect 55132 12964 55188 12974
rect 55132 12870 55188 12908
rect 55916 12404 55972 13132
rect 56140 12964 56196 12974
rect 56140 12870 56196 12908
rect 56924 12738 56980 13356
rect 57148 13076 57204 14478
rect 57148 13010 57204 13020
rect 56924 12686 56926 12738
rect 56978 12686 56980 12738
rect 55244 12292 55300 12302
rect 55916 12272 55972 12348
rect 56588 12404 56644 12414
rect 56588 12310 56644 12348
rect 55244 12198 55300 12236
rect 56476 12178 56532 12190
rect 56476 12126 56478 12178
rect 56530 12126 56532 12178
rect 55132 12068 55188 12078
rect 54908 12066 55188 12068
rect 54908 12014 55134 12066
rect 55186 12014 55188 12066
rect 54908 12012 55188 12014
rect 55132 12002 55188 12012
rect 56476 12068 56532 12126
rect 56476 12002 56532 12012
rect 56812 12178 56868 12190
rect 56812 12126 56814 12178
rect 56866 12126 56868 12178
rect 54236 11508 54292 11518
rect 53004 10782 53006 10834
rect 53058 10782 53060 10834
rect 53004 10770 53060 10782
rect 53116 11004 53732 11060
rect 54124 11394 54180 11406
rect 54124 11342 54126 11394
rect 54178 11342 54180 11394
rect 53116 10834 53172 11004
rect 53116 10782 53118 10834
rect 53170 10782 53172 10834
rect 53116 10770 53172 10782
rect 53228 10724 53284 10734
rect 54124 10724 54180 11342
rect 54236 11172 54292 11452
rect 56364 11508 56420 11518
rect 56364 11414 56420 11452
rect 56812 11396 56868 12126
rect 56924 12068 56980 12686
rect 56924 12002 56980 12012
rect 57372 12628 57428 12638
rect 57260 11508 57316 11518
rect 57036 11396 57092 11406
rect 56812 11340 57036 11396
rect 57036 11302 57092 11340
rect 54236 11116 54404 11172
rect 54236 10724 54292 10734
rect 54124 10722 54292 10724
rect 54124 10670 54238 10722
rect 54290 10670 54292 10722
rect 54124 10668 54292 10670
rect 53228 10630 53284 10668
rect 53676 10612 53732 10622
rect 54012 10612 54068 10622
rect 53676 10610 54068 10612
rect 53676 10558 53678 10610
rect 53730 10558 54014 10610
rect 54066 10558 54068 10610
rect 53676 10556 54068 10558
rect 53676 10546 53732 10556
rect 54012 10546 54068 10556
rect 54236 10612 54292 10668
rect 54348 10722 54404 11116
rect 54348 10670 54350 10722
rect 54402 10670 54404 10722
rect 54348 10658 54404 10670
rect 55020 11170 55076 11182
rect 55020 11118 55022 11170
rect 55074 11118 55076 11170
rect 54236 10546 54292 10556
rect 54796 10612 54852 10622
rect 55020 10612 55076 11118
rect 55804 10836 55860 10846
rect 55804 10742 55860 10780
rect 56476 10836 56532 10846
rect 56476 10742 56532 10780
rect 54852 10556 55076 10612
rect 56588 10612 56644 10622
rect 54796 10518 54852 10556
rect 56588 10518 56644 10556
rect 56700 10500 56756 10510
rect 56700 10406 56756 10444
rect 57260 10050 57316 11452
rect 57372 10388 57428 12572
rect 57484 12292 57540 14700
rect 57932 14308 57988 20636
rect 58492 20580 58548 21420
rect 58604 21410 58660 21420
rect 59948 21474 60004 22204
rect 60396 22372 60452 23772
rect 60732 23828 60788 24558
rect 60844 24612 60900 25228
rect 60844 24546 60900 24556
rect 60732 23762 60788 23772
rect 60844 23716 60900 23726
rect 60620 23380 60676 23390
rect 60620 23154 60676 23324
rect 60620 23102 60622 23154
rect 60674 23102 60676 23154
rect 60620 23090 60676 23102
rect 60620 22484 60676 22494
rect 60620 22390 60676 22428
rect 60172 22148 60228 22158
rect 60396 22148 60452 22316
rect 60172 22146 60452 22148
rect 60172 22094 60174 22146
rect 60226 22094 60452 22146
rect 60172 22092 60452 22094
rect 60172 22082 60228 22092
rect 59948 21422 59950 21474
rect 60002 21422 60004 21474
rect 58716 20916 58772 20926
rect 58716 20822 58772 20860
rect 59612 20916 59668 20926
rect 58604 20804 58660 20814
rect 58604 20710 58660 20748
rect 58492 20524 58772 20580
rect 58044 19236 58100 19246
rect 58044 19142 58100 19180
rect 58492 19236 58548 19246
rect 58156 18788 58212 18798
rect 58044 18450 58100 18462
rect 58044 18398 58046 18450
rect 58098 18398 58100 18450
rect 58044 17556 58100 18398
rect 58044 17462 58100 17500
rect 58156 18450 58212 18732
rect 58156 18398 58158 18450
rect 58210 18398 58212 18450
rect 58044 17332 58100 17342
rect 58156 17332 58212 18398
rect 58100 17276 58212 17332
rect 58268 18676 58324 18686
rect 58268 18450 58324 18620
rect 58268 18398 58270 18450
rect 58322 18398 58324 18450
rect 58268 17554 58324 18398
rect 58492 17778 58548 19180
rect 58492 17726 58494 17778
rect 58546 17726 58548 17778
rect 58492 17714 58548 17726
rect 58268 17502 58270 17554
rect 58322 17502 58324 17554
rect 58044 17106 58100 17276
rect 58044 17054 58046 17106
rect 58098 17054 58100 17106
rect 58044 17042 58100 17054
rect 58268 15148 58324 17502
rect 58604 17554 58660 17566
rect 58604 17502 58606 17554
rect 58658 17502 58660 17554
rect 58604 17332 58660 17502
rect 58604 17266 58660 17276
rect 58044 15092 58324 15148
rect 58044 14754 58100 15092
rect 58044 14702 58046 14754
rect 58098 14702 58100 14754
rect 58044 14690 58100 14702
rect 58156 14644 58212 14654
rect 58156 14418 58212 14588
rect 58156 14366 58158 14418
rect 58210 14366 58212 14418
rect 57484 12160 57540 12236
rect 57596 14252 57988 14308
rect 58044 14306 58100 14318
rect 58044 14254 58046 14306
rect 58098 14254 58100 14306
rect 57484 10612 57540 10650
rect 57484 10546 57540 10556
rect 57372 10332 57540 10388
rect 57260 9998 57262 10050
rect 57314 9998 57316 10050
rect 57260 9986 57316 9998
rect 52780 9650 52836 9660
rect 56700 9826 56756 9838
rect 56700 9774 56702 9826
rect 56754 9774 56756 9826
rect 52108 9604 52164 9614
rect 52108 9602 52276 9604
rect 52108 9550 52110 9602
rect 52162 9550 52276 9602
rect 52108 9548 52276 9550
rect 52108 9538 52164 9548
rect 52108 9268 52164 9278
rect 52108 9042 52164 9212
rect 52108 8990 52110 9042
rect 52162 8990 52164 9042
rect 52108 8978 52164 8990
rect 51100 8418 51156 8428
rect 51772 8372 52052 8428
rect 50540 8318 50542 8370
rect 50594 8318 50596 8370
rect 50540 8306 50596 8318
rect 50316 8194 50372 8204
rect 50764 8260 50820 8270
rect 50764 8166 50820 8204
rect 48188 7634 48244 7644
rect 48524 8146 48580 8158
rect 48524 8094 48526 8146
rect 48578 8094 48580 8146
rect 48524 8036 48580 8094
rect 51884 8146 51940 8158
rect 51884 8094 51886 8146
rect 51938 8094 51940 8146
rect 48300 7586 48356 7598
rect 48300 7534 48302 7586
rect 48354 7534 48356 7586
rect 47404 7476 47460 7486
rect 48300 7476 48356 7534
rect 47404 7474 48356 7476
rect 47404 7422 47406 7474
rect 47458 7422 48356 7474
rect 47404 7420 48356 7422
rect 47404 7410 47460 7420
rect 47292 7362 47348 7374
rect 47292 7310 47294 7362
rect 47346 7310 47348 7362
rect 47292 7252 47348 7310
rect 47292 7186 47348 7196
rect 46676 6748 46900 6804
rect 47404 6916 47460 6926
rect 45388 6466 45444 6478
rect 45388 6414 45390 6466
rect 45442 6414 45444 6466
rect 45388 5908 45444 6414
rect 46508 6468 46564 6478
rect 45948 6356 46004 6366
rect 45948 6130 46004 6300
rect 45948 6078 45950 6130
rect 46002 6078 46004 6130
rect 45948 6066 46004 6078
rect 46172 6132 46228 6142
rect 46172 6038 46228 6076
rect 45836 5908 45892 5918
rect 46284 5908 46340 5918
rect 45388 5906 45892 5908
rect 45388 5854 45838 5906
rect 45890 5854 45892 5906
rect 45388 5852 45892 5854
rect 45724 5236 45780 5246
rect 45388 5124 45444 5134
rect 45276 5122 45444 5124
rect 45276 5070 45390 5122
rect 45442 5070 45444 5122
rect 45276 5068 45444 5070
rect 45388 5058 45444 5068
rect 44940 4946 44996 4956
rect 45612 5012 45668 5022
rect 44716 4722 44772 4732
rect 44380 4284 45220 4340
rect 44044 3556 44100 4284
rect 45164 3666 45220 4284
rect 45164 3614 45166 3666
rect 45218 3614 45220 3666
rect 45164 3602 45220 3614
rect 45388 3780 45444 3790
rect 44044 3462 44100 3500
rect 44940 3554 44996 3566
rect 44940 3502 44942 3554
rect 44994 3502 44996 3554
rect 44940 3332 44996 3502
rect 45388 3554 45444 3724
rect 45500 3668 45556 3678
rect 45612 3668 45668 4956
rect 45724 5010 45780 5180
rect 45724 4958 45726 5010
rect 45778 4958 45780 5010
rect 45724 4946 45780 4958
rect 45836 4900 45892 5852
rect 46172 5906 46340 5908
rect 46172 5854 46286 5906
rect 46338 5854 46340 5906
rect 46172 5852 46340 5854
rect 46060 5796 46116 5806
rect 46060 5702 46116 5740
rect 45836 4834 45892 4844
rect 46172 5460 46228 5852
rect 46284 5842 46340 5852
rect 46508 5572 46564 6412
rect 46508 5506 46564 5516
rect 46172 4564 46228 5404
rect 46396 5348 46452 5358
rect 46396 5254 46452 5292
rect 46508 5010 46564 5022
rect 46508 4958 46510 5010
rect 46562 4958 46564 5010
rect 46396 4900 46452 4910
rect 46172 4498 46228 4508
rect 46284 4898 46452 4900
rect 46284 4846 46398 4898
rect 46450 4846 46452 4898
rect 46284 4844 46452 4846
rect 45500 3666 45668 3668
rect 45500 3614 45502 3666
rect 45554 3614 45668 3666
rect 45500 3612 45668 3614
rect 45500 3602 45556 3612
rect 45388 3502 45390 3554
rect 45442 3502 45444 3554
rect 45388 3490 45444 3502
rect 44940 3266 44996 3276
rect 45276 3444 45332 3454
rect 43932 1474 43988 1484
rect 45276 800 45332 3388
rect 46284 3442 46340 4844
rect 46396 4834 46452 4844
rect 46508 4676 46564 4958
rect 46508 4610 46564 4620
rect 46284 3390 46286 3442
rect 46338 3390 46340 3442
rect 45612 3330 45668 3342
rect 45612 3278 45614 3330
rect 45666 3278 45668 3330
rect 45612 3108 45668 3278
rect 46284 3220 46340 3390
rect 46284 3154 46340 3164
rect 45612 3042 45668 3052
rect 46620 868 46676 6748
rect 47068 6468 47124 6478
rect 47068 6374 47124 6412
rect 47404 6466 47460 6860
rect 47404 6414 47406 6466
rect 47458 6414 47460 6466
rect 46732 6020 46788 6030
rect 46732 4900 46788 5964
rect 46844 5794 46900 5806
rect 47292 5796 47348 5806
rect 46844 5742 46846 5794
rect 46898 5742 46900 5794
rect 46844 5460 46900 5742
rect 46844 5394 46900 5404
rect 47068 5794 47348 5796
rect 47068 5742 47294 5794
rect 47346 5742 47348 5794
rect 47068 5740 47348 5742
rect 46732 4834 46788 4844
rect 46844 4788 46900 4798
rect 47068 4788 47124 5740
rect 47292 5730 47348 5740
rect 46900 4732 47124 4788
rect 47180 5572 47236 5582
rect 46844 3666 46900 4732
rect 46956 4564 47012 4574
rect 46956 4470 47012 4508
rect 46844 3614 46846 3666
rect 46898 3614 46900 3666
rect 46844 3602 46900 3614
rect 47180 2548 47236 5516
rect 47404 5460 47460 6414
rect 47852 6804 47908 6814
rect 47852 6466 47908 6748
rect 48300 6692 48356 7420
rect 48412 7474 48468 7486
rect 48412 7422 48414 7474
rect 48466 7422 48468 7474
rect 48412 7252 48468 7422
rect 48412 7186 48468 7196
rect 48524 7140 48580 7980
rect 48636 8034 48692 8046
rect 48636 7982 48638 8034
rect 48690 7982 48692 8034
rect 48636 7700 48692 7982
rect 48636 7634 48692 7644
rect 48860 8034 48916 8046
rect 48860 7982 48862 8034
rect 48914 7982 48916 8034
rect 48860 7588 48916 7982
rect 49196 8036 49252 8046
rect 49196 7942 49252 7980
rect 49644 8034 49700 8046
rect 49644 7982 49646 8034
rect 49698 7982 49700 8034
rect 49644 7700 49700 7982
rect 49644 7634 49700 7644
rect 50428 8034 50484 8046
rect 50428 7982 50430 8034
rect 50482 7982 50484 8034
rect 48860 7522 48916 7532
rect 49308 7588 49364 7598
rect 48524 7074 48580 7084
rect 49196 7028 49252 7038
rect 48300 6636 48580 6692
rect 47852 6414 47854 6466
rect 47906 6414 47908 6466
rect 47852 6356 47908 6414
rect 47852 6290 47908 6300
rect 48300 6466 48356 6478
rect 48300 6414 48302 6466
rect 48354 6414 48356 6466
rect 47404 5394 47460 5404
rect 47516 6132 47572 6142
rect 47404 4564 47460 4574
rect 47292 4452 47348 4462
rect 47292 3668 47348 4396
rect 47404 4450 47460 4508
rect 47516 4562 47572 6076
rect 48300 6132 48356 6414
rect 48300 6066 48356 6076
rect 48524 6130 48580 6636
rect 48860 6580 48916 6590
rect 48748 6466 48804 6478
rect 48748 6414 48750 6466
rect 48802 6414 48804 6466
rect 48748 6356 48804 6414
rect 48524 6078 48526 6130
rect 48578 6078 48580 6130
rect 48524 6066 48580 6078
rect 48636 6132 48692 6142
rect 48636 6038 48692 6076
rect 48412 5906 48468 5918
rect 48412 5854 48414 5906
rect 48466 5854 48468 5906
rect 48188 5796 48244 5806
rect 48188 5702 48244 5740
rect 47964 5682 48020 5694
rect 47964 5630 47966 5682
rect 48018 5630 48020 5682
rect 47628 5348 47684 5358
rect 47628 5122 47684 5292
rect 47964 5348 48020 5630
rect 47964 5282 48020 5292
rect 47628 5070 47630 5122
rect 47682 5070 47684 5122
rect 47628 5058 47684 5070
rect 47740 5234 47796 5246
rect 47740 5182 47742 5234
rect 47794 5182 47796 5234
rect 47516 4510 47518 4562
rect 47570 4510 47572 4562
rect 47516 4498 47572 4510
rect 47404 4398 47406 4450
rect 47458 4398 47460 4450
rect 47404 4004 47460 4398
rect 47404 3938 47460 3948
rect 47516 4116 47572 4126
rect 47740 4116 47796 5182
rect 48412 5124 48468 5854
rect 48636 5572 48692 5582
rect 48412 5058 48468 5068
rect 48524 5348 48580 5358
rect 48412 4564 48468 4574
rect 48524 4564 48580 5292
rect 48412 4562 48580 4564
rect 48412 4510 48414 4562
rect 48466 4510 48580 4562
rect 48412 4508 48580 4510
rect 48636 4562 48692 5516
rect 48748 4676 48804 6300
rect 48748 4610 48804 4620
rect 48636 4510 48638 4562
rect 48690 4510 48692 4562
rect 48412 4498 48468 4508
rect 47516 4114 47796 4116
rect 47516 4062 47518 4114
rect 47570 4062 47796 4114
rect 47516 4060 47796 4062
rect 47404 3668 47460 3678
rect 47292 3666 47460 3668
rect 47292 3614 47406 3666
rect 47458 3614 47460 3666
rect 47292 3612 47460 3614
rect 47404 3602 47460 3612
rect 47516 3332 47572 4060
rect 47516 3266 47572 3276
rect 47628 3556 47684 3566
rect 47628 3108 47684 3500
rect 47964 3444 48020 3454
rect 47964 3350 48020 3388
rect 48636 3332 48692 4510
rect 48748 4340 48804 4350
rect 48860 4340 48916 6524
rect 49196 5346 49252 6972
rect 49308 6916 49364 7532
rect 50428 7588 50484 7982
rect 50652 8034 50708 8046
rect 50652 7982 50654 8034
rect 50706 7982 50708 8034
rect 50652 7924 50708 7982
rect 50652 7858 50708 7868
rect 51548 8034 51604 8046
rect 51548 7982 51550 8034
rect 51602 7982 51604 8034
rect 50428 7522 50484 7532
rect 49868 7474 49924 7486
rect 49868 7422 49870 7474
rect 49922 7422 49924 7474
rect 49512 7084 49776 7094
rect 49568 7028 49616 7084
rect 49672 7028 49720 7084
rect 49512 7018 49776 7028
rect 49308 6860 49588 6916
rect 49532 6802 49588 6860
rect 49532 6750 49534 6802
rect 49586 6750 49588 6802
rect 49532 6738 49588 6750
rect 49756 6244 49812 6254
rect 49644 6020 49700 6030
rect 49532 5964 49644 6020
rect 49532 5796 49588 5964
rect 49644 5926 49700 5964
rect 49756 6018 49812 6188
rect 49756 5966 49758 6018
rect 49810 5966 49812 6018
rect 49756 5954 49812 5966
rect 49868 6132 49924 7422
rect 51100 7474 51156 7486
rect 51100 7422 51102 7474
rect 51154 7422 51156 7474
rect 50092 7362 50148 7374
rect 50092 7310 50094 7362
rect 50146 7310 50148 7362
rect 50092 6916 50148 7310
rect 50092 6784 50148 6860
rect 50876 6916 50932 6926
rect 50876 6822 50932 6860
rect 49532 5730 49588 5740
rect 49644 5684 49700 5694
rect 49868 5684 49924 6076
rect 49980 6580 50036 6590
rect 49980 6020 50036 6524
rect 49980 5954 50036 5964
rect 50092 6466 50148 6478
rect 50092 6414 50094 6466
rect 50146 6414 50148 6466
rect 50092 5908 50148 6414
rect 51100 6468 51156 7422
rect 51548 7476 51604 7982
rect 51772 8034 51828 8046
rect 51772 7982 51774 8034
rect 51826 7982 51828 8034
rect 51772 7812 51828 7982
rect 51772 7746 51828 7756
rect 51324 7252 51380 7262
rect 51324 7158 51380 7196
rect 51212 6692 51268 6702
rect 51212 6598 51268 6636
rect 51548 6690 51604 7420
rect 51884 7364 51940 8094
rect 51884 7298 51940 7308
rect 51548 6638 51550 6690
rect 51602 6638 51604 6690
rect 51548 6626 51604 6638
rect 51996 6692 52052 8372
rect 51996 6626 52052 6636
rect 51436 6580 51492 6590
rect 51436 6486 51492 6524
rect 51100 6402 51156 6412
rect 51324 6466 51380 6478
rect 51324 6414 51326 6466
rect 51378 6414 51380 6466
rect 51324 6244 51380 6414
rect 52108 6466 52164 6478
rect 52108 6414 52110 6466
rect 52162 6414 52164 6466
rect 50092 5842 50148 5852
rect 51100 6188 51716 6244
rect 49644 5682 49924 5684
rect 49644 5630 49646 5682
rect 49698 5630 49924 5682
rect 49644 5628 49924 5630
rect 50204 5794 50260 5806
rect 50204 5742 50206 5794
rect 50258 5742 50260 5794
rect 49644 5618 49700 5628
rect 49512 5516 49776 5526
rect 49568 5460 49616 5516
rect 49672 5460 49720 5516
rect 49512 5450 49776 5460
rect 49196 5294 49198 5346
rect 49250 5294 49252 5346
rect 49196 5282 49252 5294
rect 49308 5124 49364 5134
rect 49308 5030 49364 5068
rect 50204 4564 50260 5742
rect 50652 5796 50708 5806
rect 50652 5702 50708 5740
rect 50428 5236 50484 5246
rect 50428 5142 50484 5180
rect 50204 4498 50260 4508
rect 50540 5124 50596 5134
rect 50540 4562 50596 5068
rect 51100 5122 51156 6188
rect 51660 6130 51716 6188
rect 51660 6078 51662 6130
rect 51714 6078 51716 6130
rect 51660 6066 51716 6078
rect 52108 6132 52164 6414
rect 52108 6066 52164 6076
rect 51436 6018 51492 6030
rect 51436 5966 51438 6018
rect 51490 5966 51492 6018
rect 51324 5906 51380 5918
rect 51324 5854 51326 5906
rect 51378 5854 51380 5906
rect 51100 5070 51102 5122
rect 51154 5070 51156 5122
rect 51100 5058 51156 5070
rect 51212 5796 51268 5806
rect 50540 4510 50542 4562
rect 50594 4510 50596 4562
rect 50540 4498 50596 4510
rect 50988 5012 51044 5022
rect 49756 4452 49812 4462
rect 49812 4396 49924 4452
rect 49756 4358 49812 4396
rect 48748 4338 48916 4340
rect 48748 4286 48750 4338
rect 48802 4286 48916 4338
rect 48748 4284 48916 4286
rect 48748 4274 48804 4284
rect 48636 3266 48692 3276
rect 48748 3442 48804 3454
rect 48748 3390 48750 3442
rect 48802 3390 48804 3442
rect 48748 3220 48804 3390
rect 48748 3154 48804 3164
rect 47180 2482 47236 2492
rect 47404 3052 47684 3108
rect 46620 802 46676 812
rect 47404 800 47460 3052
rect 48860 2996 48916 4284
rect 49512 3948 49776 3958
rect 49568 3892 49616 3948
rect 49672 3892 49720 3948
rect 49512 3882 49776 3892
rect 49868 3780 49924 4396
rect 50092 4450 50148 4462
rect 50092 4398 50094 4450
rect 50146 4398 50148 4450
rect 50092 4340 50148 4398
rect 50092 4274 50148 4284
rect 50764 4450 50820 4462
rect 50764 4398 50766 4450
rect 50818 4398 50820 4450
rect 50764 4340 50820 4398
rect 50764 4274 50820 4284
rect 50876 4338 50932 4350
rect 50876 4286 50878 4338
rect 50930 4286 50932 4338
rect 48860 2930 48916 2940
rect 49532 3724 49924 3780
rect 49532 800 49588 3724
rect 50876 3668 50932 4286
rect 50876 3602 50932 3612
rect 50988 3556 51044 4956
rect 50988 3442 51044 3500
rect 50988 3390 50990 3442
rect 51042 3390 51044 3442
rect 50988 3378 51044 3390
rect 51212 1204 51268 5740
rect 51324 5572 51380 5854
rect 51436 5684 51492 5966
rect 51436 5618 51492 5628
rect 51548 6020 51604 6030
rect 51324 4788 51380 5516
rect 51324 4722 51380 4732
rect 51548 4450 51604 5964
rect 51996 5908 52052 5918
rect 51996 5814 52052 5852
rect 52220 5684 52276 9548
rect 52556 9602 52612 9614
rect 52556 9550 52558 9602
rect 52610 9550 52612 9602
rect 52332 8034 52388 8046
rect 52332 7982 52334 8034
rect 52386 7982 52388 8034
rect 52332 7924 52388 7982
rect 52332 7858 52388 7868
rect 52444 7812 52500 7822
rect 52444 7586 52500 7756
rect 52444 7534 52446 7586
rect 52498 7534 52500 7586
rect 52444 7522 52500 7534
rect 52220 5618 52276 5628
rect 52332 7364 52388 7374
rect 52332 6804 52388 7308
rect 52556 6916 52612 9550
rect 53788 9602 53844 9614
rect 53788 9550 53790 9602
rect 53842 9550 53844 9602
rect 52780 8932 52836 8942
rect 52780 8838 52836 8876
rect 53564 8930 53620 8942
rect 53564 8878 53566 8930
rect 53618 8878 53620 8930
rect 53564 8428 53620 8878
rect 53564 8372 53732 8428
rect 53340 8034 53396 8046
rect 53340 7982 53342 8034
rect 53394 7982 53396 8034
rect 53340 7812 53396 7982
rect 53396 7756 53620 7812
rect 53340 7746 53396 7756
rect 53564 7698 53620 7756
rect 53564 7646 53566 7698
rect 53618 7646 53620 7698
rect 53564 7634 53620 7646
rect 52668 7474 52724 7486
rect 52668 7422 52670 7474
rect 52722 7422 52724 7474
rect 52668 7364 52724 7422
rect 52892 7474 52948 7486
rect 52892 7422 52894 7474
rect 52946 7422 52948 7474
rect 52668 7298 52724 7308
rect 52780 7362 52836 7374
rect 52780 7310 52782 7362
rect 52834 7310 52836 7362
rect 52556 6860 52724 6916
rect 51772 5348 51828 5358
rect 51772 5122 51828 5292
rect 51772 5070 51774 5122
rect 51826 5070 51828 5122
rect 51772 5058 51828 5070
rect 52108 5122 52164 5134
rect 52108 5070 52110 5122
rect 52162 5070 52164 5122
rect 51548 4398 51550 4450
rect 51602 4398 51604 4450
rect 51324 4340 51380 4350
rect 51324 3108 51380 4284
rect 51548 4228 51604 4398
rect 51660 4676 51716 4686
rect 51660 4450 51716 4620
rect 51660 4398 51662 4450
rect 51714 4398 51716 4450
rect 51660 4386 51716 4398
rect 52108 4340 52164 5070
rect 52332 4340 52388 6748
rect 52556 6692 52612 6702
rect 52556 6598 52612 6636
rect 52444 6244 52500 6254
rect 52444 6130 52500 6188
rect 52444 6078 52446 6130
rect 52498 6078 52500 6130
rect 52444 4676 52500 6078
rect 52444 4610 52500 4620
rect 52444 4340 52500 4350
rect 52332 4338 52500 4340
rect 52332 4286 52446 4338
rect 52498 4286 52500 4338
rect 52332 4284 52500 4286
rect 52108 4274 52164 4284
rect 52444 4274 52500 4284
rect 51548 4162 51604 4172
rect 51324 3042 51380 3052
rect 51660 3556 51716 3566
rect 51212 1138 51268 1148
rect 51660 800 51716 3500
rect 52668 3556 52724 6860
rect 52780 6692 52836 7310
rect 52892 6916 52948 7422
rect 53004 7474 53060 7486
rect 53004 7422 53006 7474
rect 53058 7422 53060 7474
rect 53004 7028 53060 7422
rect 53676 7028 53732 8372
rect 53788 8034 53844 9550
rect 54348 9604 54404 9614
rect 54460 9604 54516 9614
rect 54348 9602 54460 9604
rect 54348 9550 54350 9602
rect 54402 9550 54460 9602
rect 54348 9548 54460 9550
rect 54348 9538 54404 9548
rect 54348 9380 54404 9390
rect 54348 9154 54404 9324
rect 54348 9102 54350 9154
rect 54402 9102 54404 9154
rect 54348 9090 54404 9102
rect 53788 7982 53790 8034
rect 53842 7982 53844 8034
rect 53788 7364 53844 7982
rect 53788 7298 53844 7308
rect 54236 8148 54292 8158
rect 54236 8034 54292 8092
rect 54236 7982 54238 8034
rect 54290 7982 54292 8034
rect 53060 6972 53172 7028
rect 53004 6962 53060 6972
rect 52892 6850 52948 6860
rect 52780 6626 52836 6636
rect 52892 5794 52948 5806
rect 52892 5742 52894 5794
rect 52946 5742 52948 5794
rect 52892 5684 52948 5742
rect 52892 5618 52948 5628
rect 53004 4676 53060 4686
rect 53004 4562 53060 4620
rect 53004 4510 53006 4562
rect 53058 4510 53060 4562
rect 53004 4498 53060 4510
rect 53116 4228 53172 6972
rect 53676 6962 53732 6972
rect 54236 6916 54292 7982
rect 54348 6916 54404 6926
rect 54236 6860 54348 6916
rect 53340 6468 53396 6478
rect 53228 6466 53396 6468
rect 53228 6414 53342 6466
rect 53394 6414 53396 6466
rect 53228 6412 53396 6414
rect 53228 4452 53284 6412
rect 53340 6402 53396 6412
rect 53564 6468 53620 6478
rect 53340 6132 53396 6142
rect 53340 6038 53396 6076
rect 53228 4386 53284 4396
rect 53340 5684 53396 5694
rect 53116 4162 53172 4172
rect 53340 3666 53396 5628
rect 53564 5346 53620 6412
rect 53900 6466 53956 6478
rect 53900 6414 53902 6466
rect 53954 6414 53956 6466
rect 53900 6020 53956 6414
rect 53564 5294 53566 5346
rect 53618 5294 53620 5346
rect 53564 5124 53620 5294
rect 53564 5058 53620 5068
rect 53788 5794 53844 5806
rect 53788 5742 53790 5794
rect 53842 5742 53844 5794
rect 53676 5010 53732 5022
rect 53676 4958 53678 5010
rect 53730 4958 53732 5010
rect 53340 3614 53342 3666
rect 53394 3614 53396 3666
rect 53340 3602 53396 3614
rect 53564 4898 53620 4910
rect 53564 4846 53566 4898
rect 53618 4846 53620 4898
rect 53564 4452 53620 4846
rect 52780 3556 52836 3566
rect 52724 3554 52836 3556
rect 52724 3502 52782 3554
rect 52834 3502 52836 3554
rect 52724 3500 52836 3502
rect 51772 3444 51828 3454
rect 52668 3424 52724 3500
rect 52780 3490 52836 3500
rect 51772 3350 51828 3388
rect 53564 3332 53620 4396
rect 53676 4788 53732 4958
rect 53788 5012 53844 5742
rect 53900 5236 53956 5964
rect 54348 5796 54404 6860
rect 54460 6356 54516 9548
rect 54796 9604 54852 9614
rect 54796 9602 55076 9604
rect 54796 9550 54798 9602
rect 54850 9550 55076 9602
rect 54796 9548 55076 9550
rect 54796 9538 54852 9548
rect 54796 9156 54852 9166
rect 54684 9044 54740 9054
rect 54684 8930 54740 8988
rect 54684 8878 54686 8930
rect 54738 8878 54740 8930
rect 54684 8484 54740 8878
rect 54796 9042 54852 9100
rect 54796 8990 54798 9042
rect 54850 8990 54852 9042
rect 54796 8932 54852 8990
rect 54796 8866 54852 8876
rect 54908 8484 54964 8494
rect 54684 8482 54964 8484
rect 54684 8430 54910 8482
rect 54962 8430 54964 8482
rect 54684 8428 54964 8430
rect 54908 8418 54964 8428
rect 54572 7476 54628 7486
rect 54572 7382 54628 7420
rect 54684 7362 54740 7374
rect 54684 7310 54686 7362
rect 54738 7310 54740 7362
rect 54684 7028 54740 7310
rect 54684 6914 54740 6972
rect 54684 6862 54686 6914
rect 54738 6862 54740 6914
rect 54684 6850 54740 6862
rect 54572 6692 54628 6702
rect 54572 6690 54852 6692
rect 54572 6638 54574 6690
rect 54626 6638 54852 6690
rect 54572 6636 54852 6638
rect 54572 6626 54628 6636
rect 54460 6020 54516 6300
rect 54684 6466 54740 6478
rect 54684 6414 54686 6466
rect 54738 6414 54740 6466
rect 54684 6020 54740 6414
rect 54460 5964 54628 6020
rect 54460 5796 54516 5806
rect 54348 5794 54516 5796
rect 54348 5742 54462 5794
rect 54514 5742 54516 5794
rect 54348 5740 54516 5742
rect 53900 5170 53956 5180
rect 54012 5572 54068 5582
rect 53788 4946 53844 4956
rect 53676 4562 53732 4732
rect 53676 4510 53678 4562
rect 53730 4510 53732 4562
rect 53676 4340 53732 4510
rect 53676 4274 53732 4284
rect 53900 4676 53956 4686
rect 53900 3666 53956 4620
rect 53900 3614 53902 3666
rect 53954 3614 53956 3666
rect 53900 3602 53956 3614
rect 53564 3266 53620 3276
rect 53788 2884 53844 2894
rect 53788 800 53844 2828
rect 54012 2212 54068 5516
rect 54460 5572 54516 5740
rect 54460 5506 54516 5516
rect 54460 4900 54516 4910
rect 54348 4898 54516 4900
rect 54348 4846 54462 4898
rect 54514 4846 54516 4898
rect 54348 4844 54516 4846
rect 54124 4228 54180 4238
rect 54124 4134 54180 4172
rect 54012 2146 54068 2156
rect 54348 1652 54404 4844
rect 54460 4834 54516 4844
rect 54460 3556 54516 3566
rect 54572 3556 54628 5964
rect 54684 5954 54740 5964
rect 54796 5796 54852 6636
rect 54908 5908 54964 5918
rect 54908 5814 54964 5852
rect 54796 5730 54852 5740
rect 55020 5684 55076 9548
rect 55244 9602 55300 9614
rect 55244 9550 55246 9602
rect 55298 9550 55300 9602
rect 55244 8428 55300 9550
rect 55916 9604 55972 9614
rect 55916 9602 56308 9604
rect 55916 9550 55918 9602
rect 55970 9550 56308 9602
rect 55916 9548 56308 9550
rect 55916 9538 55972 9548
rect 56140 9156 56196 9166
rect 56140 9062 56196 9100
rect 55916 9044 55972 9054
rect 55916 8950 55972 8988
rect 56028 8932 56084 8942
rect 56028 8838 56084 8876
rect 55132 8372 55300 8428
rect 55580 8372 55636 8382
rect 55132 8148 55188 8372
rect 55580 8278 55636 8316
rect 55132 8082 55188 8092
rect 55468 8258 55524 8270
rect 55468 8206 55470 8258
rect 55522 8206 55524 8258
rect 55356 7028 55412 7038
rect 55356 6914 55412 6972
rect 55356 6862 55358 6914
rect 55410 6862 55412 6914
rect 55356 6850 55412 6862
rect 55468 6580 55524 8206
rect 56140 7474 56196 7486
rect 56140 7422 56142 7474
rect 56194 7422 56196 7474
rect 55692 7364 55748 7374
rect 55580 6692 55636 6702
rect 55580 6598 55636 6636
rect 55468 6514 55524 6524
rect 55692 6468 55748 7308
rect 55916 7028 55972 7038
rect 55916 6802 55972 6972
rect 55916 6750 55918 6802
rect 55970 6750 55972 6802
rect 55916 6738 55972 6750
rect 55804 6692 55860 6730
rect 55804 6626 55860 6636
rect 56028 6692 56084 6702
rect 56028 6598 56084 6636
rect 55580 6412 55748 6468
rect 55580 6132 55636 6412
rect 56028 6244 56084 6254
rect 55804 6132 55860 6142
rect 55580 6130 55860 6132
rect 55580 6078 55806 6130
rect 55858 6078 55860 6130
rect 55580 6076 55860 6078
rect 55804 6066 55860 6076
rect 56028 6130 56084 6188
rect 56028 6078 56030 6130
rect 56082 6078 56084 6130
rect 54908 5628 55076 5684
rect 55356 6020 55412 6030
rect 54796 5012 54852 5022
rect 54684 4900 54740 4910
rect 54684 4806 54740 4844
rect 54796 4788 54852 4956
rect 54796 4722 54852 4732
rect 54796 4452 54852 4462
rect 54796 4228 54852 4396
rect 54908 4340 54964 5628
rect 55356 5122 55412 5964
rect 56028 6020 56084 6078
rect 56140 6132 56196 7422
rect 56140 6066 56196 6076
rect 56028 5954 56084 5964
rect 55468 5908 55524 5918
rect 55468 5460 55524 5852
rect 55580 5906 55636 5918
rect 55580 5854 55582 5906
rect 55634 5854 55636 5906
rect 55580 5572 55636 5854
rect 55916 5908 55972 5918
rect 55916 5814 55972 5852
rect 56140 5906 56196 5918
rect 56140 5854 56142 5906
rect 56194 5854 56196 5906
rect 55580 5506 55636 5516
rect 56140 5684 56196 5854
rect 55468 5394 55524 5404
rect 55356 5070 55358 5122
rect 55410 5070 55412 5122
rect 55020 5012 55076 5022
rect 55020 4676 55076 4956
rect 55020 4610 55076 4620
rect 55244 4452 55300 4462
rect 55020 4340 55076 4350
rect 54908 4284 55020 4340
rect 54796 4162 54852 4172
rect 55020 3666 55076 4284
rect 55020 3614 55022 3666
rect 55074 3614 55076 3666
rect 55020 3602 55076 3614
rect 55132 4338 55188 4350
rect 55132 4286 55134 4338
rect 55186 4286 55188 4338
rect 54460 3554 54628 3556
rect 54460 3502 54462 3554
rect 54514 3502 54628 3554
rect 54460 3500 54628 3502
rect 54460 3490 54516 3500
rect 55132 2884 55188 4286
rect 55244 4116 55300 4396
rect 55244 4050 55300 4060
rect 55132 2818 55188 2828
rect 54348 1586 54404 1596
rect 55356 1092 55412 5070
rect 55580 5012 55636 5022
rect 55468 4956 55580 5012
rect 55468 3668 55524 4956
rect 55580 4946 55636 4956
rect 55916 4900 55972 4910
rect 55916 4806 55972 4844
rect 56140 4564 56196 5628
rect 56140 4498 56196 4508
rect 56140 4340 56196 4350
rect 56252 4340 56308 9548
rect 56700 9492 56756 9774
rect 57372 9826 57428 9838
rect 57372 9774 57374 9826
rect 57426 9774 57428 9826
rect 57372 9604 57428 9774
rect 57372 9538 57428 9548
rect 56700 9426 56756 9436
rect 57372 9380 57428 9390
rect 56588 9042 56644 9054
rect 56588 8990 56590 9042
rect 56642 8990 56644 9042
rect 56588 8482 56644 8990
rect 56588 8430 56590 8482
rect 56642 8430 56644 8482
rect 56588 8418 56644 8430
rect 57372 8482 57428 9324
rect 57484 9042 57540 10332
rect 57484 8990 57486 9042
rect 57538 8990 57540 9042
rect 57484 8978 57540 8990
rect 57372 8430 57374 8482
rect 57426 8430 57428 8482
rect 57372 8418 57428 8430
rect 56700 8372 56756 8382
rect 56700 8258 56756 8316
rect 56700 8206 56702 8258
rect 56754 8206 56756 8258
rect 56588 8034 56644 8046
rect 56588 7982 56590 8034
rect 56642 7982 56644 8034
rect 56476 6692 56532 6702
rect 56364 5460 56420 5470
rect 56364 5012 56420 5404
rect 56476 5348 56532 6636
rect 56588 6580 56644 7982
rect 56700 7586 56756 8206
rect 57484 8260 57540 8270
rect 57484 8166 57540 8204
rect 57372 8036 57428 8046
rect 56700 7534 56702 7586
rect 56754 7534 56756 7586
rect 56700 7522 56756 7534
rect 57260 7980 57372 8036
rect 56812 6692 56868 6702
rect 56588 6514 56644 6524
rect 56700 6578 56756 6590
rect 56700 6526 56702 6578
rect 56754 6526 56756 6578
rect 56700 6356 56756 6526
rect 56812 6578 56868 6636
rect 56812 6526 56814 6578
rect 56866 6526 56868 6578
rect 56812 6514 56868 6526
rect 56588 6300 56700 6356
rect 56588 5684 56644 6300
rect 56700 6224 56756 6300
rect 57036 6466 57092 6478
rect 57036 6414 57038 6466
rect 57090 6414 57092 6466
rect 57036 6132 57092 6414
rect 57036 6066 57092 6076
rect 56700 5796 56756 5806
rect 56700 5794 56868 5796
rect 56700 5742 56702 5794
rect 56754 5742 56868 5794
rect 56700 5740 56868 5742
rect 56700 5730 56756 5740
rect 56588 5618 56644 5628
rect 56588 5348 56644 5358
rect 56476 5292 56588 5348
rect 56588 5254 56644 5292
rect 56588 5124 56644 5134
rect 56588 5012 56644 5068
rect 56364 5010 56644 5012
rect 56364 4958 56590 5010
rect 56642 4958 56644 5010
rect 56364 4956 56644 4958
rect 56476 4562 56532 4956
rect 56588 4946 56644 4956
rect 56700 5010 56756 5022
rect 56700 4958 56702 5010
rect 56754 4958 56756 5010
rect 56476 4510 56478 4562
rect 56530 4510 56532 4562
rect 56476 4498 56532 4510
rect 56700 4676 56756 4958
rect 55916 4338 56308 4340
rect 55916 4286 56142 4338
rect 56194 4286 56308 4338
rect 55916 4284 56308 4286
rect 55580 4226 55636 4238
rect 55580 4174 55582 4226
rect 55634 4174 55636 4226
rect 55580 3892 55636 4174
rect 55580 3826 55636 3836
rect 55468 3554 55524 3612
rect 55468 3502 55470 3554
rect 55522 3502 55524 3554
rect 55468 3490 55524 3502
rect 55356 1026 55412 1036
rect 55916 800 55972 4284
rect 56140 4274 56196 4284
rect 56700 4228 56756 4620
rect 56812 4564 56868 5740
rect 57148 5122 57204 5134
rect 57148 5070 57150 5122
rect 57202 5070 57204 5122
rect 57148 5012 57204 5070
rect 57148 4946 57204 4956
rect 56812 4498 56868 4508
rect 57260 4452 57316 7980
rect 57372 7942 57428 7980
rect 57372 7364 57428 7374
rect 57596 7364 57652 14252
rect 58044 13076 58100 14254
rect 58156 13860 58212 14366
rect 58156 13794 58212 13804
rect 58044 13010 58100 13020
rect 58044 12628 58100 12638
rect 58044 12402 58100 12572
rect 58044 12350 58046 12402
rect 58098 12350 58100 12402
rect 58044 12338 58100 12350
rect 58492 12628 58548 12638
rect 58492 12402 58548 12572
rect 58492 12350 58494 12402
rect 58546 12350 58548 12402
rect 58492 12338 58548 12350
rect 57932 11508 57988 11518
rect 57932 11414 57988 11452
rect 58268 11396 58324 11406
rect 58268 11302 58324 11340
rect 58044 11170 58100 11182
rect 58044 11118 58046 11170
rect 58098 11118 58100 11170
rect 57708 10836 57764 10846
rect 57708 10742 57764 10780
rect 57820 10724 57876 10734
rect 58044 10724 58100 11118
rect 57820 10722 58100 10724
rect 57820 10670 57822 10722
rect 57874 10670 58100 10722
rect 57820 10668 58100 10670
rect 57820 10658 57876 10668
rect 58380 10500 58436 10510
rect 58380 10406 58436 10444
rect 58044 9602 58100 9614
rect 58044 9550 58046 9602
rect 58098 9550 58100 9602
rect 58044 9492 58100 9550
rect 58492 9604 58548 9614
rect 58492 9510 58548 9548
rect 58044 9426 58100 9436
rect 58044 9044 58100 9054
rect 58492 9044 58548 9054
rect 58044 9042 58548 9044
rect 58044 8990 58046 9042
rect 58098 8990 58494 9042
rect 58546 8990 58548 9042
rect 58044 8988 58548 8990
rect 58044 8978 58100 8988
rect 58380 8260 58436 8988
rect 58492 8978 58548 8988
rect 57932 8036 57988 8046
rect 57932 7476 57988 7980
rect 58380 8036 58436 8204
rect 58380 7970 58436 7980
rect 58044 7476 58100 7486
rect 57932 7420 58044 7476
rect 58044 7410 58100 7420
rect 57428 7308 57652 7364
rect 57820 7364 57876 7374
rect 58380 7364 58436 7374
rect 57820 7362 57988 7364
rect 57820 7310 57822 7362
rect 57874 7310 57988 7362
rect 57820 7308 57988 7310
rect 57372 7270 57428 7308
rect 57820 7298 57876 7308
rect 57932 7250 57988 7308
rect 58268 7308 58380 7364
rect 57932 7198 57934 7250
rect 57986 7198 57988 7250
rect 57820 6692 57876 6702
rect 57372 6468 57428 6478
rect 57372 6374 57428 6412
rect 57820 6466 57876 6636
rect 57820 6414 57822 6466
rect 57874 6414 57876 6466
rect 57820 6356 57876 6414
rect 57596 6300 57876 6356
rect 57932 6356 57988 7198
rect 57596 5796 57652 6300
rect 57932 6290 57988 6300
rect 58044 7252 58100 7262
rect 58044 6132 58100 7196
rect 57820 6076 58100 6132
rect 58156 6580 58212 6590
rect 57708 6020 57764 6030
rect 57708 5926 57764 5964
rect 57820 6018 57876 6076
rect 57820 5966 57822 6018
rect 57874 5966 57876 6018
rect 57596 5730 57652 5740
rect 57596 5236 57652 5246
rect 57596 5142 57652 5180
rect 56700 4162 56756 4172
rect 56924 4396 57316 4452
rect 57708 4900 57764 4910
rect 57708 4450 57764 4844
rect 57708 4398 57710 4450
rect 57762 4398 57764 4450
rect 56924 3554 56980 4396
rect 57708 4386 57764 4398
rect 56924 3502 56926 3554
rect 56978 3502 56980 3554
rect 56588 3330 56644 3342
rect 56588 3278 56590 3330
rect 56642 3278 56644 3330
rect 56588 1316 56644 3278
rect 56812 3332 56868 3342
rect 56812 3238 56868 3276
rect 56588 1250 56644 1260
rect 56924 980 56980 3502
rect 57484 4004 57540 4014
rect 57484 3554 57540 3948
rect 57820 4004 57876 5966
rect 58156 6020 58212 6524
rect 58156 5954 58212 5964
rect 58044 5906 58100 5918
rect 58044 5854 58046 5906
rect 58098 5854 58100 5906
rect 58044 5796 58100 5854
rect 58044 5730 58100 5740
rect 58268 5124 58324 7308
rect 58380 7270 58436 7308
rect 58716 7362 58772 20524
rect 59172 20412 59436 20422
rect 59228 20356 59276 20412
rect 59332 20356 59380 20412
rect 59172 20346 59436 20356
rect 59612 20018 59668 20860
rect 59836 20802 59892 20814
rect 59836 20750 59838 20802
rect 59890 20750 59892 20802
rect 59836 20242 59892 20750
rect 59836 20190 59838 20242
rect 59890 20190 59892 20242
rect 59836 20178 59892 20190
rect 59612 19966 59614 20018
rect 59666 19966 59668 20018
rect 59612 19954 59668 19966
rect 59948 20020 60004 21422
rect 59948 19954 60004 19964
rect 60060 21700 60116 21710
rect 60060 20804 60116 21644
rect 60060 20130 60116 20748
rect 60060 20078 60062 20130
rect 60114 20078 60116 20130
rect 60060 19458 60116 20078
rect 60060 19406 60062 19458
rect 60114 19406 60116 19458
rect 60060 19394 60116 19406
rect 60172 20018 60228 20030
rect 60172 19966 60174 20018
rect 60226 19966 60228 20018
rect 59724 19346 59780 19358
rect 59724 19294 59726 19346
rect 59778 19294 59780 19346
rect 59388 19236 59444 19246
rect 59388 19142 59444 19180
rect 59172 18844 59436 18854
rect 58940 18788 58996 18798
rect 59228 18788 59276 18844
rect 59332 18788 59380 18844
rect 59172 18778 59436 18788
rect 58940 18562 58996 18732
rect 58940 18510 58942 18562
rect 58994 18510 58996 18562
rect 58940 18498 58996 18510
rect 59164 18676 59220 18686
rect 59164 18562 59220 18620
rect 59388 18676 59444 18686
rect 59388 18582 59444 18620
rect 59164 18510 59166 18562
rect 59218 18510 59220 18562
rect 59164 18498 59220 18510
rect 59724 18452 59780 19294
rect 60172 19236 60228 19966
rect 60172 18676 60228 19180
rect 60172 18610 60228 18620
rect 60284 18452 60340 22092
rect 60508 21698 60564 21710
rect 60508 21646 60510 21698
rect 60562 21646 60564 21698
rect 60508 21476 60564 21646
rect 60732 21588 60788 21598
rect 60508 21410 60564 21420
rect 60620 21586 60788 21588
rect 60620 21534 60734 21586
rect 60786 21534 60788 21586
rect 60620 21532 60788 21534
rect 60396 20804 60452 20814
rect 60396 20710 60452 20748
rect 60620 20802 60676 21532
rect 60732 21522 60788 21532
rect 60620 20750 60622 20802
rect 60674 20750 60676 20802
rect 60620 20738 60676 20750
rect 59724 18358 59780 18396
rect 60172 18396 60340 18452
rect 59500 18226 59556 18238
rect 59500 18174 59502 18226
rect 59554 18174 59556 18226
rect 59500 17556 59556 18174
rect 59172 17276 59436 17286
rect 59228 17220 59276 17276
rect 59332 17220 59380 17276
rect 59172 17210 59436 17220
rect 59500 16322 59556 17500
rect 59500 16270 59502 16322
rect 59554 16270 59556 16322
rect 59500 16258 59556 16270
rect 59836 16210 59892 16222
rect 59836 16158 59838 16210
rect 59890 16158 59892 16210
rect 59172 15708 59436 15718
rect 59228 15652 59276 15708
rect 59332 15652 59380 15708
rect 59172 15642 59436 15652
rect 59836 15316 59892 16158
rect 59948 16100 60004 16110
rect 59948 16006 60004 16044
rect 60060 15316 60116 15326
rect 59836 15314 60116 15316
rect 59836 15262 60062 15314
rect 60114 15262 60116 15314
rect 59836 15260 60116 15262
rect 59836 15148 59892 15260
rect 60060 15250 60116 15260
rect 59612 15092 59892 15148
rect 59612 14642 59668 15092
rect 59612 14590 59614 14642
rect 59666 14590 59668 14642
rect 59612 14578 59668 14590
rect 60060 14530 60116 14542
rect 60060 14478 60062 14530
rect 60114 14478 60116 14530
rect 59172 14140 59436 14150
rect 59228 14084 59276 14140
rect 59332 14084 59380 14140
rect 59172 14074 59436 14084
rect 59276 13860 59332 13870
rect 59276 13074 59332 13804
rect 60060 13860 60116 14478
rect 60060 13794 60116 13804
rect 59836 13746 59892 13758
rect 59836 13694 59838 13746
rect 59890 13694 59892 13746
rect 59276 13022 59278 13074
rect 59330 13022 59332 13074
rect 59276 13010 59332 13022
rect 59388 13634 59444 13646
rect 59388 13582 59390 13634
rect 59442 13582 59444 13634
rect 59388 12852 59444 13582
rect 59836 13524 59892 13694
rect 59836 13458 59892 13468
rect 60172 13188 60228 18396
rect 60732 18228 60788 18238
rect 60396 17556 60452 17566
rect 60284 17108 60340 17118
rect 60284 17014 60340 17052
rect 60396 16548 60452 17500
rect 60284 16492 60452 16548
rect 60732 17108 60788 18172
rect 60284 15538 60340 16492
rect 60620 16212 60676 16222
rect 60732 16212 60788 17052
rect 60620 16210 60788 16212
rect 60620 16158 60622 16210
rect 60674 16158 60788 16210
rect 60620 16156 60788 16158
rect 60620 16146 60676 16156
rect 60284 15486 60286 15538
rect 60338 15486 60340 15538
rect 60284 15474 60340 15486
rect 60396 16100 60452 16110
rect 60396 15316 60452 16044
rect 60844 15988 60900 23660
rect 60956 21476 61012 31164
rect 61404 31108 61460 32732
rect 61516 32564 61572 32574
rect 61516 32470 61572 32508
rect 61628 32452 61684 32462
rect 61516 31780 61572 31790
rect 61628 31780 61684 32396
rect 61740 32450 61796 32732
rect 63532 32722 63588 32732
rect 62188 32564 62244 32574
rect 62188 32470 62244 32508
rect 63196 32564 63252 32574
rect 61740 32398 61742 32450
rect 61794 32398 61796 32450
rect 61740 32386 61796 32398
rect 62636 32452 62692 32462
rect 62636 32358 62692 32396
rect 61740 31892 62020 31948
rect 61740 31890 61796 31892
rect 61740 31838 61742 31890
rect 61794 31838 61796 31890
rect 61740 31826 61796 31838
rect 61516 31778 61684 31780
rect 61516 31726 61518 31778
rect 61570 31726 61684 31778
rect 61516 31724 61684 31726
rect 61516 31714 61572 31724
rect 61404 31052 61572 31108
rect 61068 30996 61124 31006
rect 61068 30994 61460 30996
rect 61068 30942 61070 30994
rect 61122 30942 61460 30994
rect 61068 30940 61460 30942
rect 61068 30930 61124 30940
rect 61404 30322 61460 30940
rect 61404 30270 61406 30322
rect 61458 30270 61460 30322
rect 61404 30258 61460 30270
rect 61404 28532 61460 28542
rect 61404 28438 61460 28476
rect 61516 28530 61572 31052
rect 61628 30994 61684 31724
rect 61852 31780 61908 31818
rect 61852 31714 61908 31724
rect 61852 31556 61908 31566
rect 61628 30942 61630 30994
rect 61682 30942 61684 30994
rect 61628 29540 61684 30942
rect 61740 31554 61908 31556
rect 61740 31502 61854 31554
rect 61906 31502 61908 31554
rect 61740 31500 61908 31502
rect 61740 30322 61796 31500
rect 61852 31490 61908 31500
rect 61964 30882 62020 31892
rect 61964 30830 61966 30882
rect 62018 30830 62020 30882
rect 61964 30660 62020 30830
rect 62300 31780 62356 31790
rect 63196 31780 63252 32508
rect 63532 32562 63588 32574
rect 63532 32510 63534 32562
rect 63586 32510 63588 32562
rect 63308 31780 63364 31790
rect 63196 31778 63364 31780
rect 63196 31726 63310 31778
rect 63362 31726 63364 31778
rect 63196 31724 63364 31726
rect 62300 30884 62356 31724
rect 63308 31714 63364 31724
rect 62188 30772 62244 30782
rect 62300 30772 62356 30828
rect 62188 30770 62356 30772
rect 62188 30718 62190 30770
rect 62242 30718 62356 30770
rect 62188 30716 62356 30718
rect 62188 30706 62244 30716
rect 61964 30594 62020 30604
rect 61740 30270 61742 30322
rect 61794 30270 61796 30322
rect 61740 30258 61796 30270
rect 62076 30212 62132 30222
rect 62076 30118 62132 30156
rect 61628 29474 61684 29484
rect 61516 28478 61518 28530
rect 61570 28478 61572 28530
rect 61516 28466 61572 28478
rect 61964 28642 62020 28654
rect 61964 28590 61966 28642
rect 62018 28590 62020 28642
rect 61628 28420 61684 28430
rect 61628 28326 61684 28364
rect 61964 28082 62020 28590
rect 61964 28030 61966 28082
rect 62018 28030 62020 28082
rect 61964 28018 62020 28030
rect 61404 27972 61460 27982
rect 61404 27878 61460 27916
rect 61852 27970 61908 27982
rect 61852 27918 61854 27970
rect 61906 27918 61908 27970
rect 61628 27858 61684 27870
rect 61628 27806 61630 27858
rect 61682 27806 61684 27858
rect 61180 27636 61236 27646
rect 61628 27636 61684 27806
rect 61852 27860 61908 27918
rect 61852 27794 61908 27804
rect 61180 27634 61684 27636
rect 61180 27582 61182 27634
rect 61234 27582 61684 27634
rect 61180 27580 61684 27582
rect 61180 27570 61236 27580
rect 61292 26964 61348 26974
rect 61180 26404 61236 26414
rect 61180 25620 61236 26348
rect 61292 26290 61348 26908
rect 61628 26964 61684 26974
rect 61628 26870 61684 26908
rect 61740 26850 61796 26862
rect 61740 26798 61742 26850
rect 61794 26798 61796 26850
rect 61292 26238 61294 26290
rect 61346 26238 61348 26290
rect 61292 26226 61348 26238
rect 61516 26292 61572 26302
rect 61740 26292 61796 26798
rect 61964 26852 62020 26862
rect 61964 26758 62020 26796
rect 61516 26290 61796 26292
rect 61516 26238 61518 26290
rect 61570 26238 61796 26290
rect 61516 26236 61796 26238
rect 62188 26292 62244 26302
rect 61292 25620 61348 25630
rect 61180 25618 61348 25620
rect 61180 25566 61294 25618
rect 61346 25566 61348 25618
rect 61180 25564 61348 25566
rect 61292 25508 61348 25564
rect 61516 25620 61572 26236
rect 62188 26198 62244 26236
rect 61516 25554 61572 25564
rect 61292 25442 61348 25452
rect 62188 25396 62244 25406
rect 62188 25302 62244 25340
rect 61852 24722 61908 24734
rect 61852 24670 61854 24722
rect 61906 24670 61908 24722
rect 61740 24610 61796 24622
rect 61740 24558 61742 24610
rect 61794 24558 61796 24610
rect 61740 23940 61796 24558
rect 61740 23846 61796 23884
rect 61852 23714 61908 24670
rect 62076 23940 62132 23950
rect 62076 23846 62132 23884
rect 61852 23662 61854 23714
rect 61906 23662 61908 23714
rect 61852 23604 61908 23662
rect 61852 23538 61908 23548
rect 61292 23380 61348 23390
rect 61292 23042 61348 23324
rect 61292 22990 61294 23042
rect 61346 22990 61348 23042
rect 61292 22978 61348 22990
rect 61404 23154 61460 23166
rect 61404 23102 61406 23154
rect 61458 23102 61460 23154
rect 61292 22148 61348 22158
rect 61404 22148 61460 23102
rect 61292 22146 61460 22148
rect 61292 22094 61294 22146
rect 61346 22094 61460 22146
rect 61292 22092 61460 22094
rect 61292 22036 61348 22092
rect 61292 21970 61348 21980
rect 61516 21700 61572 21710
rect 61516 21606 61572 21644
rect 61292 21588 61348 21598
rect 61292 21494 61348 21532
rect 61628 21586 61684 21598
rect 61628 21534 61630 21586
rect 61682 21534 61684 21586
rect 60956 21410 61012 21420
rect 61628 20804 61684 21534
rect 61628 19906 61684 20748
rect 61740 21588 61796 21598
rect 61740 20802 61796 21532
rect 62300 21026 62356 30716
rect 62524 31666 62580 31678
rect 62524 31614 62526 31666
rect 62578 31614 62580 31666
rect 62524 30212 62580 31614
rect 62636 31554 62692 31566
rect 62636 31502 62638 31554
rect 62690 31502 62692 31554
rect 62636 30996 62692 31502
rect 63532 31332 63588 32510
rect 63756 32562 63812 32574
rect 63756 32510 63758 32562
rect 63810 32510 63812 32562
rect 63756 31948 63812 32510
rect 63644 31892 63812 31948
rect 63644 31556 63700 31892
rect 63868 31890 63924 33182
rect 63980 33236 64036 33246
rect 63980 33142 64036 33180
rect 65660 33234 65716 33246
rect 65660 33182 65662 33234
rect 65714 33182 65716 33234
rect 65660 32676 65716 33182
rect 65660 32610 65716 32620
rect 63868 31838 63870 31890
rect 63922 31838 63924 31890
rect 63868 31826 63924 31838
rect 65884 31892 65940 36204
rect 67452 36036 67508 37100
rect 67452 35922 67508 35980
rect 67452 35870 67454 35922
rect 67506 35870 67508 35922
rect 67452 35858 67508 35870
rect 67564 36482 67620 36494
rect 67564 36430 67566 36482
rect 67618 36430 67620 36482
rect 66220 35700 66276 35710
rect 66220 35026 66276 35644
rect 66556 35700 66612 35710
rect 67116 35700 67172 35710
rect 66556 35698 67172 35700
rect 66556 35646 66558 35698
rect 66610 35646 67118 35698
rect 67170 35646 67172 35698
rect 66556 35644 67172 35646
rect 66556 35634 66612 35644
rect 67116 35634 67172 35644
rect 67564 35588 67620 36430
rect 67900 36260 67956 36270
rect 67900 35922 67956 36204
rect 67900 35870 67902 35922
rect 67954 35870 67956 35922
rect 67900 35858 67956 35870
rect 67564 35522 67620 35532
rect 68348 35588 68404 35598
rect 68348 35494 68404 35532
rect 66220 34974 66222 35026
rect 66274 34974 66276 35026
rect 66220 34962 66276 34974
rect 66668 35476 66724 35486
rect 65996 34914 66052 34926
rect 65996 34862 65998 34914
rect 66050 34862 66052 34914
rect 65996 34692 66052 34862
rect 66668 34914 66724 35420
rect 66668 34862 66670 34914
rect 66722 34862 66724 34914
rect 66668 34850 66724 34862
rect 67116 34916 67172 34926
rect 65996 34626 66052 34636
rect 66444 34802 66500 34814
rect 66444 34750 66446 34802
rect 66498 34750 66500 34802
rect 66444 34580 66500 34750
rect 65996 34132 66052 34142
rect 65996 34038 66052 34076
rect 66444 34132 66500 34524
rect 67116 34690 67172 34860
rect 67116 34638 67118 34690
rect 67170 34638 67172 34690
rect 66444 34066 66500 34076
rect 66668 34132 66724 34142
rect 66556 33348 66612 33358
rect 66444 33292 66556 33348
rect 66444 32674 66500 33292
rect 66556 33254 66612 33292
rect 66444 32622 66446 32674
rect 66498 32622 66500 32674
rect 66444 32610 66500 32622
rect 66668 32450 66724 34076
rect 67116 33908 67172 34638
rect 67116 33842 67172 33852
rect 67116 33346 67172 33358
rect 67116 33294 67118 33346
rect 67170 33294 67172 33346
rect 67116 32788 67172 33294
rect 68460 33348 68516 37884
rect 68572 36594 68628 38108
rect 70476 37044 70532 37054
rect 68832 36876 69096 36886
rect 68888 36820 68936 36876
rect 68992 36820 69040 36876
rect 68832 36810 69096 36820
rect 68572 36542 68574 36594
rect 68626 36542 68628 36594
rect 68572 36530 68628 36542
rect 69468 36484 69524 36494
rect 69244 36482 69524 36484
rect 69244 36430 69470 36482
rect 69522 36430 69524 36482
rect 69244 36428 69524 36430
rect 68684 36372 68740 36382
rect 68684 34916 68740 36316
rect 69020 35588 69076 35598
rect 69244 35588 69300 36428
rect 69468 36418 69524 36428
rect 70476 36372 70532 36988
rect 70700 36594 70756 39200
rect 70700 36542 70702 36594
rect 70754 36542 70756 36594
rect 70700 36530 70756 36542
rect 71148 37828 71204 37838
rect 70476 35922 70532 36316
rect 71148 36148 71204 37772
rect 71708 36708 71764 36718
rect 71148 36082 71204 36092
rect 71372 36482 71428 36494
rect 71372 36430 71374 36482
rect 71426 36430 71428 36482
rect 70476 35870 70478 35922
rect 70530 35870 70532 35922
rect 70476 35858 70532 35870
rect 70812 35698 70868 35710
rect 70812 35646 70814 35698
rect 70866 35646 70868 35698
rect 69020 35586 69300 35588
rect 69020 35534 69022 35586
rect 69074 35534 69300 35586
rect 69020 35532 69300 35534
rect 69020 35522 69076 35532
rect 68832 35308 69096 35318
rect 68888 35252 68936 35308
rect 68992 35252 69040 35308
rect 68832 35242 69096 35252
rect 68684 34850 68740 34860
rect 68832 33740 69096 33750
rect 68888 33684 68936 33740
rect 68992 33684 69040 33740
rect 68832 33674 69096 33684
rect 68460 33282 68516 33292
rect 67228 33234 67284 33246
rect 67228 33182 67230 33234
rect 67282 33182 67284 33234
rect 67228 33124 67284 33182
rect 69244 33236 69300 35532
rect 69468 35588 69524 35598
rect 69468 35252 69524 35532
rect 69692 35586 69748 35598
rect 69692 35534 69694 35586
rect 69746 35534 69748 35586
rect 69580 35476 69636 35486
rect 69580 35382 69636 35420
rect 69468 35196 69636 35252
rect 69468 35026 69524 35038
rect 69468 34974 69470 35026
rect 69522 34974 69524 35026
rect 69468 34804 69524 34974
rect 69468 34738 69524 34748
rect 69244 33170 69300 33180
rect 69580 33572 69636 35196
rect 69692 35028 69748 35534
rect 69692 34962 69748 34972
rect 69692 34802 69748 34814
rect 69692 34750 69694 34802
rect 69746 34750 69748 34802
rect 69692 34580 69748 34750
rect 70812 34692 70868 35646
rect 71260 35588 71316 35598
rect 71372 35588 71428 36430
rect 71708 35922 71764 36652
rect 73164 36596 73220 39200
rect 75628 39060 75684 39200
rect 75964 39060 76020 39228
rect 75628 39004 76020 39060
rect 75404 38052 75460 38062
rect 73164 36530 73220 36540
rect 73500 37268 73556 37278
rect 73388 36482 73444 36494
rect 73388 36430 73390 36482
rect 73442 36430 73444 36482
rect 72492 36370 72548 36382
rect 72492 36318 72494 36370
rect 72546 36318 72548 36370
rect 72492 35924 72548 36318
rect 73164 36372 73220 36382
rect 72828 36260 72884 36270
rect 72828 36166 72884 36204
rect 71708 35870 71710 35922
rect 71762 35870 71764 35922
rect 71708 35812 71764 35870
rect 72380 35868 72492 35924
rect 71708 35746 71764 35756
rect 72268 35812 72324 35822
rect 72268 35718 72324 35756
rect 71260 35586 71540 35588
rect 71260 35534 71262 35586
rect 71314 35534 71540 35586
rect 71260 35532 71540 35534
rect 71260 35522 71316 35532
rect 71372 34804 71428 34814
rect 71372 34710 71428 34748
rect 71260 34692 71316 34702
rect 70812 34690 71316 34692
rect 70812 34638 71262 34690
rect 71314 34638 71316 34690
rect 70812 34636 71316 34638
rect 71260 34626 71316 34636
rect 69692 34514 69748 34524
rect 70140 34356 70196 34366
rect 70140 34354 70532 34356
rect 70140 34302 70142 34354
rect 70194 34302 70532 34354
rect 70140 34300 70532 34302
rect 70140 34290 70196 34300
rect 70252 34130 70308 34142
rect 70252 34078 70254 34130
rect 70306 34078 70308 34130
rect 70140 33908 70196 33918
rect 70140 33814 70196 33852
rect 67228 33058 67284 33068
rect 67228 32788 67284 32798
rect 67116 32786 67284 32788
rect 67116 32734 67230 32786
rect 67282 32734 67284 32786
rect 67116 32732 67284 32734
rect 67228 32722 67284 32732
rect 69580 32786 69636 33516
rect 69580 32734 69582 32786
rect 69634 32734 69636 32786
rect 69580 32722 69636 32734
rect 70252 33346 70308 34078
rect 70252 33294 70254 33346
rect 70306 33294 70308 33346
rect 67452 32676 67508 32686
rect 66780 32564 66836 32602
rect 67452 32582 67508 32620
rect 69356 32676 69412 32686
rect 66780 32498 66836 32508
rect 67564 32564 67620 32574
rect 67564 32470 67620 32508
rect 66668 32398 66670 32450
rect 66722 32398 66724 32450
rect 66668 32386 66724 32398
rect 68832 32172 69096 32182
rect 68888 32116 68936 32172
rect 68992 32116 69040 32172
rect 68832 32106 69096 32116
rect 65884 31760 65940 31836
rect 67564 31780 67620 31790
rect 65996 31666 66052 31678
rect 65996 31614 65998 31666
rect 66050 31614 66052 31666
rect 63868 31556 63924 31566
rect 63644 31462 63700 31500
rect 63756 31554 63924 31556
rect 63756 31502 63870 31554
rect 63922 31502 63924 31554
rect 63756 31500 63924 31502
rect 63756 31332 63812 31500
rect 63868 31490 63924 31500
rect 64316 31554 64372 31566
rect 64316 31502 64318 31554
rect 64370 31502 64372 31554
rect 63532 31276 63812 31332
rect 63196 30996 63252 31006
rect 62636 30994 63252 30996
rect 62636 30942 63198 30994
rect 63250 30942 63252 30994
rect 62636 30940 63252 30942
rect 63196 30930 63252 30940
rect 63308 30772 63364 30782
rect 63308 30678 63364 30716
rect 62524 30146 62580 30156
rect 63644 29652 63700 29662
rect 63756 29652 63812 31276
rect 63868 30884 63924 30894
rect 63868 30790 63924 30828
rect 64316 30884 64372 31502
rect 64316 30818 64372 30828
rect 65436 31556 65492 31566
rect 63644 29650 63812 29652
rect 63644 29598 63646 29650
rect 63698 29598 63812 29650
rect 63644 29596 63812 29598
rect 63644 29586 63700 29596
rect 63868 29538 63924 29550
rect 63868 29486 63870 29538
rect 63922 29486 63924 29538
rect 63868 28868 63924 29486
rect 63980 29428 64036 29438
rect 64540 29428 64596 29438
rect 63980 29426 64596 29428
rect 63980 29374 63982 29426
rect 64034 29374 64542 29426
rect 64594 29374 64596 29426
rect 63980 29372 64596 29374
rect 63980 29362 64036 29372
rect 64540 29362 64596 29372
rect 64652 29316 64708 29326
rect 64652 29314 65156 29316
rect 64652 29262 64654 29314
rect 64706 29262 65156 29314
rect 64652 29260 65156 29262
rect 64652 29250 64708 29260
rect 62860 27970 62916 27982
rect 62860 27918 62862 27970
rect 62914 27918 62916 27970
rect 62636 27860 62692 27870
rect 62412 25508 62468 25518
rect 62412 25414 62468 25452
rect 62636 25508 62692 27804
rect 62748 27858 62804 27870
rect 62748 27806 62750 27858
rect 62802 27806 62804 27858
rect 62748 26292 62804 27806
rect 62860 27300 62916 27918
rect 63084 27858 63140 27870
rect 63084 27806 63086 27858
rect 63138 27806 63140 27858
rect 62972 27300 63028 27310
rect 62860 27298 63028 27300
rect 62860 27246 62974 27298
rect 63026 27246 63028 27298
rect 62860 27244 63028 27246
rect 62860 26292 62916 26302
rect 62748 26236 62860 26292
rect 62972 26292 63028 27244
rect 63084 27076 63140 27806
rect 63868 27300 63924 28812
rect 65100 28756 65156 29260
rect 64204 28642 64260 28654
rect 64204 28590 64206 28642
rect 64258 28590 64260 28642
rect 64204 27972 64260 28590
rect 64204 27906 64260 27916
rect 64652 28642 64708 28654
rect 64652 28590 64654 28642
rect 64706 28590 64708 28642
rect 65100 28624 65156 28700
rect 64428 27748 64484 27758
rect 63980 27300 64036 27310
rect 63868 27298 64036 27300
rect 63868 27246 63982 27298
rect 64034 27246 64036 27298
rect 63868 27244 64036 27246
rect 63980 27234 64036 27244
rect 63084 27010 63140 27020
rect 63868 27076 63924 27086
rect 63868 26982 63924 27020
rect 63308 26962 63364 26974
rect 63308 26910 63310 26962
rect 63362 26910 63364 26962
rect 63084 26852 63140 26862
rect 63084 26850 63252 26852
rect 63084 26798 63086 26850
rect 63138 26798 63252 26850
rect 63084 26796 63252 26798
rect 63084 26786 63140 26796
rect 63084 26292 63140 26302
rect 62972 26290 63140 26292
rect 62972 26238 63086 26290
rect 63138 26238 63140 26290
rect 62972 26236 63140 26238
rect 62860 26198 62916 26236
rect 63084 26226 63140 26236
rect 63196 26068 63252 26796
rect 63308 26516 63364 26910
rect 63308 26450 63364 26460
rect 63756 26964 63812 26974
rect 63756 26402 63812 26908
rect 63980 26852 64036 26862
rect 63980 26758 64036 26796
rect 63756 26350 63758 26402
rect 63810 26350 63812 26402
rect 63756 26338 63812 26350
rect 62748 26012 63252 26068
rect 62748 25618 62804 26012
rect 62748 25566 62750 25618
rect 62802 25566 62804 25618
rect 62748 25554 62804 25566
rect 62860 25732 62916 25742
rect 62636 25376 62692 25452
rect 62860 25506 62916 25676
rect 64204 25620 64260 25630
rect 64204 25526 64260 25564
rect 62860 25454 62862 25506
rect 62914 25454 62916 25506
rect 62860 25442 62916 25454
rect 63308 25508 63364 25518
rect 63084 25284 63140 25294
rect 62412 24836 62468 24846
rect 62412 24742 62468 24780
rect 62748 23156 62804 23166
rect 62748 23062 62804 23100
rect 63084 21588 63140 25228
rect 63308 24948 63364 25452
rect 63868 25396 63924 25406
rect 63868 25302 63924 25340
rect 63980 25172 64036 25182
rect 63420 24948 63476 24958
rect 63308 24892 63420 24948
rect 63196 21812 63252 21822
rect 63308 21812 63364 24892
rect 63420 24816 63476 24892
rect 63868 24610 63924 24622
rect 63868 24558 63870 24610
rect 63922 24558 63924 24610
rect 63868 24498 63924 24558
rect 63868 24446 63870 24498
rect 63922 24446 63924 24498
rect 63532 23042 63588 23054
rect 63532 22990 63534 23042
rect 63586 22990 63588 23042
rect 63532 22596 63588 22990
rect 63532 22530 63588 22540
rect 63756 22260 63812 22270
rect 63756 22166 63812 22204
rect 63196 21810 63364 21812
rect 63196 21758 63198 21810
rect 63250 21758 63364 21810
rect 63196 21756 63364 21758
rect 63196 21746 63252 21756
rect 63308 21700 63364 21756
rect 63756 21812 63812 21822
rect 63756 21718 63812 21756
rect 63308 21634 63364 21644
rect 63084 21532 63252 21588
rect 62300 20974 62302 21026
rect 62354 20974 62356 21026
rect 62300 20962 62356 20974
rect 61740 20750 61742 20802
rect 61794 20750 61796 20802
rect 61740 20738 61796 20750
rect 61852 20804 61908 20814
rect 61628 19854 61630 19906
rect 61682 19854 61684 19906
rect 61628 19842 61684 19854
rect 61852 19458 61908 20748
rect 61964 20802 62020 20814
rect 61964 20750 61966 20802
rect 62018 20750 62020 20802
rect 61964 20692 62020 20750
rect 62972 20804 63028 20814
rect 62972 20710 63028 20748
rect 61964 20626 62020 20636
rect 63196 20188 63252 21532
rect 63868 21364 63924 24446
rect 63980 21588 64036 25116
rect 64428 24834 64484 27692
rect 64652 27412 64708 28590
rect 65436 28082 65492 31500
rect 65772 31556 65828 31566
rect 65772 31462 65828 31500
rect 65996 31332 66052 31614
rect 66780 31666 66836 31678
rect 66780 31614 66782 31666
rect 66834 31614 66836 31666
rect 65548 31276 66052 31332
rect 66668 31554 66724 31566
rect 66668 31502 66670 31554
rect 66722 31502 66724 31554
rect 65548 31218 65604 31276
rect 66668 31220 66724 31502
rect 66780 31444 66836 31614
rect 66780 31378 66836 31388
rect 67228 31554 67284 31566
rect 67228 31502 67230 31554
rect 67282 31502 67284 31554
rect 67228 31444 67284 31502
rect 67228 31378 67284 31388
rect 67340 31556 67396 31566
rect 65548 31166 65550 31218
rect 65602 31166 65604 31218
rect 65548 31154 65604 31166
rect 65996 31164 66948 31220
rect 65996 31106 66052 31164
rect 65996 31054 65998 31106
rect 66050 31054 66052 31106
rect 65996 31042 66052 31054
rect 66892 31106 66948 31164
rect 67340 31218 67396 31500
rect 67340 31166 67342 31218
rect 67394 31166 67396 31218
rect 67340 31154 67396 31166
rect 66892 31054 66894 31106
rect 66946 31054 66948 31106
rect 66892 31042 66948 31054
rect 66108 30996 66164 31006
rect 66108 30772 66164 30940
rect 66332 30994 66388 31006
rect 66332 30942 66334 30994
rect 66386 30942 66388 30994
rect 66332 30884 66388 30942
rect 67116 30994 67172 31006
rect 67116 30942 67118 30994
rect 67170 30942 67172 30994
rect 67116 30884 67172 30942
rect 66332 30828 67172 30884
rect 67564 30996 67620 31724
rect 68236 31668 68292 31678
rect 68236 31218 68292 31612
rect 68572 31556 68628 31566
rect 68236 31166 68238 31218
rect 68290 31166 68292 31218
rect 68236 31154 68292 31166
rect 68460 31554 68628 31556
rect 68460 31502 68574 31554
rect 68626 31502 68628 31554
rect 68460 31500 68628 31502
rect 68460 31444 68516 31500
rect 68572 31490 68628 31500
rect 67564 30864 67620 30940
rect 68460 31106 68516 31388
rect 68460 31054 68462 31106
rect 68514 31054 68516 31106
rect 66108 30706 66164 30716
rect 67004 30322 67060 30334
rect 67004 30270 67006 30322
rect 67058 30270 67060 30322
rect 66108 30212 66164 30222
rect 66108 30118 66164 30156
rect 66780 30210 66836 30222
rect 66780 30158 66782 30210
rect 66834 30158 66836 30210
rect 66780 29316 66836 30158
rect 67004 29988 67060 30270
rect 67116 30212 67172 30828
rect 68460 30324 68516 31054
rect 68572 30996 68628 31006
rect 68572 30902 68628 30940
rect 69132 30996 69188 31006
rect 69132 30902 69188 30940
rect 68832 30604 69096 30614
rect 68888 30548 68936 30604
rect 68992 30548 69040 30604
rect 68832 30538 69096 30548
rect 68460 30258 68516 30268
rect 67564 30212 67620 30222
rect 67116 30210 67620 30212
rect 67116 30158 67566 30210
rect 67618 30158 67620 30210
rect 67116 30156 67620 30158
rect 67564 30146 67620 30156
rect 67788 30100 67844 30110
rect 67788 30006 67844 30044
rect 67900 30098 67956 30110
rect 67900 30046 67902 30098
rect 67954 30046 67956 30098
rect 67004 29922 67060 29932
rect 67900 29988 67956 30046
rect 68460 30100 68516 30110
rect 68460 30006 68516 30044
rect 68572 30098 68628 30110
rect 68572 30046 68574 30098
rect 68626 30046 68628 30098
rect 67788 29540 67844 29550
rect 67900 29540 67956 29932
rect 67788 29538 67900 29540
rect 67788 29486 67790 29538
rect 67842 29486 67900 29538
rect 67788 29484 67900 29486
rect 67788 29474 67844 29484
rect 67900 29474 67956 29484
rect 68236 29540 68292 29550
rect 68236 29446 68292 29484
rect 66780 29250 66836 29260
rect 67340 29316 67396 29326
rect 67340 29222 67396 29260
rect 68572 29316 68628 30046
rect 68796 29316 68852 29326
rect 68628 29314 68852 29316
rect 68628 29262 68798 29314
rect 68850 29262 68852 29314
rect 68628 29260 68852 29262
rect 68572 29184 68628 29260
rect 68796 29204 68852 29260
rect 68796 29148 69300 29204
rect 68832 29036 69096 29046
rect 68888 28980 68936 29036
rect 68992 28980 69040 29036
rect 68832 28970 69096 28980
rect 65996 28868 66052 28878
rect 65772 28756 65828 28766
rect 65772 28662 65828 28700
rect 65436 28030 65438 28082
rect 65490 28030 65492 28082
rect 65436 28018 65492 28030
rect 65884 28644 65940 28654
rect 65548 27972 65604 27982
rect 64652 27356 64932 27412
rect 64876 27300 64932 27356
rect 64876 27074 64932 27244
rect 64876 27022 64878 27074
rect 64930 27022 64932 27074
rect 64876 27010 64932 27022
rect 65212 26962 65268 26974
rect 65212 26910 65214 26962
rect 65266 26910 65268 26962
rect 65100 26850 65156 26862
rect 65100 26798 65102 26850
rect 65154 26798 65156 26850
rect 64652 26180 64708 26190
rect 65100 26180 65156 26798
rect 64540 26178 65156 26180
rect 64540 26126 64654 26178
rect 64706 26126 65156 26178
rect 64540 26124 65156 26126
rect 65212 26180 65268 26910
rect 65436 26516 65492 26526
rect 65436 26422 65492 26460
rect 65548 26402 65604 27916
rect 65772 27860 65828 27870
rect 65884 27860 65940 28588
rect 65996 28642 66052 28812
rect 65996 28590 65998 28642
rect 66050 28590 66052 28642
rect 65996 28578 66052 28590
rect 66668 28644 66724 28654
rect 66668 28530 66724 28588
rect 67340 28644 67396 28654
rect 67340 28550 67396 28588
rect 67564 28642 67620 28654
rect 67564 28590 67566 28642
rect 67618 28590 67620 28642
rect 66668 28478 66670 28530
rect 66722 28478 66724 28530
rect 66668 28466 66724 28478
rect 65996 27972 66052 27982
rect 65996 27878 66052 27916
rect 66332 27972 66388 27982
rect 65772 27858 65940 27860
rect 65772 27806 65774 27858
rect 65826 27806 65940 27858
rect 65772 27804 65940 27806
rect 65772 27794 65828 27804
rect 65996 27300 66052 27310
rect 65996 27206 66052 27244
rect 66332 27298 66388 27916
rect 67564 27972 67620 28590
rect 68236 28532 68292 28542
rect 68236 28438 68292 28476
rect 67564 27906 67620 27916
rect 69244 27524 69300 29148
rect 69356 28868 69412 32620
rect 69916 32562 69972 32574
rect 69916 32510 69918 32562
rect 69970 32510 69972 32562
rect 69916 31948 69972 32510
rect 70252 32002 70308 33294
rect 70476 33348 70532 34300
rect 71148 34244 71204 34254
rect 71148 34150 71204 34188
rect 71484 34244 71540 35532
rect 72268 35028 72324 35038
rect 71484 34178 71540 34188
rect 72156 34802 72212 34814
rect 72156 34750 72158 34802
rect 72210 34750 72212 34802
rect 70924 34132 70980 34142
rect 70924 34130 71092 34132
rect 70924 34078 70926 34130
rect 70978 34078 71092 34130
rect 70924 34076 71092 34078
rect 70924 34066 70980 34076
rect 71036 33460 71092 34076
rect 71820 34018 71876 34030
rect 71820 33966 71822 34018
rect 71874 33966 71876 34018
rect 71820 33908 71876 33966
rect 71820 33842 71876 33852
rect 72156 33908 72212 34750
rect 72156 33842 72212 33852
rect 72268 34802 72324 34972
rect 72268 34750 72270 34802
rect 72322 34750 72324 34802
rect 72268 33570 72324 34750
rect 72380 34354 72436 35868
rect 72492 35858 72548 35868
rect 72604 35812 72660 35822
rect 72604 35718 72660 35756
rect 72492 34804 72548 34814
rect 72492 34710 72548 34748
rect 72380 34302 72382 34354
rect 72434 34302 72436 34354
rect 72380 34290 72436 34302
rect 72268 33518 72270 33570
rect 72322 33518 72324 33570
rect 72268 33506 72324 33518
rect 71148 33460 71204 33470
rect 71036 33458 71204 33460
rect 71036 33406 71150 33458
rect 71202 33406 71204 33458
rect 71036 33404 71204 33406
rect 71148 33394 71204 33404
rect 73164 33458 73220 36316
rect 73388 36372 73444 36430
rect 73388 36306 73444 36316
rect 73276 36148 73332 36158
rect 73276 35922 73332 36092
rect 73276 35870 73278 35922
rect 73330 35870 73332 35922
rect 73276 34914 73332 35870
rect 73276 34862 73278 34914
rect 73330 34862 73332 34914
rect 73276 34850 73332 34862
rect 73500 34356 73556 37212
rect 74060 36596 74116 36606
rect 74060 36502 74116 36540
rect 75404 36596 75460 37996
rect 74172 36484 74228 36494
rect 74172 35698 74228 36428
rect 75404 36482 75460 36540
rect 76972 36594 77028 39228
rect 78064 39200 78176 40000
rect 77868 38500 77924 38510
rect 76972 36542 76974 36594
rect 77026 36542 77028 36594
rect 76972 36530 77028 36542
rect 77084 37380 77140 37390
rect 75404 36430 75406 36482
rect 75458 36430 75460 36482
rect 75404 36418 75460 36430
rect 76300 36482 76356 36494
rect 76300 36430 76302 36482
rect 76354 36430 76356 36482
rect 74956 36260 75012 36270
rect 74396 35812 74452 35822
rect 74396 35810 74564 35812
rect 74396 35758 74398 35810
rect 74450 35758 74564 35810
rect 74396 35756 74564 35758
rect 74396 35746 74452 35756
rect 74172 35646 74174 35698
rect 74226 35646 74228 35698
rect 74060 35028 74116 35038
rect 74172 35028 74228 35646
rect 74060 35026 74228 35028
rect 74060 34974 74062 35026
rect 74114 34974 74228 35026
rect 74060 34972 74228 34974
rect 74060 34962 74116 34972
rect 73948 34916 74004 34926
rect 73612 34692 73668 34702
rect 73612 34690 73780 34692
rect 73612 34638 73614 34690
rect 73666 34638 73780 34690
rect 73612 34636 73780 34638
rect 73612 34626 73668 34636
rect 73612 34356 73668 34366
rect 73500 34354 73668 34356
rect 73500 34302 73614 34354
rect 73666 34302 73668 34354
rect 73500 34300 73668 34302
rect 73612 34244 73668 34300
rect 73612 34178 73668 34188
rect 73164 33406 73166 33458
rect 73218 33406 73220 33458
rect 73164 33394 73220 33406
rect 70588 33348 70644 33358
rect 70476 33346 70644 33348
rect 70476 33294 70590 33346
rect 70642 33294 70644 33346
rect 70476 33292 70644 33294
rect 70476 32674 70532 33292
rect 70588 33282 70644 33292
rect 71932 33346 71988 33358
rect 71932 33294 71934 33346
rect 71986 33294 71988 33346
rect 71708 33236 71764 33246
rect 71148 33234 71764 33236
rect 71148 33182 71710 33234
rect 71762 33182 71764 33234
rect 71148 33180 71764 33182
rect 70476 32622 70478 32674
rect 70530 32622 70532 32674
rect 70476 32610 70532 32622
rect 70588 33124 70644 33134
rect 70588 32562 70644 33068
rect 70588 32510 70590 32562
rect 70642 32510 70644 32562
rect 70588 32498 70644 32510
rect 70700 32564 70756 32574
rect 70252 31950 70254 32002
rect 70306 31950 70308 32002
rect 69916 31892 70084 31948
rect 70252 31938 70308 31950
rect 69804 31780 69860 31790
rect 69804 31686 69860 31724
rect 69580 31668 69636 31678
rect 69580 31574 69636 31612
rect 70028 31444 70084 31892
rect 70028 31388 70308 31444
rect 69580 31220 69636 31230
rect 69580 31126 69636 31164
rect 70252 31106 70308 31388
rect 70700 31220 70756 32508
rect 71148 32562 71204 33180
rect 71148 32510 71150 32562
rect 71202 32510 71204 32562
rect 71148 32498 71204 32510
rect 70252 31054 70254 31106
rect 70306 31054 70308 31106
rect 70252 31042 70308 31054
rect 70588 31164 70756 31220
rect 70812 31778 70868 31790
rect 70812 31726 70814 31778
rect 70866 31726 70868 31778
rect 70812 31220 70868 31726
rect 71260 31668 71316 31678
rect 71260 31574 71316 31612
rect 69468 30994 69524 31006
rect 69468 30942 69470 30994
rect 69522 30942 69524 30994
rect 69468 30324 69524 30942
rect 69692 30996 69748 31006
rect 69692 30994 70196 30996
rect 69692 30942 69694 30994
rect 69746 30942 70196 30994
rect 69692 30940 70196 30942
rect 69692 30930 69748 30940
rect 70140 30434 70196 30940
rect 70140 30382 70142 30434
rect 70194 30382 70196 30434
rect 70140 30370 70196 30382
rect 69468 30258 69524 30268
rect 69468 30100 69524 30110
rect 69468 30006 69524 30044
rect 69580 30098 69636 30110
rect 69580 30046 69582 30098
rect 69634 30046 69636 30098
rect 69580 29540 69636 30046
rect 69692 30100 69748 30110
rect 69692 30006 69748 30044
rect 69580 29316 69636 29484
rect 70028 29316 70084 29326
rect 69580 29314 70084 29316
rect 69580 29262 70030 29314
rect 70082 29262 70084 29314
rect 69580 29260 70084 29262
rect 69468 28868 69524 28878
rect 69356 28866 69524 28868
rect 69356 28814 69470 28866
rect 69522 28814 69524 28866
rect 69356 28812 69524 28814
rect 69468 28802 69524 28812
rect 70028 28868 70084 29260
rect 70588 29204 70644 31164
rect 70812 31154 70868 31164
rect 71036 31556 71092 31566
rect 70700 30994 70756 31006
rect 70700 30942 70702 30994
rect 70754 30942 70756 30994
rect 70700 30434 70756 30942
rect 70700 30382 70702 30434
rect 70754 30382 70756 30434
rect 70700 30370 70756 30382
rect 71036 30434 71092 31500
rect 71036 30382 71038 30434
rect 71090 30382 71092 30434
rect 71036 30370 71092 30382
rect 71148 30882 71204 30894
rect 71148 30830 71150 30882
rect 71202 30830 71204 30882
rect 70812 30324 70868 30334
rect 70812 29988 70868 30268
rect 71148 30212 71204 30830
rect 71148 30146 71204 30156
rect 70812 29894 70868 29932
rect 70700 29652 70756 29662
rect 71596 29652 71652 33180
rect 71708 33170 71764 33180
rect 71932 33124 71988 33294
rect 71932 33058 71988 33068
rect 72380 33124 72436 33134
rect 72044 31668 72100 31678
rect 72044 31666 72212 31668
rect 72044 31614 72046 31666
rect 72098 31614 72212 31666
rect 72044 31612 72212 31614
rect 72044 31602 72100 31612
rect 71820 31556 71876 31566
rect 71820 31218 71876 31500
rect 71932 31554 71988 31566
rect 71932 31502 71934 31554
rect 71986 31502 71988 31554
rect 71932 31444 71988 31502
rect 71932 31378 71988 31388
rect 71820 31166 71822 31218
rect 71874 31166 71876 31218
rect 71820 31154 71876 31166
rect 71932 31220 71988 31230
rect 71932 31126 71988 31164
rect 71708 30996 71764 31006
rect 72044 30996 72100 31006
rect 71708 30434 71764 30940
rect 71932 30994 72100 30996
rect 71932 30942 72046 30994
rect 72098 30942 72100 30994
rect 71932 30940 72100 30942
rect 71932 30884 71988 30940
rect 72044 30930 72100 30940
rect 71708 30382 71710 30434
rect 71762 30382 71764 30434
rect 71708 30370 71764 30382
rect 71820 30828 71988 30884
rect 71820 29988 71876 30828
rect 72044 30772 72100 30782
rect 72044 30212 72100 30716
rect 71820 29764 71876 29932
rect 71820 29698 71876 29708
rect 71932 30210 72100 30212
rect 71932 30158 72046 30210
rect 72098 30158 72100 30210
rect 71932 30156 72100 30158
rect 71708 29652 71764 29662
rect 70700 29650 70980 29652
rect 70700 29598 70702 29650
rect 70754 29598 70980 29650
rect 70700 29596 70980 29598
rect 71596 29650 71764 29652
rect 71596 29598 71710 29650
rect 71762 29598 71764 29650
rect 71596 29596 71764 29598
rect 70700 29586 70756 29596
rect 70812 29428 70868 29438
rect 70700 29204 70756 29214
rect 70588 29202 70756 29204
rect 70588 29150 70702 29202
rect 70754 29150 70756 29202
rect 70588 29148 70756 29150
rect 70700 29138 70756 29148
rect 70028 28802 70084 28812
rect 70028 28644 70084 28654
rect 69468 28532 69524 28542
rect 69468 27858 69524 28476
rect 69468 27806 69470 27858
rect 69522 27806 69524 27858
rect 69468 27794 69524 27806
rect 69580 28530 69636 28542
rect 69580 28478 69582 28530
rect 69634 28478 69636 28530
rect 68832 27468 69096 27478
rect 68888 27412 68936 27468
rect 68992 27412 69040 27468
rect 69244 27458 69300 27468
rect 69580 27746 69636 28478
rect 70028 27970 70084 28588
rect 70812 28644 70868 29372
rect 70812 28578 70868 28588
rect 70028 27918 70030 27970
rect 70082 27918 70084 27970
rect 70028 27906 70084 27918
rect 70924 27972 70980 29596
rect 71708 29586 71764 29596
rect 71484 29540 71540 29550
rect 71484 29538 71652 29540
rect 71484 29486 71486 29538
rect 71538 29486 71652 29538
rect 71484 29484 71652 29486
rect 71484 29474 71540 29484
rect 71372 29428 71428 29438
rect 71372 29334 71428 29372
rect 71484 28754 71540 28766
rect 71484 28702 71486 28754
rect 71538 28702 71540 28754
rect 71036 28644 71092 28654
rect 71036 28550 71092 28588
rect 71484 28082 71540 28702
rect 71484 28030 71486 28082
rect 71538 28030 71540 28082
rect 71484 28018 71540 28030
rect 71372 27972 71428 27982
rect 70924 27970 71428 27972
rect 70924 27918 71374 27970
rect 71426 27918 71428 27970
rect 70924 27916 71428 27918
rect 69580 27694 69582 27746
rect 69634 27694 69636 27746
rect 68832 27402 69096 27412
rect 66332 27246 66334 27298
rect 66386 27246 66388 27298
rect 66332 27234 66388 27246
rect 68348 27076 68404 27086
rect 68348 26982 68404 27020
rect 69468 27076 69524 27086
rect 69468 26982 69524 27020
rect 65772 26964 65828 26974
rect 65772 26962 65940 26964
rect 65772 26910 65774 26962
rect 65826 26910 65940 26962
rect 65772 26908 65940 26910
rect 65772 26898 65828 26908
rect 65548 26350 65550 26402
rect 65602 26350 65604 26402
rect 65548 26338 65604 26350
rect 64540 24948 64596 26124
rect 64652 26114 64708 26124
rect 64540 24854 64596 24892
rect 64652 25732 64708 25742
rect 64652 25618 64708 25676
rect 64652 25566 64654 25618
rect 64706 25566 64708 25618
rect 64428 24782 64430 24834
rect 64482 24782 64484 24834
rect 64204 24500 64260 24510
rect 64428 24500 64484 24782
rect 64204 24498 64484 24500
rect 64204 24446 64206 24498
rect 64258 24446 64484 24498
rect 64204 24444 64484 24446
rect 64204 24434 64260 24444
rect 64428 24162 64484 24444
rect 64428 24110 64430 24162
rect 64482 24110 64484 24162
rect 64428 24098 64484 24110
rect 63980 21522 64036 21532
rect 64092 23604 64148 23614
rect 64092 23154 64148 23548
rect 64092 23102 64094 23154
rect 64146 23102 64148 23154
rect 63868 21308 64036 21364
rect 63420 20804 63476 20814
rect 63868 20804 63924 20814
rect 63420 20802 63924 20804
rect 63420 20750 63422 20802
rect 63474 20750 63870 20802
rect 63922 20750 63924 20802
rect 63420 20748 63924 20750
rect 63420 20738 63476 20748
rect 62412 20132 62468 20142
rect 61852 19406 61854 19458
rect 61906 19406 61908 19458
rect 61852 19394 61908 19406
rect 61964 20018 62020 20030
rect 61964 19966 61966 20018
rect 62018 19966 62020 20018
rect 61516 19236 61572 19246
rect 61516 19142 61572 19180
rect 61852 19236 61908 19246
rect 61964 19236 62020 19966
rect 62412 19906 62468 20076
rect 63084 20132 63140 20142
rect 63196 20132 63476 20188
rect 63084 20038 63140 20076
rect 62412 19854 62414 19906
rect 62466 19854 62468 19906
rect 62412 19842 62468 19854
rect 61852 19234 62020 19236
rect 61852 19182 61854 19234
rect 61906 19182 62020 19234
rect 61852 19180 62020 19182
rect 63196 19236 63252 19246
rect 61292 18452 61348 18462
rect 61292 18358 61348 18396
rect 60396 15184 60452 15260
rect 60620 15932 60900 15988
rect 61180 18340 61236 18350
rect 60508 14530 60564 14542
rect 60508 14478 60510 14530
rect 60562 14478 60564 14530
rect 60508 14420 60564 14478
rect 60508 14354 60564 14364
rect 60284 14308 60340 14318
rect 60284 13746 60340 14252
rect 60284 13694 60286 13746
rect 60338 13694 60340 13746
rect 60284 13682 60340 13694
rect 59388 12786 59444 12796
rect 59836 13132 60228 13188
rect 59172 12572 59436 12582
rect 59228 12516 59276 12572
rect 59332 12516 59380 12572
rect 59172 12506 59436 12516
rect 59500 12178 59556 12190
rect 59500 12126 59502 12178
rect 59554 12126 59556 12178
rect 58940 11284 58996 11294
rect 58940 11190 58996 11228
rect 59500 11284 59556 12126
rect 59500 11218 59556 11228
rect 59724 12066 59780 12078
rect 59724 12014 59726 12066
rect 59778 12014 59780 12066
rect 59724 11956 59780 12014
rect 59172 11004 59436 11014
rect 59228 10948 59276 11004
rect 59332 10948 59380 11004
rect 59172 10938 59436 10948
rect 59052 9602 59108 9614
rect 59052 9550 59054 9602
rect 59106 9550 59108 9602
rect 59052 8428 59108 9550
rect 59500 9604 59556 9614
rect 59500 9602 59668 9604
rect 59500 9550 59502 9602
rect 59554 9550 59668 9602
rect 59500 9548 59668 9550
rect 59500 9538 59556 9548
rect 59172 9436 59436 9446
rect 59228 9380 59276 9436
rect 59332 9380 59380 9436
rect 59172 9370 59436 9380
rect 59612 8428 59668 9548
rect 59724 8818 59780 11900
rect 59724 8766 59726 8818
rect 59778 8766 59780 8818
rect 59724 8754 59780 8766
rect 58940 8372 59108 8428
rect 59500 8372 59668 8428
rect 58828 8260 58884 8270
rect 58828 8034 58884 8204
rect 58828 7982 58830 8034
rect 58882 7982 58884 8034
rect 58828 7588 58884 7982
rect 58828 7522 58884 7532
rect 58716 7310 58718 7362
rect 58770 7310 58772 7362
rect 58716 7250 58772 7310
rect 58716 7198 58718 7250
rect 58770 7198 58772 7250
rect 58716 7186 58772 7198
rect 58940 7140 58996 8372
rect 59052 8148 59108 8158
rect 59052 7700 59108 8092
rect 59172 7868 59436 7878
rect 59228 7812 59276 7868
rect 59332 7812 59380 7868
rect 59172 7802 59436 7812
rect 59164 7700 59220 7710
rect 59052 7698 59220 7700
rect 59052 7646 59166 7698
rect 59218 7646 59220 7698
rect 59052 7644 59220 7646
rect 59164 7634 59220 7644
rect 59500 7364 59556 8372
rect 59612 8260 59668 8270
rect 59612 8166 59668 8204
rect 59388 7308 59556 7364
rect 59724 7362 59780 7374
rect 59724 7310 59726 7362
rect 59778 7310 59780 7362
rect 59388 7252 59444 7308
rect 59724 7252 59780 7310
rect 59388 7186 59444 7196
rect 59500 7196 59780 7252
rect 58940 7074 58996 7084
rect 59052 6804 59108 6814
rect 58268 5058 58324 5068
rect 58380 6466 58436 6478
rect 58380 6414 58382 6466
rect 58434 6414 58436 6466
rect 58380 6020 58436 6414
rect 58940 6132 58996 6142
rect 58940 6038 58996 6076
rect 59052 6130 59108 6748
rect 59164 6580 59220 6590
rect 59164 6486 59220 6524
rect 59172 6300 59436 6310
rect 59228 6244 59276 6300
rect 59332 6244 59380 6300
rect 59172 6234 59436 6244
rect 59052 6078 59054 6130
rect 59106 6078 59108 6130
rect 59052 6066 59108 6078
rect 58044 4900 58100 4910
rect 57932 4898 58100 4900
rect 57932 4846 58046 4898
rect 58098 4846 58100 4898
rect 57932 4844 58100 4846
rect 57932 4562 57988 4844
rect 58044 4834 58100 4844
rect 58380 4788 58436 5964
rect 58828 5908 58884 5918
rect 58828 5814 58884 5852
rect 59164 5906 59220 5918
rect 59164 5854 59166 5906
rect 59218 5854 59220 5906
rect 58492 5796 58548 5806
rect 58492 5702 58548 5740
rect 59052 5348 59108 5358
rect 58828 5346 59108 5348
rect 58828 5294 59054 5346
rect 59106 5294 59108 5346
rect 58828 5292 59108 5294
rect 58828 5124 58884 5292
rect 59052 5282 59108 5292
rect 58380 4722 58436 4732
rect 58604 5068 58884 5124
rect 58604 5010 58660 5068
rect 58604 4958 58606 5010
rect 58658 4958 58660 5010
rect 57932 4510 57934 4562
rect 57986 4510 57988 4562
rect 57932 4228 57988 4510
rect 58604 4564 58660 4958
rect 58044 4340 58100 4350
rect 58044 4246 58100 4284
rect 58156 4338 58212 4350
rect 58156 4286 58158 4338
rect 58210 4286 58212 4338
rect 57932 4162 57988 4172
rect 57820 3938 57876 3948
rect 58156 4004 58212 4286
rect 58380 4340 58436 4350
rect 58604 4340 58660 4508
rect 58380 4338 58660 4340
rect 58380 4286 58382 4338
rect 58434 4286 58660 4338
rect 58380 4284 58660 4286
rect 58716 4900 58772 4910
rect 58716 4452 58772 4844
rect 58828 4452 58884 5068
rect 59164 5124 59220 5854
rect 59276 5346 59332 5358
rect 59276 5294 59278 5346
rect 59330 5294 59332 5346
rect 59276 5234 59332 5294
rect 59276 5182 59278 5234
rect 59330 5182 59332 5234
rect 59276 5170 59332 5182
rect 59164 5058 59220 5068
rect 58940 4900 58996 4910
rect 58940 4806 58996 4844
rect 59172 4732 59436 4742
rect 59228 4676 59276 4732
rect 59332 4676 59380 4732
rect 59172 4666 59436 4676
rect 58940 4452 58996 4462
rect 58828 4450 58996 4452
rect 58828 4398 58942 4450
rect 58994 4398 58996 4450
rect 58828 4396 58996 4398
rect 58380 4274 58436 4284
rect 58156 3938 58212 3948
rect 57484 3502 57486 3554
rect 57538 3502 57540 3554
rect 57484 2660 57540 3502
rect 58044 3442 58100 3454
rect 58044 3390 58046 3442
rect 58098 3390 58100 3442
rect 58044 3332 58100 3390
rect 58044 3266 58100 3276
rect 58156 3444 58212 3454
rect 57484 2594 57540 2604
rect 58156 2212 58212 3388
rect 58604 3444 58660 3454
rect 58716 3444 58772 4396
rect 58940 4386 58996 4396
rect 59052 4452 59108 4462
rect 59052 4450 59220 4452
rect 59052 4398 59054 4450
rect 59106 4398 59220 4450
rect 59052 4396 59220 4398
rect 59052 4386 59108 4396
rect 59052 4114 59108 4126
rect 59052 4062 59054 4114
rect 59106 4062 59108 4114
rect 58604 3442 58772 3444
rect 58604 3390 58606 3442
rect 58658 3390 58772 3442
rect 58604 3388 58772 3390
rect 58940 3444 58996 3454
rect 58604 3378 58660 3388
rect 58940 3350 58996 3388
rect 59052 2996 59108 4062
rect 59164 4004 59220 4396
rect 59500 4228 59556 7196
rect 59724 6692 59780 6702
rect 59836 6692 59892 13132
rect 60620 13076 60676 15932
rect 60732 15314 60788 15326
rect 60732 15262 60734 15314
rect 60786 15262 60788 15314
rect 60732 13972 60788 15262
rect 60732 13916 61012 13972
rect 60956 13634 61012 13916
rect 61068 13860 61124 13870
rect 61068 13766 61124 13804
rect 60956 13582 60958 13634
rect 61010 13582 61012 13634
rect 60956 13570 61012 13582
rect 60620 13010 60676 13020
rect 59948 12962 60004 12974
rect 59948 12910 59950 12962
rect 60002 12910 60004 12962
rect 59948 12852 60004 12910
rect 59948 12786 60004 12796
rect 60172 12964 60228 12974
rect 60172 12290 60228 12908
rect 60172 12238 60174 12290
rect 60226 12238 60228 12290
rect 60172 12226 60228 12238
rect 60732 12066 60788 12078
rect 60732 12014 60734 12066
rect 60786 12014 60788 12066
rect 60508 11284 60564 11294
rect 60732 11284 60788 12014
rect 60956 11956 61012 11966
rect 60956 11862 61012 11900
rect 60564 11228 60788 11284
rect 60508 11190 60564 11228
rect 59948 9716 60004 9726
rect 60004 9660 60116 9716
rect 59948 9622 60004 9660
rect 60060 8428 60116 9660
rect 60172 9492 60228 9502
rect 60172 9042 60228 9436
rect 60172 8990 60174 9042
rect 60226 8990 60228 9042
rect 60172 8978 60228 8990
rect 60844 9042 60900 9054
rect 60844 8990 60846 9042
rect 60898 8990 60900 9042
rect 60844 8932 60900 8990
rect 60844 8866 60900 8876
rect 61180 8428 61236 18284
rect 61740 18338 61796 18350
rect 61740 18286 61742 18338
rect 61794 18286 61796 18338
rect 61740 17556 61796 18286
rect 61852 17778 61908 19180
rect 63196 19142 63252 19180
rect 62748 19012 62804 19022
rect 61852 17726 61854 17778
rect 61906 17726 61908 17778
rect 61852 17714 61908 17726
rect 62076 18450 62132 18462
rect 62076 18398 62078 18450
rect 62130 18398 62132 18450
rect 62076 17668 62132 18398
rect 62076 17536 62132 17612
rect 61740 17462 61796 17500
rect 61292 17220 61348 17230
rect 61292 16882 61348 17164
rect 61292 16830 61294 16882
rect 61346 16830 61348 16882
rect 61292 16100 61348 16830
rect 61404 17108 61460 17118
rect 61404 16994 61460 17052
rect 61404 16942 61406 16994
rect 61458 16942 61460 16994
rect 61404 16884 61460 16942
rect 61852 16996 61908 17006
rect 61404 16818 61460 16828
rect 61628 16882 61684 16894
rect 61628 16830 61630 16882
rect 61682 16830 61684 16882
rect 61628 16436 61684 16830
rect 61628 16370 61684 16380
rect 61740 16884 61796 16894
rect 61404 16100 61460 16110
rect 61292 16098 61460 16100
rect 61292 16046 61406 16098
rect 61458 16046 61460 16098
rect 61292 16044 61460 16046
rect 61740 16100 61796 16828
rect 61852 16882 61908 16940
rect 61852 16830 61854 16882
rect 61906 16830 61908 16882
rect 61852 16818 61908 16830
rect 62636 16770 62692 16782
rect 62636 16718 62638 16770
rect 62690 16718 62692 16770
rect 62300 16658 62356 16670
rect 62300 16606 62302 16658
rect 62354 16606 62356 16658
rect 62076 16436 62132 16446
rect 61964 16212 62020 16222
rect 61964 16118 62020 16156
rect 61852 16100 61908 16110
rect 61740 16098 61908 16100
rect 61740 16046 61854 16098
rect 61906 16046 61908 16098
rect 61740 16044 61908 16046
rect 61292 15538 61348 16044
rect 61404 16034 61460 16044
rect 61852 16034 61908 16044
rect 62076 16100 62132 16380
rect 62300 16324 62356 16606
rect 62636 16436 62692 16718
rect 62636 16370 62692 16380
rect 62300 16258 62356 16268
rect 62636 16212 62692 16222
rect 62636 16118 62692 16156
rect 62076 16098 62356 16100
rect 62076 16046 62078 16098
rect 62130 16046 62356 16098
rect 62076 16044 62356 16046
rect 62076 16034 62132 16044
rect 61628 15876 61684 15886
rect 61628 15782 61684 15820
rect 62076 15876 62132 15886
rect 61292 15486 61294 15538
rect 61346 15486 61348 15538
rect 61292 15474 61348 15486
rect 61964 15540 62020 15550
rect 62076 15540 62132 15820
rect 61964 15538 62132 15540
rect 61964 15486 61966 15538
rect 62018 15486 62132 15538
rect 61964 15484 62132 15486
rect 62300 15652 62356 16044
rect 62748 15652 62804 18956
rect 63420 18228 63476 20132
rect 63868 20132 63924 20748
rect 63868 20066 63924 20076
rect 63644 20020 63700 20030
rect 63644 19346 63700 19964
rect 63980 19796 64036 21308
rect 64092 20188 64148 23102
rect 64652 23154 64708 25566
rect 65212 25620 65268 26124
rect 65212 25554 65268 25564
rect 65884 25732 65940 26908
rect 68460 26852 68516 26862
rect 68460 26758 68516 26796
rect 68684 26850 68740 26862
rect 68684 26798 68686 26850
rect 68738 26798 68740 26850
rect 67004 26402 67060 26414
rect 67004 26350 67006 26402
rect 67058 26350 67060 26402
rect 65996 26180 66052 26190
rect 65996 26086 66052 26124
rect 66780 26066 66836 26078
rect 66780 26014 66782 26066
rect 66834 26014 66836 26066
rect 65884 25676 66164 25732
rect 65436 25396 65492 25406
rect 64764 24948 64820 24958
rect 65436 24948 65492 25340
rect 65548 24948 65604 24958
rect 65436 24946 65604 24948
rect 65436 24894 65550 24946
rect 65602 24894 65604 24946
rect 65436 24892 65604 24894
rect 64764 24854 64820 24892
rect 64988 24724 65044 24734
rect 64764 24162 64820 24174
rect 64764 24110 64766 24162
rect 64818 24110 64820 24162
rect 64764 24050 64820 24110
rect 64764 23998 64766 24050
rect 64818 23998 64820 24050
rect 64764 23986 64820 23998
rect 64988 23604 65044 24668
rect 65436 24724 65492 24734
rect 65436 24630 65492 24668
rect 65100 24162 65156 24174
rect 65100 24110 65102 24162
rect 65154 24110 65156 24162
rect 65100 23940 65156 24110
rect 65548 24052 65604 24892
rect 65772 24948 65828 24958
rect 65884 24948 65940 25676
rect 66108 25620 66164 25676
rect 66780 25730 66836 26014
rect 66780 25678 66782 25730
rect 66834 25678 66836 25730
rect 66780 25620 66836 25678
rect 66108 25618 66612 25620
rect 66108 25566 66110 25618
rect 66162 25566 66612 25618
rect 66108 25564 66612 25566
rect 66108 25554 66164 25564
rect 65772 24946 65940 24948
rect 65772 24894 65774 24946
rect 65826 24894 65940 24946
rect 65772 24892 65940 24894
rect 65996 25506 66052 25518
rect 65996 25454 65998 25506
rect 66050 25454 66052 25506
rect 65996 24948 66052 25454
rect 65772 24882 65828 24892
rect 65996 24882 66052 24892
rect 66332 25396 66388 25406
rect 65324 23940 65380 23950
rect 65100 23938 65380 23940
rect 65100 23886 65326 23938
rect 65378 23886 65380 23938
rect 65100 23884 65380 23886
rect 65324 23874 65380 23884
rect 65436 23828 65492 23838
rect 65548 23828 65604 23996
rect 65436 23826 65604 23828
rect 65436 23774 65438 23826
rect 65490 23774 65604 23826
rect 65436 23772 65604 23774
rect 65436 23762 65492 23772
rect 64988 23538 65044 23548
rect 65324 23604 65380 23614
rect 64652 23102 64654 23154
rect 64706 23102 64708 23154
rect 64204 22484 64260 22494
rect 64652 22484 64708 23102
rect 64204 22482 64708 22484
rect 64204 22430 64206 22482
rect 64258 22430 64708 22482
rect 64204 22428 64708 22430
rect 64204 22418 64260 22428
rect 64652 22372 64708 22428
rect 64876 23492 64932 23502
rect 64764 22372 64820 22382
rect 64652 22370 64820 22372
rect 64652 22318 64766 22370
rect 64818 22318 64820 22370
rect 64652 22316 64820 22318
rect 64764 22306 64820 22316
rect 64876 22260 64932 23436
rect 65324 23378 65380 23548
rect 65548 23492 65604 23772
rect 66332 23938 66388 25340
rect 66556 24834 66612 25564
rect 66780 25554 66836 25564
rect 67004 25396 67060 26350
rect 67900 26402 67956 26414
rect 67900 26350 67902 26402
rect 67954 26350 67956 26402
rect 67116 26068 67172 26078
rect 67116 25974 67172 26012
rect 67676 26068 67732 26078
rect 67676 25974 67732 26012
rect 67788 25620 67844 25630
rect 67788 25526 67844 25564
rect 66668 25284 66724 25294
rect 66668 24946 66724 25228
rect 66668 24894 66670 24946
rect 66722 24894 66724 24946
rect 66668 24882 66724 24894
rect 66780 24948 66836 24958
rect 66556 24782 66558 24834
rect 66610 24782 66612 24834
rect 66556 24770 66612 24782
rect 66780 24612 66836 24892
rect 66780 24546 66836 24556
rect 66332 23886 66334 23938
rect 66386 23886 66388 23938
rect 66332 23828 66388 23886
rect 66668 23940 66724 23950
rect 67004 23940 67060 25340
rect 67676 25506 67732 25518
rect 67676 25454 67678 25506
rect 67730 25454 67732 25506
rect 67676 25396 67732 25454
rect 67676 25330 67732 25340
rect 67900 25284 67956 26350
rect 68012 26292 68068 26302
rect 68684 26292 68740 26798
rect 69580 26516 69636 27694
rect 71148 27524 71204 27534
rect 69804 27076 69860 27086
rect 69692 26516 69748 26526
rect 69580 26514 69748 26516
rect 69580 26462 69694 26514
rect 69746 26462 69748 26514
rect 69580 26460 69748 26462
rect 69692 26450 69748 26460
rect 69804 26514 69860 27020
rect 69804 26462 69806 26514
rect 69858 26462 69860 26514
rect 69804 26450 69860 26462
rect 69916 27074 69972 27086
rect 69916 27022 69918 27074
rect 69970 27022 69972 27074
rect 69916 26852 69972 27022
rect 70476 27076 70532 27086
rect 69132 26292 69188 26302
rect 68684 26290 69188 26292
rect 68684 26238 69134 26290
rect 69186 26238 69188 26290
rect 68684 26236 69188 26238
rect 68012 26178 68068 26236
rect 69132 26226 69188 26236
rect 69580 26292 69636 26302
rect 69580 26198 69636 26236
rect 68012 26126 68014 26178
rect 68066 26126 68068 26178
rect 68012 26114 68068 26126
rect 68832 25900 69096 25910
rect 67900 25218 67956 25228
rect 68124 25844 68180 25854
rect 68888 25844 68936 25900
rect 68992 25844 69040 25900
rect 68832 25834 69096 25844
rect 67788 24724 67844 24734
rect 67788 24630 67844 24668
rect 67228 24612 67284 24622
rect 66668 23938 67060 23940
rect 66668 23886 66670 23938
rect 66722 23886 67060 23938
rect 66668 23884 67060 23886
rect 67116 24052 67172 24062
rect 66668 23874 66724 23884
rect 66332 23762 66388 23772
rect 65660 23716 65716 23726
rect 66444 23716 66500 23726
rect 65660 23714 66164 23716
rect 65660 23662 65662 23714
rect 65714 23662 66164 23714
rect 65660 23660 66164 23662
rect 65660 23650 65716 23660
rect 65548 23436 65716 23492
rect 65324 23326 65326 23378
rect 65378 23326 65380 23378
rect 65324 23314 65380 23326
rect 65100 22372 65156 22382
rect 65100 22278 65156 22316
rect 64876 22128 64932 22204
rect 65324 22260 65380 22270
rect 64540 21812 64596 21822
rect 64316 21588 64372 21598
rect 64316 21494 64372 21532
rect 64540 20914 64596 21756
rect 64540 20862 64542 20914
rect 64594 20862 64596 20914
rect 64540 20850 64596 20862
rect 64652 21700 64708 21710
rect 64652 20188 64708 21644
rect 64092 20132 64484 20188
rect 63980 19730 64036 19740
rect 64204 20020 64260 20030
rect 64204 19460 64260 19964
rect 64316 19460 64372 19470
rect 64204 19458 64372 19460
rect 64204 19406 64318 19458
rect 64370 19406 64372 19458
rect 64204 19404 64372 19406
rect 63644 19294 63646 19346
rect 63698 19294 63700 19346
rect 63644 19282 63700 19294
rect 63980 19348 64036 19358
rect 63980 18452 64036 19292
rect 64092 19236 64148 19246
rect 64316 19236 64372 19404
rect 64148 19180 64260 19236
rect 64092 19104 64148 19180
rect 64204 19124 64260 19180
rect 64316 19170 64372 19180
rect 64092 18452 64148 18462
rect 63980 18450 64148 18452
rect 63980 18398 64094 18450
rect 64146 18398 64148 18450
rect 63980 18396 64148 18398
rect 64092 18386 64148 18396
rect 63196 17780 63252 17790
rect 63084 17444 63140 17454
rect 62972 17442 63140 17444
rect 62972 17390 63086 17442
rect 63138 17390 63140 17442
rect 62972 17388 63140 17390
rect 62860 16212 62916 16222
rect 62860 16118 62916 16156
rect 62972 15988 63028 17388
rect 63084 17378 63140 17388
rect 63084 17108 63140 17118
rect 63196 17108 63252 17724
rect 63140 17052 63252 17108
rect 63420 17778 63476 18172
rect 63868 17892 63924 17902
rect 63420 17726 63422 17778
rect 63474 17726 63476 17778
rect 63084 17014 63140 17052
rect 63420 16884 63476 17726
rect 63420 16818 63476 16828
rect 63756 17890 63924 17892
rect 63756 17838 63870 17890
rect 63922 17838 63924 17890
rect 63756 17836 63924 17838
rect 63644 16212 63700 16222
rect 63644 16118 63700 16156
rect 62972 15922 63028 15932
rect 63196 15874 63252 15886
rect 63196 15822 63198 15874
rect 63250 15822 63252 15874
rect 62748 15596 63140 15652
rect 62300 15538 62356 15596
rect 62300 15486 62302 15538
rect 62354 15486 62356 15538
rect 61964 15474 62020 15484
rect 62300 15474 62356 15486
rect 62972 15428 63028 15438
rect 61516 15316 61572 15326
rect 61516 14642 61572 15260
rect 62972 15314 63028 15372
rect 62972 15262 62974 15314
rect 63026 15262 63028 15314
rect 62972 15250 63028 15262
rect 62860 15204 62916 15214
rect 61516 14590 61518 14642
rect 61570 14590 61572 14642
rect 61516 14578 61572 14590
rect 62748 15202 62916 15204
rect 62748 15150 62862 15202
rect 62914 15150 62916 15202
rect 62748 15148 62916 15150
rect 62076 14532 62132 14542
rect 62412 14532 62468 14542
rect 62076 14530 62468 14532
rect 62076 14478 62078 14530
rect 62130 14478 62414 14530
rect 62466 14478 62468 14530
rect 62076 14476 62468 14478
rect 62076 14466 62132 14476
rect 62412 14466 62468 14476
rect 61292 14420 61348 14430
rect 61292 13522 61348 14364
rect 62748 14418 62804 15148
rect 62860 15138 62916 15148
rect 62748 14366 62750 14418
rect 62802 14366 62804 14418
rect 61404 14308 61460 14318
rect 61404 14214 61460 14252
rect 61628 14306 61684 14318
rect 61628 14254 61630 14306
rect 61682 14254 61684 14306
rect 61292 13470 61294 13522
rect 61346 13470 61348 13522
rect 61292 13458 61348 13470
rect 61516 13860 61572 13870
rect 61516 13074 61572 13804
rect 61628 13524 61684 14254
rect 62524 14308 62580 14318
rect 62524 13858 62580 14252
rect 62524 13806 62526 13858
rect 62578 13806 62580 13858
rect 62524 13794 62580 13806
rect 62636 14306 62692 14318
rect 62636 14254 62638 14306
rect 62690 14254 62692 14306
rect 61628 13458 61684 13468
rect 61964 13634 62020 13646
rect 61964 13582 61966 13634
rect 62018 13582 62020 13634
rect 61516 13022 61518 13074
rect 61570 13022 61572 13074
rect 61516 13010 61572 13022
rect 61292 12964 61348 12974
rect 61292 12870 61348 12908
rect 61852 12962 61908 12974
rect 61852 12910 61854 12962
rect 61906 12910 61908 12962
rect 61740 12852 61796 12862
rect 61740 12758 61796 12796
rect 61292 12404 61348 12414
rect 61852 12404 61908 12910
rect 61964 12740 62020 13582
rect 62636 13524 62692 14254
rect 62748 13746 62804 14366
rect 62748 13694 62750 13746
rect 62802 13694 62804 13746
rect 62748 13682 62804 13694
rect 62972 13746 63028 13758
rect 62972 13694 62974 13746
rect 63026 13694 63028 13746
rect 62972 13524 63028 13694
rect 62636 13468 63028 13524
rect 61964 12674 62020 12684
rect 62412 12740 62468 12750
rect 62412 12646 62468 12684
rect 62860 12738 62916 12750
rect 62860 12686 62862 12738
rect 62914 12686 62916 12738
rect 61292 12402 61908 12404
rect 61292 12350 61294 12402
rect 61346 12350 61908 12402
rect 61292 12348 61908 12350
rect 62412 12516 62468 12526
rect 61292 12338 61348 12348
rect 61964 12290 62020 12302
rect 61964 12238 61966 12290
rect 62018 12238 62020 12290
rect 61964 12180 62020 12238
rect 62076 12292 62132 12302
rect 62076 12198 62132 12236
rect 61964 12114 62020 12124
rect 61964 11956 62020 11966
rect 61964 11954 62132 11956
rect 61964 11902 61966 11954
rect 62018 11902 62132 11954
rect 61964 11900 62132 11902
rect 61964 11890 62020 11900
rect 61516 11282 61572 11294
rect 61516 11230 61518 11282
rect 61570 11230 61572 11282
rect 61516 10612 61572 11230
rect 61516 9042 61572 10556
rect 61964 10722 62020 10734
rect 61964 10670 61966 10722
rect 62018 10670 62020 10722
rect 61628 10052 61684 10062
rect 61964 10052 62020 10670
rect 61684 9996 61908 10052
rect 61628 9986 61684 9996
rect 61852 9940 61908 9996
rect 61964 9986 62020 9996
rect 61852 9874 61908 9884
rect 61516 8990 61518 9042
rect 61570 8990 61572 9042
rect 61516 8978 61572 8990
rect 62076 9044 62132 11900
rect 62300 11508 62356 11518
rect 62300 11414 62356 11452
rect 62188 11394 62244 11406
rect 62188 11342 62190 11394
rect 62242 11342 62244 11394
rect 62188 10836 62244 11342
rect 62188 10770 62244 10780
rect 62300 10836 62356 10846
rect 62412 10836 62468 12460
rect 62524 12292 62580 12302
rect 62524 12198 62580 12236
rect 62860 12180 62916 12686
rect 62972 12740 63028 13468
rect 62972 12674 63028 12684
rect 63084 12628 63140 15596
rect 63196 15316 63252 15822
rect 63308 15316 63364 15326
rect 63196 15314 63588 15316
rect 63196 15262 63310 15314
rect 63362 15262 63588 15314
rect 63196 15260 63588 15262
rect 63308 15250 63364 15260
rect 63084 12562 63140 12572
rect 63308 15092 63364 15102
rect 63196 12180 63252 12190
rect 62860 12114 62916 12124
rect 63084 12178 63252 12180
rect 63084 12126 63198 12178
rect 63250 12126 63252 12178
rect 63084 12124 63252 12126
rect 62300 10834 62468 10836
rect 62300 10782 62302 10834
rect 62354 10782 62468 10834
rect 62300 10780 62468 10782
rect 63084 10834 63140 12124
rect 63196 12114 63252 12124
rect 63308 12068 63364 15036
rect 63532 14644 63588 15260
rect 63644 14644 63700 14654
rect 63532 14642 63700 14644
rect 63532 14590 63646 14642
rect 63698 14590 63700 14642
rect 63532 14588 63700 14590
rect 63644 14578 63700 14588
rect 63420 12292 63476 12302
rect 63420 12198 63476 12236
rect 63532 12180 63588 12190
rect 63532 12178 63700 12180
rect 63532 12126 63534 12178
rect 63586 12126 63700 12178
rect 63532 12124 63700 12126
rect 63532 12114 63588 12124
rect 63308 12012 63476 12068
rect 63308 11508 63364 11518
rect 63308 10948 63364 11452
rect 63308 10882 63364 10892
rect 63084 10782 63086 10834
rect 63138 10782 63140 10834
rect 62300 10770 62356 10780
rect 63084 10770 63140 10782
rect 63196 10836 63252 10846
rect 62188 10612 62244 10622
rect 62188 10518 62244 10556
rect 62412 10610 62468 10622
rect 62412 10558 62414 10610
rect 62466 10558 62468 10610
rect 62412 10050 62468 10558
rect 63196 10612 63252 10780
rect 63308 10612 63364 10622
rect 63196 10610 63364 10612
rect 63196 10558 63310 10610
rect 63362 10558 63364 10610
rect 63196 10556 63364 10558
rect 63308 10546 63364 10556
rect 63420 10610 63476 12012
rect 63532 11844 63588 11854
rect 63532 11396 63588 11788
rect 63644 11508 63700 12124
rect 63756 11956 63812 17836
rect 63868 17826 63924 17836
rect 64204 17890 64260 19068
rect 64428 19012 64484 20132
rect 64204 17838 64206 17890
rect 64258 17838 64260 17890
rect 64204 17826 64260 17838
rect 64316 18956 64484 19012
rect 64540 20132 64708 20188
rect 65212 20916 65268 20926
rect 65212 20802 65268 20860
rect 65212 20750 65214 20802
rect 65266 20750 65268 20802
rect 63868 17442 63924 17454
rect 63868 17390 63870 17442
rect 63922 17390 63924 17442
rect 63868 17220 63924 17390
rect 64316 17220 64372 18956
rect 63868 16996 63924 17164
rect 63868 16930 63924 16940
rect 63980 17164 64372 17220
rect 64428 17442 64484 17454
rect 64428 17390 64430 17442
rect 64482 17390 64484 17442
rect 63980 15652 64036 17164
rect 64428 17108 64484 17390
rect 64428 17042 64484 17052
rect 63980 15586 64036 15596
rect 64092 16996 64148 17006
rect 64092 16882 64148 16940
rect 64092 16830 64094 16882
rect 64146 16830 64148 16882
rect 63868 15428 63924 15438
rect 63868 14754 63924 15372
rect 64092 15204 64148 16830
rect 64204 16884 64260 16894
rect 64428 16884 64484 16894
rect 64204 16882 64372 16884
rect 64204 16830 64206 16882
rect 64258 16830 64372 16882
rect 64204 16828 64372 16830
rect 64204 16818 64260 16828
rect 64092 15138 64148 15148
rect 64204 16100 64260 16110
rect 63868 14702 63870 14754
rect 63922 14702 63924 14754
rect 63868 14690 63924 14702
rect 63980 14756 64036 14766
rect 63980 12964 64036 14700
rect 64204 14754 64260 16044
rect 64316 16098 64372 16828
rect 64428 16790 64484 16828
rect 64316 16046 64318 16098
rect 64370 16046 64372 16098
rect 64316 15988 64372 16046
rect 64316 15538 64372 15932
rect 64316 15486 64318 15538
rect 64370 15486 64372 15538
rect 64316 15474 64372 15486
rect 64540 14980 64596 20132
rect 64764 19908 64820 19918
rect 64764 19814 64820 19852
rect 64652 19012 64708 19022
rect 64652 19010 64820 19012
rect 64652 18958 64654 19010
rect 64706 18958 64820 19010
rect 64652 18956 64820 18958
rect 64652 18946 64708 18956
rect 64652 18450 64708 18462
rect 64652 18398 64654 18450
rect 64706 18398 64708 18450
rect 64652 17444 64708 18398
rect 64764 18452 64820 18956
rect 64764 18386 64820 18396
rect 64876 17890 64932 17902
rect 64876 17838 64878 17890
rect 64930 17838 64932 17890
rect 64876 17778 64932 17838
rect 64876 17726 64878 17778
rect 64930 17726 64932 17778
rect 64876 17714 64932 17726
rect 65212 17444 65268 20750
rect 65324 20692 65380 22204
rect 65548 22260 65604 22270
rect 65548 22166 65604 22204
rect 65660 22258 65716 23436
rect 66108 23156 66164 23660
rect 66444 23622 66500 23660
rect 67004 23716 67060 23726
rect 67116 23716 67172 23996
rect 67004 23714 67172 23716
rect 67004 23662 67006 23714
rect 67058 23662 67172 23714
rect 67004 23660 67172 23662
rect 67004 23650 67060 23660
rect 65884 23044 65940 23054
rect 65660 22206 65662 22258
rect 65714 22206 65716 22258
rect 65660 22148 65716 22206
rect 65660 22082 65716 22092
rect 65772 23042 65940 23044
rect 65772 22990 65886 23042
rect 65938 22990 65940 23042
rect 65772 22988 65940 22990
rect 65772 21924 65828 22988
rect 65884 22978 65940 22988
rect 65996 23044 66052 23054
rect 66108 23024 66164 23100
rect 67116 23042 67172 23054
rect 65772 21810 65828 21868
rect 65772 21758 65774 21810
rect 65826 21758 65828 21810
rect 65772 21746 65828 21758
rect 65884 22146 65940 22158
rect 65884 22094 65886 22146
rect 65938 22094 65940 22146
rect 65548 21700 65604 21710
rect 65548 21606 65604 21644
rect 65324 20560 65380 20636
rect 65436 21588 65492 21598
rect 65324 20244 65380 20254
rect 65436 20244 65492 21532
rect 65660 21588 65716 21598
rect 65548 20804 65604 20814
rect 65548 20710 65604 20748
rect 65324 20242 65492 20244
rect 65324 20190 65326 20242
rect 65378 20190 65492 20242
rect 65324 20188 65492 20190
rect 65660 20188 65716 21532
rect 65884 21588 65940 22094
rect 65884 21522 65940 21532
rect 65324 20178 65380 20188
rect 65548 20132 65716 20188
rect 65772 20692 65828 20702
rect 65436 19234 65492 19246
rect 65436 19182 65438 19234
rect 65490 19182 65492 19234
rect 65436 19124 65492 19182
rect 65436 19058 65492 19068
rect 65548 18674 65604 20132
rect 65772 19906 65828 20636
rect 65996 20188 66052 22988
rect 67116 22990 67118 23042
rect 67170 22990 67172 23042
rect 66444 22932 66500 22942
rect 66444 22930 66948 22932
rect 66444 22878 66446 22930
rect 66498 22878 66948 22930
rect 66444 22876 66948 22878
rect 66444 22866 66500 22876
rect 66892 22482 66948 22876
rect 66892 22430 66894 22482
rect 66946 22430 66948 22482
rect 66892 22418 66948 22430
rect 66668 22372 66724 22382
rect 66668 22278 66724 22316
rect 67116 22372 67172 22990
rect 67228 22372 67284 24556
rect 67340 24610 67396 24622
rect 67340 24558 67342 24610
rect 67394 24558 67396 24610
rect 67340 24052 67396 24558
rect 67340 23986 67396 23996
rect 67900 23828 67956 23838
rect 67452 23716 67508 23726
rect 67452 23622 67508 23660
rect 67900 23716 67956 23772
rect 67900 23714 68068 23716
rect 67900 23662 67902 23714
rect 67954 23662 68068 23714
rect 67900 23660 68068 23662
rect 67900 23650 67956 23660
rect 67452 23266 67508 23278
rect 67452 23214 67454 23266
rect 67506 23214 67508 23266
rect 67340 22372 67396 22382
rect 67228 22370 67396 22372
rect 67228 22318 67342 22370
rect 67394 22318 67396 22370
rect 67228 22316 67396 22318
rect 67116 22306 67172 22316
rect 67340 22306 67396 22316
rect 66108 22260 66164 22270
rect 66108 21812 66164 22204
rect 66108 21746 66164 21756
rect 66444 22148 66500 22158
rect 66332 21476 66388 21486
rect 66108 20914 66164 20926
rect 66108 20862 66110 20914
rect 66162 20862 66164 20914
rect 66108 20804 66164 20862
rect 66108 20738 66164 20748
rect 65772 19854 65774 19906
rect 65826 19854 65828 19906
rect 65548 18622 65550 18674
rect 65602 18622 65604 18674
rect 65548 17890 65604 18622
rect 65660 19794 65716 19806
rect 65660 19742 65662 19794
rect 65714 19742 65716 19794
rect 65660 18562 65716 19742
rect 65772 18788 65828 19854
rect 65884 20132 66052 20188
rect 66332 20690 66388 21420
rect 66332 20638 66334 20690
rect 66386 20638 66388 20690
rect 65884 19794 65940 20132
rect 65884 19742 65886 19794
rect 65938 19742 65940 19794
rect 65884 19730 65940 19742
rect 66332 19908 66388 20638
rect 66444 20188 66500 22092
rect 67116 22146 67172 22158
rect 67116 22094 67118 22146
rect 67170 22094 67172 22146
rect 66556 21588 66612 21598
rect 66556 21494 66612 21532
rect 67116 21588 67172 22094
rect 67228 22146 67284 22158
rect 67228 22094 67230 22146
rect 67282 22094 67284 22146
rect 67228 22036 67284 22094
rect 67228 21970 67284 21980
rect 67452 21924 67508 23214
rect 67900 22148 67956 22158
rect 67900 22054 67956 22092
rect 67116 21522 67172 21532
rect 67340 21868 67452 21924
rect 66892 21362 66948 21374
rect 66892 21310 66894 21362
rect 66946 21310 66948 21362
rect 66668 20804 66724 20814
rect 66444 20132 66612 20188
rect 66108 19234 66164 19246
rect 66108 19182 66110 19234
rect 66162 19182 66164 19234
rect 65772 18732 65940 18788
rect 65884 18676 65940 18732
rect 66108 18676 66164 19182
rect 65884 18620 66052 18676
rect 65660 18510 65662 18562
rect 65714 18510 65716 18562
rect 65660 18498 65716 18510
rect 65772 18450 65828 18462
rect 65772 18398 65774 18450
rect 65826 18398 65828 18450
rect 65772 18340 65828 18398
rect 65884 18452 65940 18462
rect 65884 18358 65940 18396
rect 65772 18274 65828 18284
rect 65548 17838 65550 17890
rect 65602 17838 65604 17890
rect 65548 17826 65604 17838
rect 65772 17890 65828 17902
rect 65772 17838 65774 17890
rect 65826 17838 65828 17890
rect 65772 17778 65828 17838
rect 65772 17726 65774 17778
rect 65826 17726 65828 17778
rect 65772 17714 65828 17726
rect 65996 17556 66052 18620
rect 65660 17500 66052 17556
rect 66108 18228 66164 18620
rect 66220 18228 66276 18238
rect 66108 18226 66276 18228
rect 66108 18174 66222 18226
rect 66274 18174 66276 18226
rect 66108 18172 66276 18174
rect 65324 17444 65380 17454
rect 65212 17388 65324 17444
rect 65380 17388 65492 17444
rect 64652 17378 64708 17388
rect 65324 17350 65380 17388
rect 64652 17220 64708 17230
rect 64652 16994 64708 17164
rect 64652 16942 64654 16994
rect 64706 16942 64708 16994
rect 64652 16548 64708 16942
rect 64764 16884 64820 16894
rect 64764 16770 64820 16828
rect 64764 16718 64766 16770
rect 64818 16718 64820 16770
rect 64764 16706 64820 16718
rect 64652 16492 64932 16548
rect 64876 16100 64932 16492
rect 64988 16324 65044 16334
rect 64988 16230 65044 16268
rect 65324 16100 65380 16110
rect 64876 16098 65380 16100
rect 64876 16046 65326 16098
rect 65378 16046 65380 16098
rect 64876 16044 65380 16046
rect 64876 15986 64932 16044
rect 65324 16034 65380 16044
rect 64876 15934 64878 15986
rect 64930 15934 64932 15986
rect 64876 15922 64932 15934
rect 64652 15876 64708 15886
rect 64652 15782 64708 15820
rect 65324 15204 65380 15214
rect 65324 15110 65380 15148
rect 64652 14980 64708 14990
rect 64540 14924 64652 14980
rect 64204 14702 64206 14754
rect 64258 14702 64260 14754
rect 64204 14690 64260 14702
rect 64652 13970 64708 14924
rect 65436 14084 65492 17388
rect 65548 16770 65604 16782
rect 65548 16718 65550 16770
rect 65602 16718 65604 16770
rect 65548 16324 65604 16718
rect 65548 16258 65604 16268
rect 64652 13918 64654 13970
rect 64706 13918 64708 13970
rect 64652 13860 64708 13918
rect 64652 13794 64708 13804
rect 65324 14028 65492 14084
rect 64988 13748 65044 13758
rect 64428 13076 64484 13086
rect 64428 12982 64484 13020
rect 63980 12962 64372 12964
rect 63980 12910 63982 12962
rect 64034 12910 64372 12962
rect 63980 12908 64372 12910
rect 63980 12898 64036 12908
rect 64316 12516 64372 12908
rect 64988 12962 65044 13692
rect 64988 12910 64990 12962
rect 65042 12910 65044 12962
rect 64988 12898 65044 12910
rect 65324 13076 65380 14028
rect 65436 13860 65492 13870
rect 65436 13766 65492 13804
rect 65548 13858 65604 13870
rect 65548 13806 65550 13858
rect 65602 13806 65604 13858
rect 65548 13412 65604 13806
rect 65548 13188 65604 13356
rect 65548 13122 65604 13132
rect 65436 13076 65492 13086
rect 65324 13074 65492 13076
rect 65324 13022 65438 13074
rect 65490 13022 65492 13074
rect 65324 13020 65492 13022
rect 65324 12740 65380 13020
rect 65436 13010 65492 13020
rect 65660 12852 65716 17500
rect 65772 16996 65828 17006
rect 65772 16882 65828 16940
rect 65772 16830 65774 16882
rect 65826 16830 65828 16882
rect 65772 16818 65828 16830
rect 65884 15876 65940 15886
rect 66108 15876 66164 18172
rect 66220 18162 66276 18172
rect 66220 16100 66276 16110
rect 66220 16006 66276 16044
rect 66108 15820 66276 15876
rect 65884 15538 65940 15820
rect 65884 15486 65886 15538
rect 65938 15486 65940 15538
rect 65884 15474 65940 15486
rect 65324 12674 65380 12684
rect 65436 12796 65716 12852
rect 65772 15428 65828 15438
rect 65772 13746 65828 15372
rect 66108 14420 66164 14430
rect 66108 14326 66164 14364
rect 65772 13694 65774 13746
rect 65826 13694 65828 13746
rect 64316 12460 64708 12516
rect 63756 11890 63812 11900
rect 63868 12292 63924 12302
rect 63868 12068 63924 12236
rect 63980 12068 64036 12078
rect 63868 12066 64036 12068
rect 63868 12014 63982 12066
rect 64034 12014 64036 12066
rect 63868 12012 64036 12014
rect 63756 11508 63812 11518
rect 63644 11452 63756 11508
rect 63756 11414 63812 11452
rect 63532 11340 63700 11396
rect 63532 10948 63588 10958
rect 63532 10834 63588 10892
rect 63532 10782 63534 10834
rect 63586 10782 63588 10834
rect 63532 10770 63588 10782
rect 63420 10558 63422 10610
rect 63474 10558 63476 10610
rect 63420 10546 63476 10558
rect 62412 9998 62414 10050
rect 62466 9998 62468 10050
rect 62412 9986 62468 9998
rect 63420 10052 63476 10062
rect 63420 9958 63476 9996
rect 62412 9826 62468 9838
rect 62412 9774 62414 9826
rect 62466 9774 62468 9826
rect 62412 9716 62468 9774
rect 62300 9044 62356 9054
rect 62076 9042 62356 9044
rect 62076 8990 62302 9042
rect 62354 8990 62356 9042
rect 62076 8988 62356 8990
rect 59780 6636 59892 6692
rect 59948 8372 60116 8428
rect 60396 8372 60452 8382
rect 59948 6692 60004 8372
rect 60396 8278 60452 8316
rect 60844 8372 61236 8428
rect 61628 8372 61684 8382
rect 60284 8260 60340 8270
rect 60284 8166 60340 8204
rect 60732 7700 60788 7710
rect 59724 6598 59780 6636
rect 59948 6626 60004 6636
rect 60060 7362 60116 7374
rect 60060 7310 60062 7362
rect 60114 7310 60116 7362
rect 60060 7252 60116 7310
rect 60060 6356 60116 7196
rect 60508 7362 60564 7374
rect 60508 7310 60510 7362
rect 60562 7310 60564 7362
rect 60508 7250 60564 7310
rect 60508 7198 60510 7250
rect 60562 7198 60564 7250
rect 60284 7140 60340 7150
rect 60172 6468 60228 6478
rect 60172 6374 60228 6412
rect 60060 6290 60116 6300
rect 60060 5906 60116 5918
rect 60060 5854 60062 5906
rect 60114 5854 60116 5906
rect 59948 5796 60004 5806
rect 59948 5702 60004 5740
rect 60060 5348 60116 5854
rect 60060 5282 60116 5292
rect 60172 5348 60228 5358
rect 60284 5348 60340 7084
rect 60508 6580 60564 7198
rect 60620 7364 60676 7374
rect 60620 6802 60676 7308
rect 60620 6750 60622 6802
rect 60674 6750 60676 6802
rect 60620 6738 60676 6750
rect 60508 6514 60564 6524
rect 60732 6020 60788 7644
rect 60172 5346 60340 5348
rect 60172 5294 60174 5346
rect 60226 5294 60340 5346
rect 60172 5292 60340 5294
rect 60508 5964 60788 6020
rect 60172 5282 60228 5292
rect 60508 5236 60564 5964
rect 59612 5124 59668 5134
rect 59612 4562 59668 5068
rect 60396 5012 60452 5022
rect 60396 4918 60452 4956
rect 60508 5010 60564 5180
rect 60508 4958 60510 5010
rect 60562 4958 60564 5010
rect 60508 4946 60564 4958
rect 60732 5124 60788 5134
rect 60844 5124 60900 8372
rect 61628 8278 61684 8316
rect 61068 8260 61124 8270
rect 61068 7698 61124 8204
rect 62076 8258 62132 8988
rect 62300 8978 62356 8988
rect 62412 8932 62468 9660
rect 62748 9714 62804 9726
rect 62748 9662 62750 9714
rect 62802 9662 62804 9714
rect 62748 9492 62804 9662
rect 63420 9716 63476 9726
rect 63420 9622 63476 9660
rect 63532 9714 63588 9726
rect 63532 9662 63534 9714
rect 63586 9662 63588 9714
rect 62748 9426 62804 9436
rect 63084 9492 63140 9502
rect 62860 9380 62916 9390
rect 62748 9268 62804 9278
rect 62748 9174 62804 9212
rect 62860 9266 62916 9324
rect 62860 9214 62862 9266
rect 62914 9214 62916 9266
rect 62860 9202 62916 9214
rect 62972 9042 63028 9054
rect 62972 8990 62974 9042
rect 63026 8990 63028 9042
rect 62412 8866 62468 8876
rect 62524 8930 62580 8942
rect 62524 8878 62526 8930
rect 62578 8878 62580 8930
rect 62524 8428 62580 8878
rect 62412 8372 62580 8428
rect 62972 8372 63028 8990
rect 62412 8306 62468 8316
rect 62972 8306 63028 8316
rect 63084 8370 63140 9436
rect 63532 9492 63588 9662
rect 63532 9426 63588 9436
rect 63532 9268 63588 9278
rect 63532 9174 63588 9212
rect 63084 8318 63086 8370
rect 63138 8318 63140 8370
rect 63084 8306 63140 8318
rect 62076 8206 62078 8258
rect 62130 8206 62132 8258
rect 62076 8194 62132 8206
rect 63308 8258 63364 8270
rect 63308 8206 63310 8258
rect 63362 8206 63364 8258
rect 62524 8148 62580 8158
rect 63308 8148 63364 8206
rect 62524 8146 63364 8148
rect 62524 8094 62526 8146
rect 62578 8094 63364 8146
rect 62524 8092 63364 8094
rect 62524 8082 62580 8092
rect 61068 7646 61070 7698
rect 61122 7646 61124 7698
rect 61068 7634 61124 7646
rect 61292 7812 61348 7822
rect 61292 7476 61348 7756
rect 63084 7700 63140 7710
rect 60732 5122 60900 5124
rect 60732 5070 60734 5122
rect 60786 5070 60900 5122
rect 60732 5068 60900 5070
rect 61068 6692 61124 6702
rect 61068 5796 61124 6636
rect 61292 6690 61348 7420
rect 62636 7474 62692 7486
rect 62636 7422 62638 7474
rect 62690 7422 62692 7474
rect 61404 7362 61460 7374
rect 61404 7310 61406 7362
rect 61458 7310 61460 7362
rect 61404 7140 61460 7310
rect 61404 7074 61460 7084
rect 61852 7362 61908 7374
rect 61852 7310 61854 7362
rect 61906 7310 61908 7362
rect 61852 7250 61908 7310
rect 61852 7198 61854 7250
rect 61906 7198 61908 7250
rect 61292 6638 61294 6690
rect 61346 6638 61348 6690
rect 61292 6626 61348 6638
rect 61852 6244 61908 7198
rect 62076 7028 62132 7038
rect 62076 6690 62132 6972
rect 62076 6638 62078 6690
rect 62130 6638 62132 6690
rect 62076 6626 62132 6638
rect 62188 6802 62244 6814
rect 62188 6750 62190 6802
rect 62242 6750 62244 6802
rect 61852 6178 61908 6188
rect 62188 6020 62244 6750
rect 62636 6130 62692 7422
rect 62636 6078 62638 6130
rect 62690 6078 62692 6130
rect 62636 6066 62692 6078
rect 62860 7028 62916 7038
rect 62860 6130 62916 6972
rect 62972 6692 63028 6702
rect 63084 6692 63140 7644
rect 63308 7586 63364 8092
rect 63532 8258 63588 8270
rect 63532 8206 63534 8258
rect 63586 8206 63588 8258
rect 63532 7700 63588 8206
rect 63532 7634 63588 7644
rect 63308 7534 63310 7586
rect 63362 7534 63364 7586
rect 63308 7522 63364 7534
rect 63196 7364 63252 7374
rect 63196 7270 63252 7308
rect 62972 6690 63140 6692
rect 62972 6638 62974 6690
rect 63026 6638 63140 6690
rect 62972 6636 63140 6638
rect 62972 6626 63028 6636
rect 63420 6466 63476 6478
rect 63420 6414 63422 6466
rect 63474 6414 63476 6466
rect 63420 6356 63476 6414
rect 63420 6290 63476 6300
rect 63644 6244 63700 11340
rect 63868 11394 63924 12012
rect 63980 12002 64036 12012
rect 63868 11342 63870 11394
rect 63922 11342 63924 11394
rect 63868 11172 63924 11342
rect 63868 11106 63924 11116
rect 64540 10052 64596 12460
rect 64652 12402 64708 12460
rect 64652 12350 64654 12402
rect 64706 12350 64708 12402
rect 64652 12338 64708 12350
rect 65436 12180 65492 12796
rect 64764 11172 64820 11182
rect 64764 11078 64820 11116
rect 65436 10612 65492 12124
rect 65548 12068 65604 12078
rect 65548 11974 65604 12012
rect 65548 10612 65604 10622
rect 65436 10610 65604 10612
rect 65436 10558 65550 10610
rect 65602 10558 65604 10610
rect 65436 10556 65604 10558
rect 65548 10546 65604 10556
rect 64652 10498 64708 10510
rect 64652 10446 64654 10498
rect 64706 10446 64708 10498
rect 64652 10276 64708 10446
rect 64652 10210 64708 10220
rect 64540 9986 64596 9996
rect 65548 9940 65604 9950
rect 65548 9846 65604 9884
rect 65100 9602 65156 9614
rect 65772 9604 65828 13694
rect 66108 13636 66164 13646
rect 66108 13542 66164 13580
rect 66220 13412 66276 15820
rect 66332 15428 66388 19852
rect 66444 16996 66500 17006
rect 66444 16770 66500 16940
rect 66444 16718 66446 16770
rect 66498 16718 66500 16770
rect 66444 16210 66500 16718
rect 66444 16158 66446 16210
rect 66498 16158 66500 16210
rect 66444 16146 66500 16158
rect 66556 15988 66612 20132
rect 66668 20018 66724 20748
rect 66668 19966 66670 20018
rect 66722 19966 66724 20018
rect 66668 19954 66724 19966
rect 66892 20018 66948 21310
rect 67228 20468 67284 20478
rect 67228 20130 67284 20412
rect 67340 20242 67396 21868
rect 67452 21858 67508 21868
rect 67564 21588 67620 21598
rect 67452 21476 67508 21486
rect 67452 21382 67508 21420
rect 67564 20802 67620 21532
rect 67788 21474 67844 21486
rect 67788 21422 67790 21474
rect 67842 21422 67844 21474
rect 67788 20916 67844 21422
rect 67788 20850 67844 20860
rect 68012 20916 68068 23660
rect 68012 20850 68068 20860
rect 67564 20750 67566 20802
rect 67618 20750 67620 20802
rect 67564 20738 67620 20750
rect 67340 20190 67342 20242
rect 67394 20190 67396 20242
rect 67340 20178 67396 20190
rect 68124 20188 68180 25788
rect 69804 25620 69860 25630
rect 69916 25620 69972 26796
rect 70364 26962 70420 26974
rect 70364 26910 70366 26962
rect 70418 26910 70420 26962
rect 70364 26402 70420 26910
rect 70476 26514 70532 27020
rect 71036 27076 71092 27086
rect 71036 26982 71092 27020
rect 70476 26462 70478 26514
rect 70530 26462 70532 26514
rect 70476 26450 70532 26462
rect 70364 26350 70366 26402
rect 70418 26350 70420 26402
rect 70364 26338 70420 26350
rect 69804 25618 69972 25620
rect 69804 25566 69806 25618
rect 69858 25566 69972 25618
rect 69804 25564 69972 25566
rect 69804 25554 69860 25564
rect 69244 25506 69300 25518
rect 69244 25454 69246 25506
rect 69298 25454 69300 25506
rect 68572 25396 68628 25406
rect 68572 25302 68628 25340
rect 69020 24836 69076 24846
rect 69020 24742 69076 24780
rect 68832 24332 69096 24342
rect 68888 24276 68936 24332
rect 68992 24276 69040 24332
rect 68832 24266 69096 24276
rect 69244 23940 69300 25454
rect 69916 25396 69972 25406
rect 69916 25302 69972 25340
rect 70588 25396 70644 25406
rect 69692 25284 69748 25294
rect 69692 25282 69860 25284
rect 69692 25230 69694 25282
rect 69746 25230 69860 25282
rect 69692 25228 69860 25230
rect 69692 25218 69748 25228
rect 69804 24836 69860 25228
rect 69804 24742 69860 24780
rect 70588 24610 70644 25340
rect 70700 24836 70756 24846
rect 70700 24722 70756 24780
rect 70700 24670 70702 24722
rect 70754 24670 70756 24722
rect 70700 24658 70756 24670
rect 70588 24558 70590 24610
rect 70642 24558 70644 24610
rect 70588 24546 70644 24558
rect 71148 24500 71204 27468
rect 71372 27300 71428 27916
rect 71596 27972 71652 29484
rect 71932 28642 71988 30156
rect 72044 30146 72100 30156
rect 72156 30212 72212 31612
rect 72268 31444 72324 31454
rect 72268 31218 72324 31388
rect 72268 31166 72270 31218
rect 72322 31166 72324 31218
rect 72268 30322 72324 31166
rect 72268 30270 72270 30322
rect 72322 30270 72324 30322
rect 72268 30258 72324 30270
rect 72156 30146 72212 30156
rect 71932 28590 71934 28642
rect 71986 28590 71988 28642
rect 71932 28578 71988 28590
rect 72044 29314 72100 29326
rect 72044 29262 72046 29314
rect 72098 29262 72100 29314
rect 72044 27972 72100 29262
rect 72380 29204 72436 33068
rect 73388 32564 73444 32574
rect 73388 32002 73444 32508
rect 73388 31950 73390 32002
rect 73442 31950 73444 32002
rect 73388 31938 73444 31950
rect 73500 31666 73556 31678
rect 73500 31614 73502 31666
rect 73554 31614 73556 31666
rect 73388 31554 73444 31566
rect 73388 31502 73390 31554
rect 73442 31502 73444 31554
rect 73388 31220 73444 31502
rect 73500 31332 73556 31614
rect 73500 31266 73556 31276
rect 73388 31154 73444 31164
rect 72380 29138 72436 29148
rect 72716 30100 72772 30110
rect 72716 29986 72772 30044
rect 72716 29934 72718 29986
rect 72770 29934 72772 29986
rect 72716 28644 72772 29934
rect 72716 28578 72772 28588
rect 71596 27970 72100 27972
rect 71596 27918 71598 27970
rect 71650 27918 72100 27970
rect 71596 27916 72100 27918
rect 71596 27906 71652 27916
rect 71372 27234 71428 27244
rect 72044 27746 72100 27916
rect 72044 27694 72046 27746
rect 72098 27694 72100 27746
rect 71260 27074 71316 27086
rect 71260 27022 71262 27074
rect 71314 27022 71316 27074
rect 71260 26292 71316 27022
rect 71260 26226 71316 26236
rect 71932 27076 71988 27086
rect 71932 26290 71988 27020
rect 71932 26238 71934 26290
rect 71986 26238 71988 26290
rect 71932 26226 71988 26238
rect 72044 26068 72100 27694
rect 73052 27300 73108 27310
rect 73052 27206 73108 27244
rect 72492 27076 72548 27086
rect 72716 27076 72772 27086
rect 72492 26982 72548 27020
rect 72604 27074 72772 27076
rect 72604 27022 72718 27074
rect 72770 27022 72772 27074
rect 72604 27020 72772 27022
rect 72044 26002 72100 26012
rect 72268 26964 72324 26974
rect 72268 26066 72324 26908
rect 72268 26014 72270 26066
rect 72322 26014 72324 26066
rect 72268 26002 72324 26014
rect 72380 26292 72436 26302
rect 72604 26292 72660 27020
rect 72716 27010 72772 27020
rect 72380 26290 72660 26292
rect 72380 26238 72382 26290
rect 72434 26238 72660 26290
rect 72380 26236 72660 26238
rect 72380 25730 72436 26236
rect 72380 25678 72382 25730
rect 72434 25678 72436 25730
rect 72380 25666 72436 25678
rect 72492 25396 72548 25406
rect 72492 25394 73332 25396
rect 72492 25342 72494 25394
rect 72546 25342 73332 25394
rect 72492 25340 73332 25342
rect 72492 25330 72548 25340
rect 72380 25284 72436 25294
rect 72268 25282 72436 25284
rect 72268 25230 72382 25282
rect 72434 25230 72436 25282
rect 72268 25228 72436 25230
rect 72268 24946 72324 25228
rect 72380 25218 72436 25228
rect 72268 24894 72270 24946
rect 72322 24894 72324 24946
rect 72268 24882 72324 24894
rect 73276 24946 73332 25340
rect 73276 24894 73278 24946
rect 73330 24894 73332 24946
rect 73276 24882 73332 24894
rect 72044 24836 72100 24846
rect 72044 24834 72212 24836
rect 72044 24782 72046 24834
rect 72098 24782 72212 24834
rect 72044 24780 72212 24782
rect 72044 24770 72100 24780
rect 71372 24722 71428 24734
rect 71932 24724 71988 24734
rect 71372 24670 71374 24722
rect 71426 24670 71428 24722
rect 71372 24612 71428 24670
rect 71820 24722 71988 24724
rect 71820 24670 71934 24722
rect 71986 24670 71988 24722
rect 71820 24668 71988 24670
rect 71820 24612 71876 24668
rect 71932 24658 71988 24668
rect 71372 24556 71876 24612
rect 71148 24444 71652 24500
rect 69244 23874 69300 23884
rect 68572 23156 68628 23166
rect 68572 23062 68628 23100
rect 71260 23154 71316 23166
rect 71260 23102 71262 23154
rect 71314 23102 71316 23154
rect 69244 23042 69300 23054
rect 69244 22990 69246 23042
rect 69298 22990 69300 23042
rect 68832 22764 69096 22774
rect 68888 22708 68936 22764
rect 68992 22708 69040 22764
rect 68832 22698 69096 22708
rect 69244 22484 69300 22990
rect 69244 22418 69300 22428
rect 70588 23044 70644 23054
rect 70588 22482 70644 22988
rect 71260 23044 71316 23102
rect 70588 22430 70590 22482
rect 70642 22430 70644 22482
rect 70588 22418 70644 22430
rect 71148 22596 71204 22606
rect 71148 22370 71204 22540
rect 71148 22318 71150 22370
rect 71202 22318 71204 22370
rect 71148 22306 71204 22318
rect 68348 22260 68404 22270
rect 68348 22166 68404 22204
rect 71260 22258 71316 22988
rect 71372 23042 71428 23054
rect 71372 22990 71374 23042
rect 71426 22990 71428 23042
rect 71372 22708 71428 22990
rect 71372 22642 71428 22652
rect 71484 22596 71540 22606
rect 71484 22370 71540 22540
rect 71484 22318 71486 22370
rect 71538 22318 71540 22370
rect 71484 22306 71540 22318
rect 71260 22206 71262 22258
rect 71314 22206 71316 22258
rect 71260 22194 71316 22206
rect 71036 22148 71092 22158
rect 71596 22148 71652 24444
rect 71820 24050 71876 24556
rect 71820 23998 71822 24050
rect 71874 23998 71876 24050
rect 71820 23986 71876 23998
rect 72156 23938 72212 24780
rect 72156 23886 72158 23938
rect 72210 23886 72212 23938
rect 72156 23380 72212 23886
rect 73500 24834 73556 24846
rect 73500 24782 73502 24834
rect 73554 24782 73556 24834
rect 73500 24612 73556 24782
rect 72604 23826 72660 23838
rect 72604 23774 72606 23826
rect 72658 23774 72660 23826
rect 72604 23492 72660 23774
rect 73500 23604 73556 24556
rect 72604 23426 72660 23436
rect 73276 23548 73556 23604
rect 73612 24722 73668 24734
rect 73612 24670 73614 24722
rect 73666 24670 73668 24722
rect 72156 23314 72212 23324
rect 72156 23156 72212 23166
rect 72156 22372 72212 23100
rect 73276 23044 73332 23548
rect 73612 23492 73668 24670
rect 73612 23426 73668 23436
rect 73500 23380 73556 23390
rect 73500 23286 73556 23324
rect 72492 22484 72548 22494
rect 72492 22390 72548 22428
rect 72268 22372 72324 22382
rect 72156 22370 72324 22372
rect 72156 22318 72270 22370
rect 72322 22318 72324 22370
rect 72156 22316 72324 22318
rect 72268 22306 72324 22316
rect 72940 22372 72996 22382
rect 72940 22278 72996 22316
rect 69468 21474 69524 21486
rect 69468 21422 69470 21474
rect 69522 21422 69524 21474
rect 68832 21196 69096 21206
rect 68888 21140 68936 21196
rect 68992 21140 69040 21196
rect 68832 21130 69096 21140
rect 69244 20916 69300 20926
rect 68236 20692 68292 20702
rect 68236 20598 68292 20636
rect 68124 20132 68292 20188
rect 67228 20078 67230 20130
rect 67282 20078 67284 20130
rect 67228 20066 67284 20078
rect 67116 20020 67172 20030
rect 66892 19966 66894 20018
rect 66946 19966 66948 20018
rect 66892 19954 66948 19966
rect 67004 20018 67172 20020
rect 67004 19966 67118 20018
rect 67170 19966 67172 20018
rect 67004 19964 67172 19966
rect 67004 19908 67060 19964
rect 67116 19954 67172 19964
rect 66780 19236 66836 19246
rect 66780 19142 66836 19180
rect 67004 19012 67060 19852
rect 67900 19908 67956 19918
rect 67900 19814 67956 19852
rect 67564 19124 67620 19134
rect 67564 19030 67620 19068
rect 66780 18956 67060 19012
rect 68012 19010 68068 19022
rect 68012 18958 68014 19010
rect 68066 18958 68068 19010
rect 66668 18340 66724 18350
rect 66668 18246 66724 18284
rect 66332 15362 66388 15372
rect 66444 15932 66612 15988
rect 65100 9550 65102 9602
rect 65154 9550 65156 9602
rect 64092 9044 64148 9054
rect 64092 8428 64148 8988
rect 64540 8930 64596 8942
rect 64540 8878 64542 8930
rect 64594 8878 64596 8930
rect 63756 8372 63812 8382
rect 64092 8372 64260 8428
rect 63756 6692 63812 8316
rect 63868 7362 63924 7374
rect 63868 7310 63870 7362
rect 63922 7310 63924 7362
rect 63868 6916 63924 7310
rect 63868 6850 63924 6860
rect 63980 7250 64036 7262
rect 63980 7198 63982 7250
rect 64034 7198 64036 7250
rect 63756 6626 63812 6636
rect 63868 6468 63924 6478
rect 63980 6468 64036 7198
rect 63868 6466 64036 6468
rect 63868 6414 63870 6466
rect 63922 6414 64036 6466
rect 63868 6412 64036 6414
rect 62860 6078 62862 6130
rect 62914 6078 62916 6130
rect 62860 6066 62916 6078
rect 63532 6188 63700 6244
rect 63756 6244 63812 6254
rect 59612 4510 59614 4562
rect 59666 4510 59668 4562
rect 59612 4498 59668 4510
rect 59724 4898 59780 4910
rect 59724 4846 59726 4898
rect 59778 4846 59780 4898
rect 59500 4162 59556 4172
rect 59164 3938 59220 3948
rect 59724 3892 59780 4846
rect 59948 4564 60004 4574
rect 59836 4452 59892 4462
rect 59836 4358 59892 4396
rect 59948 4450 60004 4508
rect 59948 4398 59950 4450
rect 60002 4398 60004 4450
rect 59724 3826 59780 3836
rect 59612 3780 59668 3790
rect 59612 3686 59668 3724
rect 59500 3556 59556 3566
rect 59500 3462 59556 3500
rect 59948 3556 60004 4398
rect 60396 4452 60452 4462
rect 60396 4228 60452 4396
rect 60396 4162 60452 4172
rect 60732 3892 60788 5068
rect 61068 4564 61124 5740
rect 61516 5906 61572 5918
rect 61516 5854 61518 5906
rect 61570 5854 61572 5906
rect 62188 5888 62244 5964
rect 62972 6020 63028 6030
rect 62972 5926 63028 5964
rect 62524 5908 62580 5918
rect 61292 4900 61348 4910
rect 61068 4498 61124 4508
rect 61180 4898 61348 4900
rect 61180 4846 61294 4898
rect 61346 4846 61348 4898
rect 61180 4844 61348 4846
rect 60732 3826 60788 3836
rect 59948 3490 60004 3500
rect 60172 3556 60228 3566
rect 59612 3332 59668 3342
rect 59612 3238 59668 3276
rect 59172 3164 59436 3174
rect 59228 3108 59276 3164
rect 59332 3108 59380 3164
rect 59172 3098 59436 3108
rect 59052 2930 59108 2940
rect 56924 914 56980 924
rect 58044 2156 58212 2212
rect 58044 800 58100 2156
rect 60172 800 60228 3500
rect 60508 3332 60564 3342
rect 60508 3238 60564 3276
rect 61180 2884 61236 4844
rect 61292 4834 61348 4844
rect 61516 4900 61572 5854
rect 62076 5684 62132 5694
rect 61292 4676 61348 4686
rect 61292 4338 61348 4620
rect 61516 4562 61572 4844
rect 61964 5236 62020 5246
rect 61964 4900 62020 5180
rect 61964 4834 62020 4844
rect 61516 4510 61518 4562
rect 61570 4510 61572 4562
rect 61516 4498 61572 4510
rect 61292 4286 61294 4338
rect 61346 4286 61348 4338
rect 61292 3780 61348 4286
rect 61628 4340 61684 4350
rect 61628 4246 61684 4284
rect 61964 4340 62020 4350
rect 62076 4340 62132 5628
rect 62524 5122 62580 5852
rect 62524 5070 62526 5122
rect 62578 5070 62580 5122
rect 61964 4338 62132 4340
rect 61964 4286 61966 4338
rect 62018 4286 62132 4338
rect 61964 4284 62132 4286
rect 62300 4452 62356 4462
rect 61964 4274 62020 4284
rect 61292 3714 61348 3724
rect 61404 4226 61460 4238
rect 61404 4174 61406 4226
rect 61458 4174 61460 4226
rect 61404 3332 61460 4174
rect 61404 3266 61460 3276
rect 61180 2818 61236 2828
rect 62300 800 62356 4396
rect 62524 4226 62580 5070
rect 63420 5124 63476 5134
rect 63532 5124 63588 6188
rect 63644 6018 63700 6030
rect 63644 5966 63646 6018
rect 63698 5966 63700 6018
rect 63644 5908 63700 5966
rect 63756 6018 63812 6188
rect 63756 5966 63758 6018
rect 63810 5966 63812 6018
rect 63756 5954 63812 5966
rect 63644 5842 63700 5852
rect 63644 5684 63700 5694
rect 63644 5590 63700 5628
rect 63868 5124 63924 6412
rect 64204 6020 64260 8372
rect 64316 7362 64372 7374
rect 64316 7310 64318 7362
rect 64370 7310 64372 7362
rect 64316 7028 64372 7310
rect 64316 6972 64484 7028
rect 64428 6578 64484 6972
rect 64540 6692 64596 8878
rect 65100 8820 65156 9550
rect 65660 9548 65828 9604
rect 65884 13356 66276 13412
rect 66332 14644 66388 14654
rect 65436 9044 65492 9054
rect 65436 8950 65492 8988
rect 65100 8754 65156 8764
rect 65212 8932 65268 8942
rect 64988 8260 65044 8270
rect 64988 8166 65044 8204
rect 64652 8034 64708 8046
rect 64652 7982 64654 8034
rect 64706 7982 64708 8034
rect 64652 7588 64708 7982
rect 65212 8034 65268 8876
rect 65212 7982 65214 8034
rect 65266 7982 65268 8034
rect 64652 7532 65044 7588
rect 64988 7476 65044 7532
rect 64652 7362 64708 7374
rect 64652 7310 64654 7362
rect 64706 7310 64708 7362
rect 64652 7250 64708 7310
rect 64652 7198 64654 7250
rect 64706 7198 64708 7250
rect 64652 7186 64708 7198
rect 64876 7140 64932 7150
rect 64764 6692 64820 6702
rect 64540 6636 64708 6692
rect 64428 6526 64430 6578
rect 64482 6526 64484 6578
rect 63420 5122 63588 5124
rect 63420 5070 63422 5122
rect 63474 5070 63588 5122
rect 63420 5068 63588 5070
rect 63756 5068 63924 5124
rect 64092 5964 64260 6020
rect 64316 6244 64372 6254
rect 63084 5010 63140 5022
rect 63084 4958 63086 5010
rect 63138 4958 63140 5010
rect 63084 4564 63140 4958
rect 63196 4900 63252 4910
rect 63196 4806 63252 4844
rect 63084 4498 63140 4508
rect 62524 4174 62526 4226
rect 62578 4174 62580 4226
rect 62524 4162 62580 4174
rect 63420 4228 63476 5068
rect 63756 4900 63812 5068
rect 63756 4834 63812 4844
rect 63868 4898 63924 4910
rect 63868 4846 63870 4898
rect 63922 4846 63924 4898
rect 63868 4788 63924 4846
rect 63532 4452 63588 4462
rect 63532 4358 63588 4396
rect 63420 4162 63476 4172
rect 63868 4116 63924 4732
rect 64092 4788 64148 5964
rect 64092 4722 64148 4732
rect 64204 5794 64260 5806
rect 64204 5742 64206 5794
rect 64258 5742 64260 5794
rect 64204 5012 64260 5742
rect 64316 5234 64372 6188
rect 64316 5182 64318 5234
rect 64370 5182 64372 5234
rect 64316 5170 64372 5182
rect 64428 6020 64484 6526
rect 64428 5012 64484 5964
rect 63868 4050 63924 4060
rect 63532 3668 63588 3678
rect 63532 3574 63588 3612
rect 64204 3668 64260 4956
rect 64204 3602 64260 3612
rect 64316 4956 64484 5012
rect 64540 6468 64596 6478
rect 62972 3556 63028 3566
rect 62972 3442 63028 3500
rect 62972 3390 62974 3442
rect 63026 3390 63028 3442
rect 62972 3378 63028 3390
rect 64316 2772 64372 4956
rect 64540 4900 64596 6412
rect 64652 6020 64708 6636
rect 64764 6598 64820 6636
rect 64652 5964 64820 6020
rect 64652 5796 64708 5806
rect 64652 5702 64708 5740
rect 64540 4834 64596 4844
rect 64428 4564 64484 4574
rect 64428 4470 64484 4508
rect 64764 3556 64820 5964
rect 64876 5234 64932 7084
rect 64988 6244 65044 7420
rect 65212 6468 65268 7982
rect 65324 8820 65380 8830
rect 65324 8484 65380 8764
rect 65324 8146 65380 8428
rect 65324 8094 65326 8146
rect 65378 8094 65380 8146
rect 65324 7028 65380 8094
rect 65548 7924 65604 7934
rect 65548 7698 65604 7868
rect 65548 7646 65550 7698
rect 65602 7646 65604 7698
rect 65548 7634 65604 7646
rect 65436 7476 65492 7486
rect 65436 7382 65492 7420
rect 65660 7140 65716 9548
rect 65772 8932 65828 8942
rect 65772 8838 65828 8876
rect 65772 8484 65828 8494
rect 65772 8370 65828 8428
rect 65772 8318 65774 8370
rect 65826 8318 65828 8370
rect 65772 8306 65828 8318
rect 65772 7700 65828 7710
rect 65884 7700 65940 13356
rect 66332 13074 66388 14588
rect 66332 13022 66334 13074
rect 66386 13022 66388 13074
rect 66332 13010 66388 13022
rect 66220 12740 66276 12750
rect 65996 12628 66052 12638
rect 65996 12402 66052 12572
rect 65996 12350 65998 12402
rect 66050 12350 66052 12402
rect 65996 12338 66052 12350
rect 66220 11506 66276 12684
rect 66220 11454 66222 11506
rect 66274 11454 66276 11506
rect 66220 11442 66276 11454
rect 65996 10610 66052 10622
rect 65996 10558 65998 10610
rect 66050 10558 66052 10610
rect 65996 10276 66052 10558
rect 65996 10210 66052 10220
rect 66444 9940 66500 15932
rect 66780 14308 66836 18956
rect 67228 18676 67284 18686
rect 67116 18452 67172 18462
rect 67228 18452 67284 18620
rect 68012 18676 68068 18958
rect 68012 18610 68068 18620
rect 67116 18450 67284 18452
rect 67116 18398 67118 18450
rect 67170 18398 67284 18450
rect 67116 18396 67284 18398
rect 68124 18564 68180 18574
rect 67116 18386 67172 18396
rect 67228 17780 67284 17790
rect 66892 16884 66948 16894
rect 66892 16790 66948 16828
rect 66892 15986 66948 15998
rect 66892 15934 66894 15986
rect 66946 15934 66948 15986
rect 66892 14532 66948 15934
rect 67004 14644 67060 14654
rect 67004 14550 67060 14588
rect 66892 14400 66948 14476
rect 66780 14252 66948 14308
rect 66556 13748 66612 13758
rect 66556 13654 66612 13692
rect 66780 12964 66836 12974
rect 66668 12740 66724 12750
rect 66556 12628 66612 12638
rect 66556 11506 66612 12572
rect 66668 12290 66724 12684
rect 66780 12516 66836 12908
rect 66780 12450 66836 12460
rect 66668 12238 66670 12290
rect 66722 12238 66724 12290
rect 66668 12226 66724 12238
rect 66780 12292 66836 12302
rect 66780 11956 66836 12236
rect 66780 11890 66836 11900
rect 66556 11454 66558 11506
rect 66610 11454 66612 11506
rect 66556 11172 66612 11454
rect 66556 11106 66612 11116
rect 66668 11508 66724 11518
rect 66668 10722 66724 11452
rect 66668 10670 66670 10722
rect 66722 10670 66724 10722
rect 66668 10658 66724 10670
rect 66444 9874 66500 9884
rect 66668 10052 66724 10062
rect 66108 9602 66164 9614
rect 66108 9550 66110 9602
rect 66162 9550 66164 9602
rect 66108 8932 66164 9550
rect 66332 8932 66388 8942
rect 66108 8930 66388 8932
rect 66108 8878 66334 8930
rect 66386 8878 66388 8930
rect 66108 8876 66388 8878
rect 66332 8596 66388 8876
rect 66332 8530 66388 8540
rect 66668 8484 66724 9996
rect 66780 9156 66836 9166
rect 66780 9062 66836 9100
rect 66668 8258 66724 8428
rect 66668 8206 66670 8258
rect 66722 8206 66724 8258
rect 66668 8194 66724 8206
rect 66780 8596 66836 8606
rect 66780 8146 66836 8540
rect 66892 8428 66948 14252
rect 67116 14196 67172 14206
rect 67116 13858 67172 14140
rect 67228 14196 67284 17724
rect 67564 16996 67620 17006
rect 67564 16902 67620 16940
rect 67340 16882 67396 16894
rect 67340 16830 67342 16882
rect 67394 16830 67396 16882
rect 67340 16100 67396 16830
rect 67452 16884 67508 16894
rect 67452 16790 67508 16828
rect 67340 16034 67396 16044
rect 67900 15316 67956 15326
rect 67676 14644 67732 14654
rect 67676 14530 67732 14588
rect 67900 14642 67956 15260
rect 67900 14590 67902 14642
rect 67954 14590 67956 14642
rect 67900 14578 67956 14590
rect 67676 14478 67678 14530
rect 67730 14478 67732 14530
rect 67676 14466 67732 14478
rect 68012 14532 68068 14542
rect 68012 14438 68068 14476
rect 67228 14130 67284 14140
rect 67452 14084 67508 14094
rect 67228 13972 67284 13982
rect 67228 13878 67284 13916
rect 67452 13970 67508 14028
rect 67452 13918 67454 13970
rect 67506 13918 67508 13970
rect 67452 13906 67508 13918
rect 67788 13972 67844 13982
rect 67788 13878 67844 13916
rect 67116 13806 67118 13858
rect 67170 13806 67172 13858
rect 67116 13794 67172 13806
rect 68012 13636 68068 13646
rect 67004 13188 67060 13198
rect 67004 12404 67060 13132
rect 67228 13076 67284 13086
rect 67228 12982 67284 13020
rect 67900 12964 67956 12974
rect 67900 12870 67956 12908
rect 67004 12338 67060 12348
rect 67004 12180 67060 12190
rect 67676 12180 67732 12190
rect 67004 12178 67172 12180
rect 67004 12126 67006 12178
rect 67058 12126 67172 12178
rect 67004 12124 67172 12126
rect 67004 12114 67060 12124
rect 67004 11956 67060 11966
rect 67004 11506 67060 11900
rect 67004 11454 67006 11506
rect 67058 11454 67060 11506
rect 67004 11442 67060 11454
rect 67116 10612 67172 12124
rect 67452 12178 67732 12180
rect 67452 12126 67678 12178
rect 67730 12126 67732 12178
rect 67452 12124 67732 12126
rect 67452 11956 67508 12124
rect 67676 12114 67732 12124
rect 67452 11506 67508 11900
rect 67452 11454 67454 11506
rect 67506 11454 67508 11506
rect 67452 11442 67508 11454
rect 67452 11172 67508 11182
rect 67340 10612 67396 10622
rect 67116 10556 67340 10612
rect 67340 10518 67396 10556
rect 67004 10500 67060 10510
rect 67004 9826 67060 10444
rect 67340 10276 67396 10286
rect 67004 9774 67006 9826
rect 67058 9774 67060 9826
rect 67004 9762 67060 9774
rect 67228 9938 67284 9950
rect 67228 9886 67230 9938
rect 67282 9886 67284 9938
rect 67228 9266 67284 9886
rect 67228 9214 67230 9266
rect 67282 9214 67284 9266
rect 67228 9202 67284 9214
rect 66892 8372 67060 8428
rect 66780 8094 66782 8146
rect 66834 8094 66836 8146
rect 66780 8082 66836 8094
rect 67004 8036 67060 8372
rect 67004 8034 67172 8036
rect 67004 7982 67006 8034
rect 67058 7982 67172 8034
rect 67004 7980 67172 7982
rect 67004 7970 67060 7980
rect 65772 7698 65940 7700
rect 65772 7646 65774 7698
rect 65826 7646 65940 7698
rect 65772 7644 65940 7646
rect 66556 7924 66612 7934
rect 66556 7700 66612 7868
rect 66556 7698 66724 7700
rect 66556 7646 66558 7698
rect 66610 7646 66724 7698
rect 66556 7644 66724 7646
rect 65772 7634 65828 7644
rect 66556 7634 66612 7644
rect 66108 7476 66164 7486
rect 66108 7382 66164 7420
rect 65660 7074 65716 7084
rect 65324 6972 65604 7028
rect 65212 6402 65268 6412
rect 64988 6178 65044 6188
rect 64876 5182 64878 5234
rect 64930 5182 64932 5234
rect 64876 5170 64932 5182
rect 65436 5908 65492 5918
rect 65436 5010 65492 5852
rect 65548 5794 65604 6972
rect 66444 6916 66500 6926
rect 66444 6822 66500 6860
rect 65772 6802 65828 6814
rect 65772 6750 65774 6802
rect 65826 6750 65828 6802
rect 65660 6692 65716 6702
rect 65660 6598 65716 6636
rect 65548 5742 65550 5794
rect 65602 5742 65604 5794
rect 65548 5730 65604 5742
rect 65772 6468 65828 6750
rect 65436 4958 65438 5010
rect 65490 4958 65492 5010
rect 64316 2706 64372 2716
rect 64428 3554 64820 3556
rect 64428 3502 64766 3554
rect 64818 3502 64820 3554
rect 64428 3500 64820 3502
rect 64428 800 64484 3500
rect 64764 3490 64820 3500
rect 65100 4900 65156 4910
rect 65100 3666 65156 4844
rect 65100 3614 65102 3666
rect 65154 3614 65156 3666
rect 65100 1540 65156 3614
rect 65100 1474 65156 1484
rect 65436 1428 65492 4958
rect 65548 5236 65604 5246
rect 65548 5010 65604 5180
rect 65548 4958 65550 5010
rect 65602 4958 65604 5010
rect 65548 4946 65604 4958
rect 65660 5124 65716 5134
rect 65660 4338 65716 5068
rect 65772 5122 65828 6412
rect 66668 6356 66724 7644
rect 66556 6244 66612 6254
rect 66556 6020 66612 6188
rect 65884 5908 65940 5946
rect 66556 5926 66612 5964
rect 66668 6130 66724 6300
rect 66668 6078 66670 6130
rect 66722 6078 66724 6130
rect 65884 5842 65940 5852
rect 65772 5070 65774 5122
rect 65826 5070 65828 5122
rect 65772 5058 65828 5070
rect 65884 5684 65940 5694
rect 65660 4286 65662 4338
rect 65714 4286 65716 4338
rect 65660 4274 65716 4286
rect 65884 4226 65940 5628
rect 66332 5348 66388 5358
rect 65884 4174 65886 4226
rect 65938 4174 65940 4226
rect 65884 4162 65940 4174
rect 66108 5236 66164 5246
rect 65660 3444 65716 3454
rect 66108 3444 66164 5180
rect 66220 5010 66276 5022
rect 66220 4958 66222 5010
rect 66274 4958 66276 5010
rect 66220 4788 66276 4958
rect 66332 4900 66388 5292
rect 66668 5236 66724 6078
rect 67004 6466 67060 6478
rect 67004 6414 67006 6466
rect 67058 6414 67060 6466
rect 66892 5908 66948 5918
rect 66892 5814 66948 5852
rect 67004 5348 67060 6414
rect 67116 6020 67172 7980
rect 67340 7700 67396 10220
rect 67452 9380 67508 11116
rect 67564 10498 67620 10510
rect 67564 10446 67566 10498
rect 67618 10446 67620 10498
rect 67564 10388 67620 10446
rect 67564 10050 67620 10332
rect 67564 9998 67566 10050
rect 67618 9998 67620 10050
rect 67564 9986 67620 9998
rect 68012 9828 68068 13580
rect 68124 13412 68180 18508
rect 68236 14420 68292 20132
rect 69020 20020 69076 20030
rect 69020 19926 69076 19964
rect 68684 19908 68740 19918
rect 68684 19814 68740 19852
rect 68832 19628 69096 19638
rect 68888 19572 68936 19628
rect 68992 19572 69040 19628
rect 68832 19562 69096 19572
rect 68572 19012 68628 19022
rect 68684 19012 68740 19022
rect 68572 19010 68684 19012
rect 68572 18958 68574 19010
rect 68626 18958 68684 19010
rect 68572 18956 68684 18958
rect 68572 18946 68628 18956
rect 68348 18340 68404 18350
rect 68348 17780 68404 18284
rect 68348 17714 68404 17724
rect 68236 14354 68292 14364
rect 68348 14418 68404 14430
rect 68348 14366 68350 14418
rect 68402 14366 68404 14418
rect 68236 14196 68292 14206
rect 68236 13860 68292 14140
rect 68236 13766 68292 13804
rect 68124 13356 68292 13412
rect 68124 13076 68180 13086
rect 68124 12962 68180 13020
rect 68124 12910 68126 12962
rect 68178 12910 68180 12962
rect 68124 12292 68180 12910
rect 68124 12226 68180 12236
rect 68236 12404 68292 13356
rect 68348 13188 68404 14366
rect 68460 13188 68516 13198
rect 68348 13186 68516 13188
rect 68348 13134 68462 13186
rect 68514 13134 68516 13186
rect 68348 13132 68516 13134
rect 68460 13122 68516 13132
rect 68236 12178 68292 12348
rect 68236 12126 68238 12178
rect 68290 12126 68292 12178
rect 68236 12114 68292 12126
rect 68572 10612 68628 10650
rect 68572 10546 68628 10556
rect 68348 10500 68404 10510
rect 68236 10388 68292 10398
rect 68236 10294 68292 10332
rect 68348 9940 68404 10444
rect 68572 10388 68628 10398
rect 68572 10294 68628 10332
rect 68348 9938 68516 9940
rect 68348 9886 68350 9938
rect 68402 9886 68516 9938
rect 68348 9884 68516 9886
rect 68348 9874 68404 9884
rect 67788 9772 68068 9828
rect 67452 9324 67620 9380
rect 67564 9268 67620 9324
rect 67452 9156 67508 9166
rect 67452 9062 67508 9100
rect 67564 9154 67620 9212
rect 67564 9102 67566 9154
rect 67618 9102 67620 9154
rect 67564 9090 67620 9102
rect 67564 8372 67620 8382
rect 67452 7700 67508 7710
rect 67340 7644 67452 7700
rect 67452 7568 67508 7644
rect 67564 7588 67620 8316
rect 67564 7522 67620 7532
rect 67340 7476 67396 7486
rect 67340 7382 67396 7420
rect 67676 7476 67732 7486
rect 67676 7382 67732 7420
rect 67676 7140 67732 7150
rect 67676 6466 67732 7084
rect 67788 6690 67844 9772
rect 68236 9156 68292 9166
rect 67900 9154 68292 9156
rect 67900 9102 68238 9154
rect 68290 9102 68292 9154
rect 67900 9100 68292 9102
rect 67900 7924 67956 9100
rect 68236 9090 68292 9100
rect 68348 9044 68404 9054
rect 68348 8950 68404 8988
rect 67900 7858 67956 7868
rect 68012 8932 68068 8942
rect 68012 8034 68068 8876
rect 68236 8820 68292 8830
rect 68460 8820 68516 9884
rect 68236 8818 68516 8820
rect 68236 8766 68238 8818
rect 68290 8766 68516 8818
rect 68236 8764 68516 8766
rect 68236 8754 68292 8764
rect 68684 8428 68740 18956
rect 68908 18562 68964 18574
rect 68908 18510 68910 18562
rect 68962 18510 68964 18562
rect 68908 18340 68964 18510
rect 68908 18274 68964 18284
rect 69244 18340 69300 20860
rect 69356 20690 69412 20702
rect 69356 20638 69358 20690
rect 69410 20638 69412 20690
rect 69356 19908 69412 20638
rect 69468 20580 69524 21422
rect 69804 21474 69860 21486
rect 69804 21422 69806 21474
rect 69858 21422 69860 21474
rect 69580 20916 69636 20926
rect 69580 20802 69636 20860
rect 69804 20804 69860 21422
rect 70812 21474 70868 21486
rect 70812 21422 70814 21474
rect 70866 21422 70868 21474
rect 69916 21028 69972 21038
rect 69916 20934 69972 20972
rect 70812 21028 70868 21422
rect 70812 20962 70868 20972
rect 71036 20914 71092 22092
rect 71484 22092 71652 22148
rect 71036 20862 71038 20914
rect 71090 20862 71092 20914
rect 71036 20850 71092 20862
rect 71148 21586 71204 21598
rect 71148 21534 71150 21586
rect 71202 21534 71204 21586
rect 69580 20750 69582 20802
rect 69634 20750 69636 20802
rect 69580 20738 69636 20750
rect 69692 20748 69804 20804
rect 69468 20514 69524 20524
rect 69356 19842 69412 19852
rect 69468 20356 69524 20366
rect 69468 19458 69524 20300
rect 69692 20188 69748 20748
rect 69804 20738 69860 20748
rect 70364 20804 70420 20814
rect 70364 20710 70420 20748
rect 70812 20690 70868 20702
rect 70812 20638 70814 20690
rect 70866 20638 70868 20690
rect 69804 20580 69860 20590
rect 70476 20580 70532 20590
rect 69860 20524 69972 20580
rect 69804 20486 69860 20524
rect 69468 19406 69470 19458
rect 69522 19406 69524 19458
rect 69468 19394 69524 19406
rect 69580 20132 69748 20188
rect 69356 19124 69412 19134
rect 69356 19030 69412 19068
rect 69468 19012 69524 19022
rect 69468 18918 69524 18956
rect 69356 18340 69412 18350
rect 69244 18338 69412 18340
rect 69244 18286 69358 18338
rect 69410 18286 69412 18338
rect 69244 18284 69412 18286
rect 68832 18060 69096 18070
rect 68888 18004 68936 18060
rect 68992 18004 69040 18060
rect 68832 17994 69096 18004
rect 68832 16492 69096 16502
rect 68888 16436 68936 16492
rect 68992 16436 69040 16492
rect 68832 16426 69096 16436
rect 69244 15876 69300 18284
rect 69356 18274 69412 18284
rect 69580 18228 69636 20132
rect 69916 20020 69972 20524
rect 69916 19954 69972 19964
rect 70028 20132 70084 20142
rect 69580 18162 69636 18172
rect 69692 19908 69748 19918
rect 69692 17780 69748 19852
rect 70028 18562 70084 20076
rect 70364 20132 70420 20142
rect 70476 20132 70532 20524
rect 70364 20130 70532 20132
rect 70364 20078 70366 20130
rect 70418 20078 70532 20130
rect 70364 20076 70532 20078
rect 70364 20066 70420 20076
rect 70812 20020 70868 20638
rect 70924 20580 70980 20590
rect 70924 20486 70980 20524
rect 71148 20578 71204 21534
rect 71148 20526 71150 20578
rect 71202 20526 71204 20578
rect 71148 20468 71204 20526
rect 71148 20402 71204 20412
rect 70252 19908 70308 19918
rect 70252 19814 70308 19852
rect 70476 19346 70532 19358
rect 70476 19294 70478 19346
rect 70530 19294 70532 19346
rect 70364 19234 70420 19246
rect 70364 19182 70366 19234
rect 70418 19182 70420 19234
rect 70364 19012 70420 19182
rect 70476 19124 70532 19294
rect 70476 19058 70532 19068
rect 70364 18946 70420 18956
rect 70028 18510 70030 18562
rect 70082 18510 70084 18562
rect 70028 18498 70084 18510
rect 70140 18564 70196 18574
rect 70140 18004 70196 18508
rect 70700 18452 70756 18462
rect 70700 18358 70756 18396
rect 69580 17724 69748 17780
rect 70028 17948 70196 18004
rect 69356 17668 69412 17678
rect 69356 17574 69412 17612
rect 69468 16884 69524 16894
rect 69468 16790 69524 16828
rect 69244 15810 69300 15820
rect 69468 16660 69524 16670
rect 68908 15652 68964 15662
rect 68908 15314 68964 15596
rect 69468 15538 69524 16604
rect 69468 15486 69470 15538
rect 69522 15486 69524 15538
rect 69468 15428 69524 15486
rect 69468 15362 69524 15372
rect 68908 15262 68910 15314
rect 68962 15262 68964 15314
rect 68908 15250 68964 15262
rect 68832 14924 69096 14934
rect 68888 14868 68936 14924
rect 68992 14868 69040 14924
rect 68832 14858 69096 14868
rect 69356 13748 69412 13758
rect 68832 13356 69096 13366
rect 68888 13300 68936 13356
rect 68992 13300 69040 13356
rect 68832 13290 69096 13300
rect 69244 12738 69300 12750
rect 69244 12686 69246 12738
rect 69298 12686 69300 12738
rect 68796 12292 68852 12302
rect 68796 12198 68852 12236
rect 69244 12292 69300 12686
rect 69244 12226 69300 12236
rect 68832 11788 69096 11798
rect 68888 11732 68936 11788
rect 68992 11732 69040 11788
rect 68832 11722 69096 11732
rect 69356 11060 69412 13692
rect 69580 12068 69636 17724
rect 69804 17668 69860 17678
rect 69692 17556 69748 17566
rect 69692 16882 69748 17500
rect 69692 16830 69694 16882
rect 69746 16830 69748 16882
rect 69692 16818 69748 16830
rect 69804 16884 69860 17612
rect 70028 17106 70084 17948
rect 70140 17778 70196 17790
rect 70140 17726 70142 17778
rect 70194 17726 70196 17778
rect 70140 17556 70196 17726
rect 70140 17490 70196 17500
rect 70364 17556 70420 17566
rect 70028 17054 70030 17106
rect 70082 17054 70084 17106
rect 70028 17042 70084 17054
rect 70252 17444 70308 17454
rect 69804 16818 69860 16828
rect 69916 16100 69972 16110
rect 69916 16098 70084 16100
rect 69916 16046 69918 16098
rect 69970 16046 70084 16098
rect 69916 16044 70084 16046
rect 69916 16034 69972 16044
rect 69916 15428 69972 15438
rect 69692 14642 69748 14654
rect 69692 14590 69694 14642
rect 69746 14590 69748 14642
rect 69692 14084 69748 14590
rect 69692 14018 69748 14028
rect 69804 13634 69860 13646
rect 69804 13582 69806 13634
rect 69858 13582 69860 13634
rect 69804 13188 69860 13582
rect 69804 13122 69860 13132
rect 69580 11974 69636 12012
rect 69916 11396 69972 15372
rect 70028 15316 70084 16044
rect 70028 15250 70084 15260
rect 70140 16098 70196 16110
rect 70140 16046 70142 16098
rect 70194 16046 70196 16098
rect 70140 15204 70196 16046
rect 70252 15538 70308 17388
rect 70364 16210 70420 17500
rect 70812 17332 70868 19964
rect 71260 20020 71316 20030
rect 71260 19234 71316 19964
rect 71260 19182 71262 19234
rect 71314 19182 71316 19234
rect 71260 19170 71316 19182
rect 71484 18676 71540 22092
rect 73276 22036 73332 22988
rect 73388 23154 73444 23166
rect 73388 23102 73390 23154
rect 73442 23102 73444 23154
rect 73388 22484 73444 23102
rect 73612 23156 73668 23166
rect 73612 23062 73668 23100
rect 73388 22418 73444 22428
rect 73276 21970 73332 21980
rect 72156 21812 72212 21822
rect 71708 21700 71764 21710
rect 71708 21606 71764 21644
rect 72156 20914 72212 21756
rect 73724 21588 73780 34636
rect 73948 33570 74004 34860
rect 74060 34244 74116 34254
rect 74396 34244 74452 34254
rect 74060 34150 74116 34188
rect 74172 34242 74452 34244
rect 74172 34190 74398 34242
rect 74450 34190 74452 34242
rect 74172 34188 74452 34190
rect 73948 33518 73950 33570
rect 74002 33518 74004 33570
rect 73948 33506 74004 33518
rect 73948 33348 74004 33358
rect 73948 33254 74004 33292
rect 74172 31948 74228 34188
rect 74396 34178 74452 34188
rect 74508 34132 74564 35756
rect 74956 35698 75012 36204
rect 75180 36260 75236 36270
rect 75180 36258 75348 36260
rect 75180 36206 75182 36258
rect 75234 36206 75348 36258
rect 75180 36204 75348 36206
rect 75180 36194 75236 36204
rect 74956 35646 74958 35698
rect 75010 35646 75012 35698
rect 74956 35634 75012 35646
rect 74956 34916 75012 34926
rect 74956 34822 75012 34860
rect 74956 34132 75012 34142
rect 74508 34130 75012 34132
rect 74508 34078 74958 34130
rect 75010 34078 75012 34130
rect 74508 34076 75012 34078
rect 74956 34066 75012 34076
rect 74396 33570 74452 33582
rect 74396 33518 74398 33570
rect 74450 33518 74452 33570
rect 74396 33458 74452 33518
rect 74396 33406 74398 33458
rect 74450 33406 74452 33458
rect 74396 33394 74452 33406
rect 75068 33348 75124 33358
rect 74732 33346 75124 33348
rect 74732 33294 75070 33346
rect 75122 33294 75124 33346
rect 74732 33292 75124 33294
rect 74284 32788 74340 32798
rect 74284 32694 74340 32732
rect 74732 32674 74788 33292
rect 75068 33282 75124 33292
rect 74844 33124 74900 33134
rect 74844 33030 74900 33068
rect 74732 32622 74734 32674
rect 74786 32622 74788 32674
rect 74732 32610 74788 32622
rect 74844 32564 74900 32574
rect 74844 32470 74900 32508
rect 75180 32562 75236 32574
rect 75180 32510 75182 32562
rect 75234 32510 75236 32562
rect 75180 31948 75236 32510
rect 74060 31892 74228 31948
rect 74284 31892 75236 31948
rect 73836 28868 73892 28878
rect 73836 28754 73892 28812
rect 73836 28702 73838 28754
rect 73890 28702 73892 28754
rect 73836 28690 73892 28702
rect 73836 26964 73892 26974
rect 73836 26402 73892 26908
rect 73836 26350 73838 26402
rect 73890 26350 73892 26402
rect 73836 26338 73892 26350
rect 73948 26628 74004 26638
rect 73948 24388 74004 26572
rect 74060 24836 74116 31892
rect 74284 31890 74340 31892
rect 74284 31838 74286 31890
rect 74338 31838 74340 31890
rect 74284 31826 74340 31838
rect 74396 31666 74452 31678
rect 74396 31614 74398 31666
rect 74450 31614 74452 31666
rect 74172 31554 74228 31566
rect 74172 31502 74174 31554
rect 74226 31502 74228 31554
rect 74172 29988 74228 31502
rect 74396 31556 74452 31614
rect 74396 31490 74452 31500
rect 74620 31220 74676 31230
rect 74620 31126 74676 31164
rect 74844 31106 74900 31118
rect 74844 31054 74846 31106
rect 74898 31054 74900 31106
rect 74396 30324 74452 30334
rect 74396 30230 74452 30268
rect 74508 30324 74564 30334
rect 74844 30324 74900 31054
rect 74508 30322 74900 30324
rect 74508 30270 74510 30322
rect 74562 30270 74900 30322
rect 74508 30268 74900 30270
rect 74956 30994 75012 31006
rect 74956 30942 74958 30994
rect 75010 30942 75012 30994
rect 74172 29922 74228 29932
rect 74284 29986 74340 29998
rect 74284 29934 74286 29986
rect 74338 29934 74340 29986
rect 74284 29876 74340 29934
rect 74284 29810 74340 29820
rect 74508 28868 74564 30268
rect 74956 30100 75012 30942
rect 75068 30212 75124 30222
rect 75068 30118 75124 30156
rect 74956 30034 75012 30044
rect 74508 28802 74564 28812
rect 74844 29876 74900 29886
rect 74620 28754 74676 28766
rect 74620 28702 74622 28754
rect 74674 28702 74676 28754
rect 74508 28642 74564 28654
rect 74508 28590 74510 28642
rect 74562 28590 74564 28642
rect 74508 27972 74564 28590
rect 74508 27906 74564 27916
rect 74172 27860 74228 27870
rect 74172 27746 74228 27804
rect 74172 27694 74174 27746
rect 74226 27694 74228 27746
rect 74172 27188 74228 27694
rect 74508 27748 74564 27758
rect 74620 27748 74676 28702
rect 74508 27746 74676 27748
rect 74508 27694 74510 27746
rect 74562 27694 74676 27746
rect 74508 27692 74676 27694
rect 74508 27524 74564 27692
rect 74508 27458 74564 27468
rect 74172 27132 74676 27188
rect 74172 26962 74228 26974
rect 74172 26910 74174 26962
rect 74226 26910 74228 26962
rect 74172 26628 74228 26910
rect 74620 26908 74676 27132
rect 74844 27186 74900 29820
rect 75068 29764 75124 29774
rect 75068 28082 75124 29708
rect 75180 29428 75236 29438
rect 75292 29428 75348 36204
rect 75740 36036 75796 36046
rect 75628 33460 75684 33470
rect 75628 33366 75684 33404
rect 75740 32788 75796 35980
rect 76300 36036 76356 36430
rect 76300 35970 76356 35980
rect 76076 35924 76132 35934
rect 76076 35810 76132 35868
rect 76076 35758 76078 35810
rect 76130 35758 76132 35810
rect 76076 35746 76132 35758
rect 76748 35812 76804 35822
rect 76748 35698 76804 35756
rect 76748 35646 76750 35698
rect 76802 35646 76804 35698
rect 76748 35634 76804 35646
rect 76076 35028 76132 35038
rect 76076 34934 76132 34972
rect 77084 34804 77140 37324
rect 77868 35810 77924 38444
rect 77980 36596 78036 36606
rect 77980 36502 78036 36540
rect 77868 35758 77870 35810
rect 77922 35758 77924 35810
rect 77868 35746 77924 35758
rect 77532 35252 77588 35262
rect 76748 34244 76804 34254
rect 76748 34150 76804 34188
rect 77084 34242 77140 34748
rect 77084 34190 77086 34242
rect 77138 34190 77140 34242
rect 77084 34178 77140 34190
rect 77308 34802 77364 34814
rect 77308 34750 77310 34802
rect 77362 34750 77364 34802
rect 76076 34018 76132 34030
rect 76076 33966 76078 34018
rect 76130 33966 76132 34018
rect 76076 33684 76132 33966
rect 76076 33618 76132 33628
rect 76412 33460 76468 33470
rect 76412 33346 76468 33404
rect 76412 33294 76414 33346
rect 76466 33294 76468 33346
rect 76412 33282 76468 33294
rect 77308 33348 77364 34750
rect 77532 34132 77588 35196
rect 77980 35140 78036 35150
rect 77644 34692 77700 34702
rect 77644 34690 77924 34692
rect 77644 34638 77646 34690
rect 77698 34638 77924 34690
rect 77644 34636 77924 34638
rect 77644 34626 77700 34636
rect 77644 34244 77700 34254
rect 77644 34242 77812 34244
rect 77644 34190 77646 34242
rect 77698 34190 77812 34242
rect 77644 34188 77812 34190
rect 77644 34178 77700 34188
rect 77532 34066 77588 34076
rect 77308 33282 77364 33292
rect 77532 33346 77588 33358
rect 77532 33294 77534 33346
rect 77586 33294 77588 33346
rect 75740 32722 75796 32732
rect 76188 33122 76244 33134
rect 76188 33070 76190 33122
rect 76242 33070 76244 33122
rect 75516 31890 75572 31902
rect 75516 31838 75518 31890
rect 75570 31838 75572 31890
rect 75404 31556 75460 31566
rect 75404 30884 75460 31500
rect 75516 31108 75572 31838
rect 76188 31778 76244 33070
rect 77308 33124 77364 33134
rect 77308 33122 77476 33124
rect 77308 33070 77310 33122
rect 77362 33070 77476 33122
rect 77308 33068 77476 33070
rect 77308 33058 77364 33068
rect 76524 32674 76580 32686
rect 76524 32622 76526 32674
rect 76578 32622 76580 32674
rect 76188 31726 76190 31778
rect 76242 31726 76244 31778
rect 76188 31714 76244 31726
rect 76300 32338 76356 32350
rect 76300 32286 76302 32338
rect 76354 32286 76356 32338
rect 76300 31220 76356 32286
rect 76300 31154 76356 31164
rect 75516 31042 75572 31052
rect 75964 30994 76020 31006
rect 75964 30942 75966 30994
rect 76018 30942 76020 30994
rect 75516 30884 75572 30894
rect 75404 30882 75572 30884
rect 75404 30830 75518 30882
rect 75570 30830 75572 30882
rect 75404 30828 75572 30830
rect 75516 30818 75572 30828
rect 75964 30772 76020 30942
rect 75964 30706 76020 30716
rect 76076 30994 76132 31006
rect 76076 30942 76078 30994
rect 76130 30942 76132 30994
rect 75404 30324 75460 30334
rect 75404 30230 75460 30268
rect 75516 30212 75572 30222
rect 75516 30118 75572 30156
rect 76076 30212 76132 30942
rect 76076 30146 76132 30156
rect 76188 30994 76244 31006
rect 76188 30942 76190 30994
rect 76242 30942 76244 30994
rect 76188 29876 76244 30942
rect 76188 29810 76244 29820
rect 76412 30434 76468 30446
rect 76412 30382 76414 30434
rect 76466 30382 76468 30434
rect 75180 29426 75348 29428
rect 75180 29374 75182 29426
rect 75234 29374 75348 29426
rect 75180 29372 75348 29374
rect 75180 29362 75236 29372
rect 76076 29314 76132 29326
rect 76076 29262 76078 29314
rect 76130 29262 76132 29314
rect 75516 28756 75572 28766
rect 75404 28644 75460 28654
rect 75404 28550 75460 28588
rect 75068 28030 75070 28082
rect 75122 28030 75124 28082
rect 75068 28018 75124 28030
rect 75516 27970 75572 28700
rect 76076 28644 76132 29262
rect 76076 28578 76132 28588
rect 76188 28754 76244 28766
rect 76188 28702 76190 28754
rect 76242 28702 76244 28754
rect 76188 28196 76244 28702
rect 76300 28756 76356 28766
rect 76300 28642 76356 28700
rect 76300 28590 76302 28642
rect 76354 28590 76356 28642
rect 76300 28578 76356 28590
rect 76412 28308 76468 30382
rect 76524 30100 76580 32622
rect 77196 32674 77252 32686
rect 77196 32622 77198 32674
rect 77250 32622 77252 32674
rect 76636 32338 76692 32350
rect 76636 32286 76638 32338
rect 76690 32286 76692 32338
rect 76636 31892 76692 32286
rect 76636 31826 76692 31836
rect 76860 31108 76916 31118
rect 76748 31106 76916 31108
rect 76748 31054 76862 31106
rect 76914 31054 76916 31106
rect 76748 31052 76916 31054
rect 76748 30434 76804 31052
rect 76860 31042 76916 31052
rect 77084 30996 77140 31006
rect 77084 30902 77140 30940
rect 76748 30382 76750 30434
rect 76802 30382 76804 30434
rect 76748 30370 76804 30382
rect 76524 30034 76580 30044
rect 76636 29986 76692 29998
rect 76636 29934 76638 29986
rect 76690 29934 76692 29986
rect 76636 29540 76692 29934
rect 76636 29484 77028 29540
rect 76748 29316 76804 29326
rect 76188 28130 76244 28140
rect 76300 28252 76468 28308
rect 76636 29314 76804 29316
rect 76636 29262 76750 29314
rect 76802 29262 76804 29314
rect 76636 29260 76804 29262
rect 76636 29202 76692 29260
rect 76748 29250 76804 29260
rect 76972 29316 77028 29484
rect 77084 29316 77140 29326
rect 76972 29314 77140 29316
rect 76972 29262 77086 29314
rect 77138 29262 77140 29314
rect 76972 29260 77140 29262
rect 76636 29150 76638 29202
rect 76690 29150 76692 29202
rect 75516 27918 75518 27970
rect 75570 27918 75572 27970
rect 75516 27906 75572 27918
rect 75740 27972 75796 27982
rect 75740 27878 75796 27916
rect 75628 27858 75684 27870
rect 75628 27806 75630 27858
rect 75682 27806 75684 27858
rect 75628 27524 75684 27806
rect 75628 27458 75684 27468
rect 74844 27134 74846 27186
rect 74898 27134 74900 27186
rect 74844 27122 74900 27134
rect 76188 27188 76244 27198
rect 75628 27074 75684 27086
rect 75628 27022 75630 27074
rect 75682 27022 75684 27074
rect 74172 26562 74228 26572
rect 74508 26852 74676 26908
rect 74732 26962 74788 26974
rect 74732 26910 74734 26962
rect 74786 26910 74788 26962
rect 74284 26516 74340 26526
rect 74172 26292 74228 26302
rect 74172 26198 74228 26236
rect 74284 26068 74340 26460
rect 74284 26002 74340 26012
rect 74396 26290 74452 26302
rect 74396 26238 74398 26290
rect 74450 26238 74452 26290
rect 74396 25956 74452 26238
rect 74396 25890 74452 25900
rect 74060 24780 74228 24836
rect 74060 24612 74116 24622
rect 74060 24518 74116 24556
rect 73948 24332 74116 24388
rect 73948 23154 74004 23166
rect 73948 23102 73950 23154
rect 74002 23102 74004 23154
rect 73948 22596 74004 23102
rect 73948 22530 74004 22540
rect 73724 21522 73780 21532
rect 72156 20862 72158 20914
rect 72210 20862 72212 20914
rect 72156 20850 72212 20862
rect 72716 20916 72772 20926
rect 72716 20822 72772 20860
rect 74060 20914 74116 24332
rect 74172 21028 74228 24780
rect 74396 22370 74452 22382
rect 74396 22318 74398 22370
rect 74450 22318 74452 22370
rect 74396 22260 74452 22318
rect 74396 22194 74452 22204
rect 74396 21588 74452 21598
rect 74396 21494 74452 21532
rect 74172 20962 74228 20972
rect 74060 20862 74062 20914
rect 74114 20862 74116 20914
rect 74060 20850 74116 20862
rect 71596 20802 71652 20814
rect 71596 20750 71598 20802
rect 71650 20750 71652 20802
rect 71596 20356 71652 20750
rect 73724 20804 73780 20814
rect 73724 20710 73780 20748
rect 74284 20802 74340 20814
rect 74284 20750 74286 20802
rect 74338 20750 74340 20802
rect 71596 20290 71652 20300
rect 71708 20692 71764 20702
rect 71708 20018 71764 20636
rect 72268 20692 72324 20702
rect 72268 20598 72324 20636
rect 73836 20690 73892 20702
rect 73836 20638 73838 20690
rect 73890 20638 73892 20690
rect 71708 19966 71710 20018
rect 71762 19966 71764 20018
rect 71708 19954 71764 19966
rect 72044 20578 72100 20590
rect 72044 20526 72046 20578
rect 72098 20526 72100 20578
rect 72044 20020 72100 20526
rect 72044 19954 72100 19964
rect 71932 19908 71988 19918
rect 71932 19814 71988 19852
rect 72492 19908 72548 19918
rect 72044 19796 72100 19806
rect 71708 19012 71764 19022
rect 71708 18918 71764 18956
rect 71708 18676 71764 18686
rect 71484 18674 71764 18676
rect 71484 18622 71710 18674
rect 71762 18622 71764 18674
rect 71484 18620 71764 18622
rect 71708 18610 71764 18620
rect 71372 18564 71428 18574
rect 71428 18508 71652 18564
rect 71372 18498 71428 18508
rect 71596 18450 71652 18508
rect 71596 18398 71598 18450
rect 71650 18398 71652 18450
rect 71596 18386 71652 18398
rect 71820 18450 71876 18462
rect 71820 18398 71822 18450
rect 71874 18398 71876 18450
rect 70924 18338 70980 18350
rect 70924 18286 70926 18338
rect 70978 18286 70980 18338
rect 70924 17780 70980 18286
rect 71148 17780 71204 17790
rect 70924 17778 71204 17780
rect 70924 17726 71150 17778
rect 71202 17726 71204 17778
rect 70924 17724 71204 17726
rect 71148 17714 71204 17724
rect 71260 17668 71316 17678
rect 71260 17574 71316 17612
rect 71484 17668 71540 17678
rect 71820 17668 71876 18398
rect 72044 18228 72100 19740
rect 72156 18452 72212 18462
rect 72156 18358 72212 18396
rect 72044 18172 72212 18228
rect 71484 17666 71876 17668
rect 71484 17614 71486 17666
rect 71538 17614 71876 17666
rect 71484 17612 71876 17614
rect 71036 17556 71092 17566
rect 71036 17462 71092 17500
rect 71484 17444 71540 17612
rect 71484 17378 71540 17388
rect 70812 17276 71092 17332
rect 70364 16158 70366 16210
rect 70418 16158 70420 16210
rect 70364 16146 70420 16158
rect 70812 15874 70868 15886
rect 70812 15822 70814 15874
rect 70866 15822 70868 15874
rect 70812 15652 70868 15822
rect 70924 15652 70980 15662
rect 70812 15596 70924 15652
rect 70252 15486 70254 15538
rect 70306 15486 70308 15538
rect 70252 15474 70308 15486
rect 70924 15426 70980 15596
rect 71036 15540 71092 17276
rect 71260 15874 71316 15886
rect 71260 15822 71262 15874
rect 71314 15822 71316 15874
rect 71260 15540 71316 15822
rect 71092 15484 71316 15540
rect 71036 15446 71092 15484
rect 70924 15374 70926 15426
rect 70978 15374 70980 15426
rect 70924 15362 70980 15374
rect 71596 15428 71652 15438
rect 71596 15334 71652 15372
rect 71260 15314 71316 15326
rect 71260 15262 71262 15314
rect 71314 15262 71316 15314
rect 70364 15204 70420 15214
rect 70140 15202 70420 15204
rect 70140 15150 70366 15202
rect 70418 15150 70420 15202
rect 70140 15148 70420 15150
rect 70364 15092 70420 15148
rect 70364 15026 70420 15036
rect 70028 14756 70084 14766
rect 70028 14530 70084 14700
rect 71260 14756 71316 15262
rect 71260 14690 71316 14700
rect 71820 14756 71876 14766
rect 70028 14478 70030 14530
rect 70082 14478 70084 14530
rect 70028 14466 70084 14478
rect 70476 14532 70532 14542
rect 70476 14438 70532 14476
rect 71484 14532 71540 14542
rect 71484 14438 71540 14476
rect 71708 14530 71764 14542
rect 71708 14478 71710 14530
rect 71762 14478 71764 14530
rect 71708 14196 71764 14478
rect 71372 14140 71764 14196
rect 70140 13860 70196 13870
rect 70140 12852 70196 13804
rect 70364 13636 70420 13646
rect 70364 13542 70420 13580
rect 70812 13636 70868 13646
rect 70812 13542 70868 13580
rect 71372 13636 71428 14140
rect 71708 13860 71764 13870
rect 71484 13748 71540 13758
rect 71484 13654 71540 13692
rect 71372 13542 71428 13580
rect 70140 12758 70196 12796
rect 70252 13188 70308 13198
rect 70252 12850 70308 13132
rect 71708 13074 71764 13804
rect 71708 13022 71710 13074
rect 71762 13022 71764 13074
rect 71708 13010 71764 13022
rect 70252 12798 70254 12850
rect 70306 12798 70308 12850
rect 70252 12786 70308 12798
rect 71148 12962 71204 12974
rect 71148 12910 71150 12962
rect 71202 12910 71204 12962
rect 70476 12740 70532 12750
rect 70476 12646 70532 12684
rect 71148 12740 71204 12910
rect 70476 12178 70532 12190
rect 70476 12126 70478 12178
rect 70530 12126 70532 12178
rect 70028 12068 70084 12078
rect 70028 11618 70084 12012
rect 70364 12068 70420 12078
rect 70364 11974 70420 12012
rect 70028 11566 70030 11618
rect 70082 11566 70084 11618
rect 70028 11554 70084 11566
rect 70140 11396 70196 11406
rect 69916 11340 70140 11396
rect 70140 11264 70196 11340
rect 69468 11172 69524 11182
rect 70028 11172 70084 11182
rect 69468 11170 70084 11172
rect 69468 11118 69470 11170
rect 69522 11118 70030 11170
rect 70082 11118 70084 11170
rect 69468 11116 70084 11118
rect 69468 11106 69524 11116
rect 69356 10994 69412 11004
rect 69356 10836 69412 10846
rect 69356 10742 69412 10780
rect 69468 10722 69524 10734
rect 69468 10670 69470 10722
rect 69522 10670 69524 10722
rect 69244 10388 69300 10398
rect 69244 10294 69300 10332
rect 68832 10220 69096 10230
rect 68888 10164 68936 10220
rect 68992 10164 69040 10220
rect 68832 10154 69096 10164
rect 69468 9938 69524 10670
rect 69468 9886 69470 9938
rect 69522 9886 69524 9938
rect 69468 9874 69524 9886
rect 69692 9828 69748 9838
rect 69692 9734 69748 9772
rect 69020 9716 69076 9726
rect 68908 9492 68964 9502
rect 68908 8820 68964 9436
rect 69020 9268 69076 9660
rect 70028 9716 70084 11116
rect 70140 11060 70196 11070
rect 70140 10722 70196 11004
rect 70476 10834 70532 12126
rect 71148 11506 71204 12684
rect 71372 12962 71428 12974
rect 71372 12910 71374 12962
rect 71426 12910 71428 12962
rect 71260 12292 71316 12302
rect 71372 12292 71428 12910
rect 71820 12962 71876 14700
rect 72044 14532 72100 14542
rect 72044 13970 72100 14476
rect 72044 13918 72046 13970
rect 72098 13918 72100 13970
rect 72044 13906 72100 13918
rect 72156 13970 72212 18172
rect 72492 16212 72548 19852
rect 73276 19906 73332 19918
rect 73276 19854 73278 19906
rect 73330 19854 73332 19906
rect 73276 19796 73332 19854
rect 73276 19730 73332 19740
rect 73836 19796 73892 20638
rect 73836 19348 73892 19740
rect 73836 19282 73892 19292
rect 73948 20580 74004 20590
rect 73724 18564 73780 18574
rect 73724 18338 73780 18508
rect 73724 18286 73726 18338
rect 73778 18286 73780 18338
rect 73724 18274 73780 18286
rect 73836 18562 73892 18574
rect 73836 18510 73838 18562
rect 73890 18510 73892 18562
rect 73836 18340 73892 18510
rect 73836 18274 73892 18284
rect 73948 18004 74004 20524
rect 74060 20018 74116 20030
rect 74060 19966 74062 20018
rect 74114 19966 74116 20018
rect 74060 19796 74116 19966
rect 74060 19730 74116 19740
rect 74172 20018 74228 20030
rect 74172 19966 74174 20018
rect 74226 19966 74228 20018
rect 74172 19684 74228 19966
rect 74284 19908 74340 20750
rect 74396 20244 74452 20254
rect 74508 20244 74564 26852
rect 74732 26628 74788 26910
rect 74732 26562 74788 26572
rect 74956 26850 75012 26862
rect 74956 26798 74958 26850
rect 75010 26798 75012 26850
rect 74956 25732 75012 26798
rect 74956 25666 75012 25676
rect 75068 26292 75124 26302
rect 74844 25172 74900 25182
rect 74844 23378 74900 25116
rect 74956 24948 75012 24958
rect 75068 24948 75124 26236
rect 75628 26292 75684 27022
rect 75628 26226 75684 26236
rect 75852 26962 75908 26974
rect 75852 26910 75854 26962
rect 75906 26910 75908 26962
rect 75516 26180 75572 26190
rect 75516 26086 75572 26124
rect 75852 25956 75908 26910
rect 75964 26964 76020 26974
rect 75964 26870 76020 26908
rect 76188 26290 76244 27132
rect 76188 26238 76190 26290
rect 76242 26238 76244 26290
rect 76188 26226 76244 26238
rect 75852 25890 75908 25900
rect 74956 24946 75124 24948
rect 74956 24894 74958 24946
rect 75010 24894 75124 24946
rect 74956 24892 75124 24894
rect 75852 25506 75908 25518
rect 75852 25454 75854 25506
rect 75906 25454 75908 25506
rect 75852 25172 75908 25454
rect 74956 24882 75012 24892
rect 75180 24834 75236 24846
rect 75180 24782 75182 24834
rect 75234 24782 75236 24834
rect 75180 24612 75236 24782
rect 75852 24836 75908 25116
rect 76300 24948 76356 28252
rect 76524 28196 76580 28206
rect 76524 28082 76580 28140
rect 76524 28030 76526 28082
rect 76578 28030 76580 28082
rect 76524 28018 76580 28030
rect 76412 27860 76468 27870
rect 76636 27860 76692 29150
rect 76972 28980 77028 29260
rect 77084 29250 77140 29260
rect 76748 27972 76804 27982
rect 76748 27878 76804 27916
rect 76412 27858 76692 27860
rect 76412 27806 76414 27858
rect 76466 27806 76692 27858
rect 76412 27804 76692 27806
rect 76972 27860 77028 28924
rect 76412 27524 76468 27804
rect 76412 27458 76468 27468
rect 76412 27300 76468 27310
rect 76412 27206 76468 27244
rect 76972 27076 77028 27804
rect 76972 27010 77028 27020
rect 76524 25620 76580 25630
rect 76524 25526 76580 25564
rect 75852 24770 75908 24780
rect 75964 24892 76356 24948
rect 76412 25506 76468 25518
rect 76412 25454 76414 25506
rect 76466 25454 76468 25506
rect 76412 24948 76468 25454
rect 76412 24892 76916 24948
rect 75292 24724 75348 24734
rect 75292 24630 75348 24668
rect 75180 24546 75236 24556
rect 75516 24050 75572 24062
rect 75516 23998 75518 24050
rect 75570 23998 75572 24050
rect 75516 23716 75572 23998
rect 75516 23650 75572 23660
rect 74844 23326 74846 23378
rect 74898 23326 74900 23378
rect 74844 23314 74900 23326
rect 75628 23492 75684 23502
rect 74732 23042 74788 23054
rect 74732 22990 74734 23042
rect 74786 22990 74788 23042
rect 74620 22370 74676 22382
rect 74620 22318 74622 22370
rect 74674 22318 74676 22370
rect 74620 21700 74676 22318
rect 74732 22148 74788 22990
rect 75628 23042 75684 23436
rect 75628 22990 75630 23042
rect 75682 22990 75684 23042
rect 75628 22978 75684 22990
rect 75740 23154 75796 23166
rect 75740 23102 75742 23154
rect 75794 23102 75796 23154
rect 75740 23044 75796 23102
rect 75740 22978 75796 22988
rect 75628 22372 75684 22382
rect 75628 22278 75684 22316
rect 75852 22370 75908 22382
rect 75852 22318 75854 22370
rect 75906 22318 75908 22370
rect 74732 22082 74788 22092
rect 74844 22258 74900 22270
rect 74844 22206 74846 22258
rect 74898 22206 74900 22258
rect 74620 21634 74676 21644
rect 74844 20916 74900 22206
rect 75404 22260 75460 22270
rect 75404 22166 75460 22204
rect 75852 21812 75908 22318
rect 75852 21746 75908 21756
rect 74956 21588 75012 21598
rect 74956 21494 75012 21532
rect 74844 20850 74900 20860
rect 75068 21028 75124 21038
rect 74396 20242 74564 20244
rect 74396 20190 74398 20242
rect 74450 20190 74564 20242
rect 74396 20188 74564 20190
rect 74732 20690 74788 20702
rect 74732 20638 74734 20690
rect 74786 20638 74788 20690
rect 74396 20178 74452 20188
rect 74620 20132 74676 20142
rect 74284 19842 74340 19852
rect 74396 20020 74452 20030
rect 74620 20020 74676 20076
rect 74172 19618 74228 19628
rect 74396 19348 74452 19964
rect 74396 19216 74452 19292
rect 74508 20018 74676 20020
rect 74508 19966 74622 20018
rect 74674 19966 74676 20018
rect 74508 19964 74676 19966
rect 74060 18228 74116 18238
rect 74060 18134 74116 18172
rect 73948 17948 74116 18004
rect 73948 17556 74004 17566
rect 73500 17444 73556 17454
rect 73948 17444 74004 17500
rect 73500 17442 74004 17444
rect 73500 17390 73502 17442
rect 73554 17390 74004 17442
rect 73500 17388 74004 17390
rect 73500 17378 73556 17388
rect 72492 16210 73220 16212
rect 72492 16158 72494 16210
rect 72546 16158 73220 16210
rect 72492 16156 73220 16158
rect 72492 16146 72548 16156
rect 72380 16100 72436 16110
rect 72268 16098 72436 16100
rect 72268 16046 72382 16098
rect 72434 16046 72436 16098
rect 72268 16044 72436 16046
rect 72268 15428 72324 16044
rect 72380 16034 72436 16044
rect 73164 15428 73220 16156
rect 73276 16100 73332 16110
rect 73276 16006 73332 16044
rect 73388 15428 73444 15438
rect 73164 15426 73444 15428
rect 73164 15374 73390 15426
rect 73442 15374 73444 15426
rect 73164 15372 73444 15374
rect 72268 14084 72324 15372
rect 73388 15362 73444 15372
rect 73500 15428 73556 15438
rect 73500 15334 73556 15372
rect 73612 15316 73668 17388
rect 74060 17106 74116 17948
rect 74508 17890 74564 19964
rect 74620 19954 74676 19964
rect 74732 19908 74788 20638
rect 74732 19842 74788 19852
rect 74620 18452 74676 18462
rect 74620 18358 74676 18396
rect 74508 17838 74510 17890
rect 74562 17838 74564 17890
rect 74508 17826 74564 17838
rect 74620 17668 74676 17678
rect 74620 17574 74676 17612
rect 74508 17556 74564 17566
rect 74508 17462 74564 17500
rect 74060 17054 74062 17106
rect 74114 17054 74116 17106
rect 74060 17042 74116 17054
rect 73724 16994 73780 17006
rect 73724 16942 73726 16994
rect 73778 16942 73780 16994
rect 73724 15538 73780 16942
rect 73948 16882 74004 16894
rect 73948 16830 73950 16882
rect 74002 16830 74004 16882
rect 73948 16100 74004 16830
rect 74172 16884 74228 16894
rect 74172 16882 74340 16884
rect 74172 16830 74174 16882
rect 74226 16830 74340 16882
rect 74172 16828 74340 16830
rect 74172 16818 74228 16828
rect 74284 16212 74340 16828
rect 74396 16212 74452 16222
rect 74284 16210 74452 16212
rect 74284 16158 74398 16210
rect 74450 16158 74452 16210
rect 74284 16156 74452 16158
rect 74172 16100 74228 16110
rect 74004 16098 74228 16100
rect 74004 16046 74174 16098
rect 74226 16046 74228 16098
rect 74004 16044 74228 16046
rect 73948 15968 74004 16044
rect 74172 16034 74228 16044
rect 73724 15486 73726 15538
rect 73778 15486 73780 15538
rect 73724 15474 73780 15486
rect 74060 15428 74116 15438
rect 74060 15334 74116 15372
rect 73612 15260 73780 15316
rect 72492 15204 72548 15214
rect 72380 15202 72548 15204
rect 72380 15150 72494 15202
rect 72546 15150 72548 15202
rect 72380 15148 72548 15150
rect 72380 14644 72436 15148
rect 72492 15138 72548 15148
rect 72604 15092 72660 15102
rect 72604 15090 73668 15092
rect 72604 15038 72606 15090
rect 72658 15038 73668 15090
rect 72604 15036 73668 15038
rect 72604 15026 72660 15036
rect 72380 14550 72436 14588
rect 73052 14644 73108 14654
rect 73052 14550 73108 14588
rect 73500 14530 73556 14542
rect 73500 14478 73502 14530
rect 73554 14478 73556 14530
rect 72268 14028 72660 14084
rect 72156 13918 72158 13970
rect 72210 13918 72212 13970
rect 72156 13906 72212 13918
rect 72268 13748 72324 13758
rect 72268 13654 72324 13692
rect 71820 12910 71822 12962
rect 71874 12910 71876 12962
rect 71820 12898 71876 12910
rect 72380 12852 72436 12862
rect 71260 12290 71428 12292
rect 71260 12238 71262 12290
rect 71314 12238 71428 12290
rect 71260 12236 71428 12238
rect 71260 12226 71316 12236
rect 71148 11454 71150 11506
rect 71202 11454 71204 11506
rect 71148 11442 71204 11454
rect 71260 11618 71316 11630
rect 71260 11566 71262 11618
rect 71314 11566 71316 11618
rect 70476 10782 70478 10834
rect 70530 10782 70532 10834
rect 70476 10770 70532 10782
rect 70812 11396 70868 11406
rect 70812 10834 70868 11340
rect 70812 10782 70814 10834
rect 70866 10782 70868 10834
rect 70812 10770 70868 10782
rect 71036 11060 71092 11070
rect 70140 10670 70142 10722
rect 70194 10670 70196 10722
rect 70140 10658 70196 10670
rect 70252 10724 70308 10734
rect 70252 10722 70420 10724
rect 70252 10670 70254 10722
rect 70306 10670 70420 10722
rect 70252 10668 70420 10670
rect 70252 10658 70308 10668
rect 70028 9650 70084 9660
rect 70252 9714 70308 9726
rect 70252 9662 70254 9714
rect 70306 9662 70308 9714
rect 69468 9602 69524 9614
rect 69468 9550 69470 9602
rect 69522 9550 69524 9602
rect 69468 9492 69524 9550
rect 69468 9426 69524 9436
rect 70028 9492 70084 9502
rect 69580 9268 69636 9278
rect 69020 9266 69300 9268
rect 69020 9214 69022 9266
rect 69074 9214 69300 9266
rect 69020 9212 69300 9214
rect 69020 9156 69076 9212
rect 69020 9090 69076 9100
rect 69132 9044 69188 9054
rect 69132 8950 69188 8988
rect 69020 8820 69076 8830
rect 68908 8818 69076 8820
rect 68908 8766 69022 8818
rect 69074 8766 69076 8818
rect 68908 8764 69076 8766
rect 69020 8754 69076 8764
rect 68832 8652 69096 8662
rect 68888 8596 68936 8652
rect 68992 8596 69040 8652
rect 68832 8586 69096 8596
rect 68460 8372 68740 8428
rect 68460 8260 68516 8372
rect 69244 8370 69300 9212
rect 69244 8318 69246 8370
rect 69298 8318 69300 8370
rect 69244 8306 69300 8318
rect 69468 9212 69580 9268
rect 68012 7982 68014 8034
rect 68066 7982 68068 8034
rect 68012 7250 68068 7982
rect 68236 8204 68516 8260
rect 68124 7588 68180 7598
rect 68124 7494 68180 7532
rect 68012 7198 68014 7250
rect 68066 7198 68068 7250
rect 68012 7186 68068 7198
rect 67788 6638 67790 6690
rect 67842 6638 67844 6690
rect 67788 6626 67844 6638
rect 68012 6690 68068 6702
rect 68012 6638 68014 6690
rect 68066 6638 68068 6690
rect 67676 6414 67678 6466
rect 67730 6414 67732 6466
rect 67676 6356 67732 6414
rect 67900 6468 67956 6478
rect 67900 6374 67956 6412
rect 67676 6290 67732 6300
rect 67116 5954 67172 5964
rect 67228 6132 67284 6142
rect 67228 5684 67284 6076
rect 67564 6132 67620 6142
rect 68012 6132 68068 6638
rect 67564 6130 68068 6132
rect 67564 6078 67566 6130
rect 67618 6078 68068 6130
rect 67564 6076 68068 6078
rect 67564 6066 67620 6076
rect 67452 6020 67508 6030
rect 67452 5908 67508 5964
rect 67900 5908 67956 5918
rect 67452 5906 67956 5908
rect 67452 5854 67902 5906
rect 67954 5854 67956 5906
rect 67452 5852 67956 5854
rect 67900 5842 67956 5852
rect 68124 5908 68180 5918
rect 68124 5814 68180 5852
rect 67228 5618 67284 5628
rect 67004 5282 67060 5292
rect 66668 5170 66724 5180
rect 66556 5124 66612 5134
rect 66556 5030 66612 5068
rect 67676 5122 67732 5134
rect 67900 5124 67956 5134
rect 67676 5070 67678 5122
rect 67730 5070 67732 5122
rect 67676 5012 67732 5070
rect 67676 4946 67732 4956
rect 67788 5122 67956 5124
rect 67788 5070 67902 5122
rect 67954 5070 67956 5122
rect 67788 5068 67956 5070
rect 66332 4806 66388 4844
rect 66556 4900 66612 4910
rect 66220 4722 66276 4732
rect 66556 3554 66612 4844
rect 66892 4898 66948 4910
rect 66892 4846 66894 4898
rect 66946 4846 66948 4898
rect 66892 4564 66948 4846
rect 66892 4498 66948 4508
rect 67004 4788 67060 4798
rect 66556 3502 66558 3554
rect 66610 3502 66612 3554
rect 66220 3444 66276 3454
rect 66108 3442 66276 3444
rect 66108 3390 66222 3442
rect 66274 3390 66276 3442
rect 66108 3388 66276 3390
rect 65660 3350 65716 3388
rect 66220 3378 66276 3388
rect 65436 1362 65492 1372
rect 66556 800 66612 3502
rect 67004 4338 67060 4732
rect 67004 4286 67006 4338
rect 67058 4286 67060 4338
rect 67004 2996 67060 4286
rect 67116 4676 67172 4686
rect 67116 3666 67172 4620
rect 67340 4340 67396 4350
rect 67340 3892 67396 4284
rect 67676 4116 67732 4126
rect 67676 4022 67732 4060
rect 67340 3778 67396 3836
rect 67340 3726 67342 3778
rect 67394 3726 67396 3778
rect 67340 3714 67396 3726
rect 67676 3780 67732 3790
rect 67788 3780 67844 5068
rect 67900 5058 67956 5068
rect 68236 5010 68292 8204
rect 68460 8034 68516 8046
rect 68460 7982 68462 8034
rect 68514 7982 68516 8034
rect 68460 7924 68516 7982
rect 68460 7858 68516 7868
rect 68460 7700 68516 7710
rect 68460 7606 68516 7644
rect 69356 7476 69412 7486
rect 69356 7382 69412 7420
rect 68460 7250 68516 7262
rect 68460 7198 68462 7250
rect 68514 7198 68516 7250
rect 68348 6692 68404 6702
rect 68348 6598 68404 6636
rect 68236 4958 68238 5010
rect 68290 4958 68292 5010
rect 68236 4946 68292 4958
rect 68124 4898 68180 4910
rect 68124 4846 68126 4898
rect 68178 4846 68180 4898
rect 68124 4788 68180 4846
rect 68124 4564 68180 4732
rect 68124 4498 68180 4508
rect 68348 4898 68404 4910
rect 68348 4846 68350 4898
rect 68402 4846 68404 4898
rect 68348 4788 68404 4846
rect 68236 4452 68292 4462
rect 68236 4358 68292 4396
rect 68348 4228 68404 4732
rect 68348 4162 68404 4172
rect 67676 3778 67844 3780
rect 67676 3726 67678 3778
rect 67730 3726 67844 3778
rect 67676 3724 67844 3726
rect 67676 3714 67732 3724
rect 67116 3614 67118 3666
rect 67170 3614 67172 3666
rect 67116 3602 67172 3614
rect 68460 3668 68516 7198
rect 68832 7084 69096 7094
rect 68888 7028 68936 7084
rect 68992 7028 69040 7084
rect 68832 7018 69096 7028
rect 68572 6692 68628 6702
rect 68572 6130 68628 6636
rect 68572 6078 68574 6130
rect 68626 6078 68628 6130
rect 68572 6066 68628 6078
rect 68908 6468 68964 6478
rect 68796 6018 68852 6030
rect 68796 5966 68798 6018
rect 68850 5966 68852 6018
rect 68796 5684 68852 5966
rect 68908 6018 68964 6412
rect 69468 6468 69524 9212
rect 69580 9174 69636 9212
rect 70028 9266 70084 9436
rect 70028 9214 70030 9266
rect 70082 9214 70084 9266
rect 70028 9202 70084 9214
rect 70252 9268 70308 9662
rect 70364 9604 70420 10668
rect 70588 9828 70644 9838
rect 71036 9828 71092 11004
rect 70588 9734 70644 9772
rect 70924 9826 71092 9828
rect 70924 9774 71038 9826
rect 71090 9774 71092 9826
rect 70924 9772 71092 9774
rect 70364 9602 70532 9604
rect 70364 9550 70366 9602
rect 70418 9550 70532 9602
rect 70364 9548 70532 9550
rect 70364 9538 70420 9548
rect 70252 9202 70308 9212
rect 70364 9044 70420 9054
rect 69804 8932 69860 8942
rect 69692 8260 69748 8270
rect 69692 7812 69748 8204
rect 69804 8148 69860 8876
rect 70364 8372 70420 8988
rect 70476 8932 70532 9548
rect 70476 8838 70532 8876
rect 70924 9266 70980 9772
rect 71036 9762 71092 9772
rect 71148 9716 71204 9726
rect 71148 9622 71204 9660
rect 70924 9214 70926 9266
rect 70978 9214 70980 9266
rect 70924 8932 70980 9214
rect 70924 8866 70980 8876
rect 71260 8428 71316 11566
rect 71372 11394 71428 12236
rect 71372 11342 71374 11394
rect 71426 11342 71428 11394
rect 71372 11330 71428 11342
rect 71596 12738 71652 12750
rect 71596 12686 71598 12738
rect 71650 12686 71652 12738
rect 71596 10836 71652 12686
rect 72380 12738 72436 12796
rect 72380 12686 72382 12738
rect 72434 12686 72436 12738
rect 72380 11956 72436 12686
rect 72380 11890 72436 11900
rect 72268 11170 72324 11182
rect 72268 11118 72270 11170
rect 72322 11118 72324 11170
rect 72268 11060 72324 11118
rect 72268 10994 72324 11004
rect 71372 10780 71876 10836
rect 71372 9826 71428 10780
rect 71820 10500 71876 10780
rect 72156 10610 72212 10622
rect 72156 10558 72158 10610
rect 72210 10558 72212 10610
rect 71820 10498 72100 10500
rect 71820 10446 71822 10498
rect 71874 10446 72100 10498
rect 71820 10444 72100 10446
rect 71820 10434 71876 10444
rect 72044 10050 72100 10444
rect 72044 9998 72046 10050
rect 72098 9998 72100 10050
rect 72044 9986 72100 9998
rect 71372 9774 71374 9826
rect 71426 9774 71428 9826
rect 71372 9762 71428 9774
rect 72156 9828 72212 10558
rect 72492 10500 72548 10510
rect 72492 10406 72548 10444
rect 72156 9716 72212 9772
rect 72380 9938 72436 9950
rect 72380 9886 72382 9938
rect 72434 9886 72436 9938
rect 72268 9716 72324 9726
rect 72156 9714 72324 9716
rect 72156 9662 72270 9714
rect 72322 9662 72324 9714
rect 72156 9660 72324 9662
rect 72380 9716 72436 9886
rect 72492 9716 72548 9726
rect 72380 9714 72548 9716
rect 72380 9662 72494 9714
rect 72546 9662 72548 9714
rect 72380 9660 72548 9662
rect 72268 9650 72324 9660
rect 72492 9650 72548 9660
rect 71708 9268 71764 9278
rect 70476 8372 70532 8382
rect 70364 8370 70532 8372
rect 70364 8318 70478 8370
rect 70530 8318 70532 8370
rect 70364 8316 70532 8318
rect 70476 8306 70532 8316
rect 71148 8372 71316 8428
rect 71372 9266 71764 9268
rect 71372 9214 71710 9266
rect 71762 9214 71764 9266
rect 71372 9212 71764 9214
rect 71148 8258 71204 8372
rect 71148 8206 71150 8258
rect 71202 8206 71204 8258
rect 69804 8054 69860 8092
rect 70364 8148 70420 8158
rect 70364 8054 70420 8092
rect 71148 8148 71204 8206
rect 71148 8082 71204 8092
rect 71372 8258 71428 9212
rect 71708 9202 71764 9212
rect 72268 9268 72324 9278
rect 72268 9174 72324 9212
rect 71596 9044 71652 9054
rect 71596 8950 71652 8988
rect 71932 9044 71988 9054
rect 71932 8950 71988 8988
rect 71372 8206 71374 8258
rect 71426 8206 71428 8258
rect 69692 7700 69748 7756
rect 69804 7700 69860 7710
rect 69692 7698 69860 7700
rect 69692 7646 69806 7698
rect 69858 7646 69860 7698
rect 69692 7644 69860 7646
rect 69804 7634 69860 7644
rect 69916 7700 69972 7710
rect 69916 7606 69972 7644
rect 71372 7700 71428 8206
rect 72044 8260 72100 8270
rect 72044 8166 72100 8204
rect 71372 7634 71428 7644
rect 70588 7588 70644 7598
rect 70588 7494 70644 7532
rect 70028 7476 70084 7486
rect 69916 7474 70084 7476
rect 69916 7422 70030 7474
rect 70082 7422 70084 7474
rect 69916 7420 70084 7422
rect 69580 7364 69636 7374
rect 69580 6916 69636 7308
rect 69580 6850 69636 6860
rect 69468 6402 69524 6412
rect 69692 6580 69748 6590
rect 69916 6580 69972 7420
rect 70028 7410 70084 7420
rect 71708 7476 71764 7486
rect 71708 7382 71764 7420
rect 71820 7364 71876 7374
rect 71820 7270 71876 7308
rect 72268 7250 72324 7262
rect 72268 7198 72270 7250
rect 72322 7198 72324 7250
rect 70028 6692 70084 6702
rect 70028 6598 70084 6636
rect 70924 6692 70980 6702
rect 69692 6578 69972 6580
rect 69692 6526 69694 6578
rect 69746 6526 69972 6578
rect 69692 6524 69972 6526
rect 70252 6580 70308 6590
rect 68908 5966 68910 6018
rect 68962 5966 68964 6018
rect 68908 5954 68964 5966
rect 69692 5908 69748 6524
rect 69804 6132 69860 6142
rect 69804 6038 69860 6076
rect 70252 6130 70308 6524
rect 70700 6356 70756 6366
rect 70252 6078 70254 6130
rect 70306 6078 70308 6130
rect 70252 6066 70308 6078
rect 70588 6132 70644 6142
rect 69692 5842 69748 5852
rect 68796 5618 68852 5628
rect 69356 5796 69412 5806
rect 68832 5516 69096 5526
rect 68888 5460 68936 5516
rect 68992 5460 69040 5516
rect 68832 5450 69096 5460
rect 69244 5236 69300 5246
rect 69356 5236 69412 5740
rect 69244 5234 69412 5236
rect 69244 5182 69246 5234
rect 69298 5182 69412 5234
rect 69244 5180 69412 5182
rect 69692 5236 69748 5246
rect 69244 5170 69300 5180
rect 69692 5142 69748 5180
rect 70588 5234 70644 6076
rect 70700 6130 70756 6300
rect 70700 6078 70702 6130
rect 70754 6078 70756 6130
rect 70700 6066 70756 6078
rect 70924 6020 70980 6636
rect 72156 6690 72212 6702
rect 72156 6638 72158 6690
rect 72210 6638 72212 6690
rect 70924 5954 70980 5964
rect 71036 6468 71092 6478
rect 70588 5182 70590 5234
rect 70642 5182 70644 5234
rect 70588 5170 70644 5182
rect 70252 5122 70308 5134
rect 70252 5070 70254 5122
rect 70306 5070 70308 5122
rect 69132 5012 69188 5022
rect 69132 4226 69188 4956
rect 69580 4676 69636 4686
rect 69580 4452 69636 4620
rect 70252 4564 70308 5070
rect 70252 4498 70308 4508
rect 69580 4338 69636 4396
rect 69580 4286 69582 4338
rect 69634 4286 69636 4338
rect 69580 4274 69636 4286
rect 70924 4340 70980 4350
rect 70924 4246 70980 4284
rect 69132 4174 69134 4226
rect 69186 4174 69188 4226
rect 69132 4162 69188 4174
rect 68832 3948 69096 3958
rect 68888 3892 68936 3948
rect 68992 3892 69040 3948
rect 68832 3882 69096 3892
rect 68908 3668 68964 3678
rect 68460 3666 68964 3668
rect 68460 3614 68910 3666
rect 68962 3614 68964 3666
rect 68460 3612 68964 3614
rect 68908 3602 68964 3612
rect 70252 3668 70308 3678
rect 68348 3556 68404 3566
rect 68348 3462 68404 3500
rect 67004 2930 67060 2940
rect 68684 3444 68740 3454
rect 68684 800 68740 3388
rect 70252 3444 70308 3612
rect 70252 3312 70308 3388
rect 70812 3444 70868 3454
rect 70812 800 70868 3388
rect 71036 3330 71092 6412
rect 71484 6468 71540 6478
rect 71484 6374 71540 6412
rect 72044 5908 72100 5918
rect 72044 5814 72100 5852
rect 72044 5572 72100 5582
rect 71708 5236 71764 5246
rect 71372 5234 71988 5236
rect 71372 5182 71710 5234
rect 71762 5182 71988 5234
rect 71372 5180 71988 5182
rect 71372 4450 71428 5180
rect 71708 5170 71764 5180
rect 71372 4398 71374 4450
rect 71426 4398 71428 4450
rect 71932 4506 71988 5180
rect 71932 4454 71934 4506
rect 71986 4454 71988 4506
rect 71932 4442 71988 4454
rect 72044 5122 72100 5516
rect 72044 5070 72046 5122
rect 72098 5070 72100 5122
rect 72044 4450 72100 5070
rect 71372 4386 71428 4398
rect 72044 4398 72046 4450
rect 72098 4398 72100 4450
rect 72044 4340 72100 4398
rect 71932 4284 72100 4340
rect 71372 3444 71428 3454
rect 71372 3350 71428 3388
rect 71036 3278 71038 3330
rect 71090 3278 71092 3330
rect 71036 3266 71092 3278
rect 71932 3332 71988 4284
rect 72044 4116 72100 4126
rect 72156 4116 72212 6638
rect 72268 6580 72324 7198
rect 72604 6690 72660 14028
rect 73500 13860 73556 14478
rect 73500 13766 73556 13804
rect 73612 13858 73668 15036
rect 73612 13806 73614 13858
rect 73666 13806 73668 13858
rect 73612 13794 73668 13806
rect 72716 13748 72772 13758
rect 73276 13748 73332 13758
rect 72716 13746 73332 13748
rect 72716 13694 72718 13746
rect 72770 13694 73278 13746
rect 73330 13694 73332 13746
rect 72716 13692 73332 13694
rect 72716 13682 72772 13692
rect 73276 13682 73332 13692
rect 73724 13636 73780 15260
rect 74396 15148 74452 16156
rect 74844 16100 74900 16110
rect 74844 16006 74900 16044
rect 74508 15428 74564 15438
rect 74508 15334 74564 15372
rect 73948 15092 74452 15148
rect 73948 14642 74004 15092
rect 73948 14590 73950 14642
rect 74002 14590 74004 14642
rect 73948 14578 74004 14590
rect 74508 14644 74564 14654
rect 75068 14644 75124 20972
rect 75516 20916 75572 20926
rect 75516 20822 75572 20860
rect 75180 20802 75236 20814
rect 75180 20750 75182 20802
rect 75234 20750 75236 20802
rect 75180 20580 75236 20750
rect 75180 20514 75236 20524
rect 75292 20020 75348 20030
rect 75292 19926 75348 19964
rect 75404 19908 75460 19918
rect 75404 19814 75460 19852
rect 75628 19796 75684 19806
rect 75628 19702 75684 19740
rect 75516 19346 75572 19358
rect 75516 19294 75518 19346
rect 75570 19294 75572 19346
rect 75516 19012 75572 19294
rect 75516 18946 75572 18956
rect 75180 18450 75236 18462
rect 75180 18398 75182 18450
rect 75234 18398 75236 18450
rect 75180 18228 75236 18398
rect 75180 17780 75236 18172
rect 75180 17686 75236 17724
rect 75628 17666 75684 17678
rect 75628 17614 75630 17666
rect 75682 17614 75684 17666
rect 75628 17556 75684 17614
rect 75628 17490 75684 17500
rect 75180 17444 75236 17454
rect 75180 16882 75236 17388
rect 75180 16830 75182 16882
rect 75234 16830 75236 16882
rect 75180 16818 75236 16830
rect 75516 17444 75572 17454
rect 75292 16548 75348 16558
rect 74508 14642 75124 14644
rect 74508 14590 74510 14642
rect 74562 14590 75124 14642
rect 74508 14588 75124 14590
rect 74508 14578 74564 14588
rect 75068 14530 75124 14588
rect 75068 14478 75070 14530
rect 75122 14478 75124 14530
rect 75068 14466 75124 14478
rect 75180 15316 75236 15326
rect 73612 13580 73780 13636
rect 74620 14420 74676 14430
rect 73500 12404 73556 12414
rect 73500 12310 73556 12348
rect 73388 12178 73444 12190
rect 73388 12126 73390 12178
rect 73442 12126 73444 12178
rect 73388 11396 73444 12126
rect 73388 11330 73444 11340
rect 73388 10500 73444 10510
rect 73388 10406 73444 10444
rect 73500 10498 73556 10510
rect 73500 10446 73502 10498
rect 73554 10446 73556 10498
rect 73276 10052 73332 10062
rect 73500 10052 73556 10446
rect 73276 10050 73556 10052
rect 73276 9998 73278 10050
rect 73330 9998 73556 10050
rect 73276 9996 73556 9998
rect 73276 9986 73332 9996
rect 73612 9940 73668 13580
rect 74060 12404 74116 12414
rect 74060 12310 74116 12348
rect 73724 12178 73780 12190
rect 73724 12126 73726 12178
rect 73778 12126 73780 12178
rect 73724 10612 73780 12126
rect 73836 11396 73892 11406
rect 73892 11340 74116 11396
rect 73836 11302 73892 11340
rect 73724 10518 73780 10556
rect 73500 9884 73668 9940
rect 72940 9826 72996 9838
rect 72940 9774 72942 9826
rect 72994 9774 72996 9826
rect 72828 9716 72884 9726
rect 72940 9716 72996 9774
rect 72828 9714 72996 9716
rect 72828 9662 72830 9714
rect 72882 9662 72996 9714
rect 72828 9660 72996 9662
rect 73164 9716 73220 9726
rect 73388 9716 73444 9726
rect 73164 9714 73444 9716
rect 73164 9662 73166 9714
rect 73218 9662 73390 9714
rect 73442 9662 73444 9714
rect 73164 9660 73444 9662
rect 72828 9650 72884 9660
rect 73052 8932 73108 8942
rect 72716 8260 72772 8270
rect 72716 8166 72772 8204
rect 72604 6638 72606 6690
rect 72658 6638 72660 6690
rect 72604 6626 72660 6638
rect 72268 6514 72324 6524
rect 72380 6468 72436 6478
rect 72380 5906 72436 6412
rect 72380 5854 72382 5906
rect 72434 5854 72436 5906
rect 72380 5842 72436 5854
rect 72492 6466 72548 6478
rect 72492 6414 72494 6466
rect 72546 6414 72548 6466
rect 72492 5908 72548 6414
rect 72716 6468 72772 6478
rect 72716 6374 72772 6412
rect 73052 5908 73108 8876
rect 73164 8258 73220 9660
rect 73388 9650 73444 9660
rect 73500 9266 73556 9884
rect 73500 9214 73502 9266
rect 73554 9214 73556 9266
rect 73500 9202 73556 9214
rect 73612 9714 73668 9726
rect 73612 9662 73614 9714
rect 73666 9662 73668 9714
rect 73612 9266 73668 9662
rect 73724 9716 73780 9726
rect 73724 9622 73780 9660
rect 73612 9214 73614 9266
rect 73666 9214 73668 9266
rect 73612 9202 73668 9214
rect 73164 8206 73166 8258
rect 73218 8206 73220 8258
rect 73164 8194 73220 8206
rect 73388 9154 73444 9166
rect 73388 9102 73390 9154
rect 73442 9102 73444 9154
rect 73388 8260 73444 9102
rect 73948 9044 74004 9054
rect 73948 8950 74004 8988
rect 74060 8428 74116 11340
rect 74508 11170 74564 11182
rect 74508 11118 74510 11170
rect 74562 11118 74564 11170
rect 74508 10388 74564 11118
rect 74508 10322 74564 10332
rect 74620 9940 74676 14364
rect 75180 14084 75236 15260
rect 74844 14028 75236 14084
rect 74844 11506 74900 14028
rect 75292 13972 75348 16492
rect 75404 16212 75460 16222
rect 75404 15540 75460 16156
rect 75516 16210 75572 17388
rect 75964 16548 76020 24892
rect 76860 24836 76916 24892
rect 76300 24722 76356 24734
rect 76300 24670 76302 24722
rect 76354 24670 76356 24722
rect 76300 24612 76356 24670
rect 76300 24546 76356 24556
rect 76412 24724 76468 24734
rect 76860 24704 76916 24780
rect 76412 24610 76468 24668
rect 76412 24558 76414 24610
rect 76466 24558 76468 24610
rect 76188 23940 76244 23950
rect 76188 23846 76244 23884
rect 76412 23266 76468 24558
rect 76412 23214 76414 23266
rect 76466 23214 76468 23266
rect 76412 23202 76468 23214
rect 76860 23044 76916 23054
rect 76860 22950 76916 22988
rect 76748 22372 76804 22382
rect 76748 21698 76804 22316
rect 77084 22148 77140 22158
rect 76860 21812 76916 21822
rect 76860 21718 76916 21756
rect 77084 21810 77140 22092
rect 77084 21758 77086 21810
rect 77138 21758 77140 21810
rect 77084 21746 77140 21758
rect 76748 21646 76750 21698
rect 76802 21646 76804 21698
rect 76748 21634 76804 21646
rect 76076 21474 76132 21486
rect 76076 21422 76078 21474
rect 76130 21422 76132 21474
rect 76076 21252 76132 21422
rect 76076 21186 76132 21196
rect 76972 20132 77028 20142
rect 76972 20038 77028 20076
rect 76748 20020 76804 20030
rect 76636 20018 76804 20020
rect 76636 19966 76750 20018
rect 76802 19966 76804 20018
rect 76636 19964 76804 19966
rect 76636 19684 76692 19964
rect 76748 19954 76804 19964
rect 77084 20018 77140 20030
rect 77084 19966 77086 20018
rect 77138 19966 77140 20018
rect 77084 19796 77140 19966
rect 77084 19730 77140 19740
rect 76188 19236 76244 19246
rect 76188 19142 76244 19180
rect 76636 18564 76692 19628
rect 77196 19348 77252 32622
rect 77420 31948 77476 33068
rect 77532 32900 77588 33294
rect 77756 33012 77812 34188
rect 77532 32834 77588 32844
rect 77644 32956 77812 33012
rect 77532 32676 77588 32686
rect 77532 32582 77588 32620
rect 77308 31892 77364 31902
rect 77420 31892 77588 31948
rect 77308 31798 77364 31836
rect 77532 31780 77588 31892
rect 77532 31714 77588 31724
rect 77420 31668 77476 31678
rect 77420 31574 77476 31612
rect 77532 31556 77588 31566
rect 77532 31462 77588 31500
rect 77644 31220 77700 32956
rect 77868 31948 77924 34636
rect 77980 34356 78036 35084
rect 78092 35028 78148 39200
rect 78492 36092 78756 36102
rect 78548 36036 78596 36092
rect 78652 36036 78700 36092
rect 78492 36026 78756 36036
rect 78092 34962 78148 34972
rect 78092 34804 78148 34814
rect 78092 34710 78148 34748
rect 78492 34524 78756 34534
rect 78548 34468 78596 34524
rect 78652 34468 78700 34524
rect 78492 34458 78756 34468
rect 77980 34300 78148 34356
rect 77980 34132 78036 34142
rect 77980 34038 78036 34076
rect 78092 33348 78148 34300
rect 78876 34244 78932 34254
rect 77980 33292 78148 33348
rect 78204 34132 78260 34142
rect 77980 32676 78036 33292
rect 78092 33122 78148 33134
rect 78092 33070 78094 33122
rect 78146 33070 78148 33122
rect 78092 32900 78148 33070
rect 78092 32834 78148 32844
rect 77980 32544 78036 32620
rect 78204 31948 78260 34076
rect 78492 32956 78756 32966
rect 78548 32900 78596 32956
rect 78652 32900 78700 32956
rect 78492 32890 78756 32900
rect 77420 31164 77700 31220
rect 77756 31892 77924 31948
rect 78092 31892 78260 31948
rect 77308 30772 77364 30782
rect 77308 30210 77364 30716
rect 77308 30158 77310 30210
rect 77362 30158 77364 30210
rect 77308 30146 77364 30158
rect 77308 28868 77364 28878
rect 77308 28774 77364 28812
rect 77308 27972 77364 27982
rect 77308 27298 77364 27916
rect 77308 27246 77310 27298
rect 77362 27246 77364 27298
rect 77308 27234 77364 27246
rect 77308 27076 77364 27114
rect 77420 27076 77476 31164
rect 77644 30996 77700 31006
rect 77644 30902 77700 30940
rect 77756 30324 77812 31892
rect 78092 31890 78148 31892
rect 78092 31838 78094 31890
rect 78146 31838 78148 31890
rect 78092 31826 78148 31838
rect 77644 30268 77812 30324
rect 78204 31780 78260 31790
rect 77532 30098 77588 30110
rect 77532 30046 77534 30098
rect 77586 30046 77588 30098
rect 77532 29876 77588 30046
rect 77532 29810 77588 29820
rect 77644 29540 77700 30268
rect 77868 30212 77924 30222
rect 77756 30100 77812 30110
rect 77756 30006 77812 30044
rect 77868 30098 77924 30156
rect 77868 30046 77870 30098
rect 77922 30046 77924 30098
rect 77644 29484 77812 29540
rect 77644 29314 77700 29326
rect 77644 29262 77646 29314
rect 77698 29262 77700 29314
rect 77644 29202 77700 29262
rect 77644 29150 77646 29202
rect 77698 29150 77700 29202
rect 77644 29138 77700 29150
rect 77644 28756 77700 28766
rect 77644 28642 77700 28700
rect 77644 28590 77646 28642
rect 77698 28590 77700 28642
rect 77644 27748 77700 28590
rect 77756 28196 77812 29484
rect 77868 29092 77924 30046
rect 77980 29316 78036 29326
rect 77980 29314 78148 29316
rect 77980 29262 77982 29314
rect 78034 29262 78148 29314
rect 77980 29260 78148 29262
rect 77980 29250 78036 29260
rect 77868 29036 78036 29092
rect 77868 28868 77924 28878
rect 77868 28754 77924 28812
rect 77868 28702 77870 28754
rect 77922 28702 77924 28754
rect 77868 28690 77924 28702
rect 77980 28756 78036 29036
rect 77980 28690 78036 28700
rect 78092 28532 78148 29260
rect 78092 28466 78148 28476
rect 77756 28130 77812 28140
rect 77868 28420 77924 28430
rect 77756 27972 77812 27982
rect 77868 27972 77924 28364
rect 77756 27970 77924 27972
rect 77756 27918 77758 27970
rect 77810 27918 77924 27970
rect 77756 27916 77924 27918
rect 77980 28308 78036 28318
rect 77756 27906 77812 27916
rect 77868 27748 77924 27758
rect 77980 27748 78036 28252
rect 77644 27692 77812 27748
rect 77532 27634 77588 27646
rect 77532 27582 77534 27634
rect 77586 27582 77588 27634
rect 77532 27300 77588 27582
rect 77532 27234 77588 27244
rect 77420 27020 77588 27076
rect 77308 27010 77364 27020
rect 77308 26628 77364 26638
rect 77308 26178 77364 26572
rect 77308 26126 77310 26178
rect 77362 26126 77364 26178
rect 77308 26114 77364 26126
rect 77420 26290 77476 26302
rect 77420 26238 77422 26290
rect 77474 26238 77476 26290
rect 77308 25732 77364 25742
rect 77308 25638 77364 25676
rect 77420 25620 77476 26238
rect 77420 25488 77476 25564
rect 77532 25060 77588 27020
rect 77644 26964 77700 26974
rect 77644 26870 77700 26908
rect 77756 26178 77812 27692
rect 77868 27746 78036 27748
rect 77868 27694 77870 27746
rect 77922 27694 78036 27746
rect 77868 27692 78036 27694
rect 78092 28196 78148 28206
rect 77868 27682 77924 27692
rect 77980 27524 78036 27534
rect 77756 26126 77758 26178
rect 77810 26126 77812 26178
rect 77756 26114 77812 26126
rect 77868 26628 77924 26638
rect 77308 25004 77588 25060
rect 77756 25956 77812 25966
rect 77308 24050 77364 25004
rect 77532 24834 77588 24846
rect 77532 24782 77534 24834
rect 77586 24782 77588 24834
rect 77532 24724 77588 24782
rect 77644 24836 77700 24846
rect 77644 24742 77700 24780
rect 77532 24658 77588 24668
rect 77308 23998 77310 24050
rect 77362 23998 77364 24050
rect 77308 23940 77364 23998
rect 77308 23874 77364 23884
rect 77420 24612 77476 24622
rect 77420 22482 77476 24556
rect 77532 24500 77588 24510
rect 77756 24500 77812 25900
rect 77868 25618 77924 26572
rect 77868 25566 77870 25618
rect 77922 25566 77924 25618
rect 77868 25554 77924 25566
rect 77532 24498 77812 24500
rect 77532 24446 77534 24498
rect 77586 24446 77812 24498
rect 77532 24444 77812 24446
rect 77532 24434 77588 24444
rect 77980 22596 78036 27468
rect 78092 27188 78148 28140
rect 78092 27056 78148 27132
rect 77420 22430 77422 22482
rect 77474 22430 77476 22482
rect 77420 22418 77476 22430
rect 77644 22540 78036 22596
rect 77532 22260 77588 22270
rect 77532 22166 77588 22204
rect 77308 22146 77364 22158
rect 77308 22094 77310 22146
rect 77362 22094 77364 22146
rect 77308 21700 77364 22094
rect 77308 21634 77364 21644
rect 77532 20916 77588 20926
rect 77532 20822 77588 20860
rect 77308 20802 77364 20814
rect 77308 20750 77310 20802
rect 77362 20750 77364 20802
rect 77308 20580 77364 20750
rect 77308 20514 77364 20524
rect 77532 20132 77588 20142
rect 77532 20038 77588 20076
rect 77308 19348 77364 19358
rect 77196 19346 77364 19348
rect 77196 19294 77310 19346
rect 77362 19294 77364 19346
rect 77196 19292 77364 19294
rect 77196 19236 77252 19292
rect 77308 19282 77364 19292
rect 77196 19170 77252 19180
rect 77644 18674 77700 22540
rect 77756 22148 77812 22158
rect 77756 22054 77812 22092
rect 77868 20804 77924 20814
rect 77868 20710 77924 20748
rect 77644 18622 77646 18674
rect 77698 18622 77700 18674
rect 77644 18610 77700 18622
rect 76524 18508 76692 18564
rect 77532 18564 77588 18574
rect 76076 18450 76132 18462
rect 76076 18398 76078 18450
rect 76130 18398 76132 18450
rect 76076 18340 76132 18398
rect 76076 18274 76132 18284
rect 76076 17668 76132 17678
rect 76076 17574 76132 17612
rect 76076 16884 76132 16922
rect 76076 16818 76132 16828
rect 75964 16482 76020 16492
rect 76076 16660 76132 16670
rect 75516 16158 75518 16210
rect 75570 16158 75572 16210
rect 75516 16146 75572 16158
rect 75964 16100 76020 16110
rect 75964 16006 76020 16044
rect 76076 15986 76132 16604
rect 76300 16100 76356 16110
rect 76524 16100 76580 18508
rect 77532 18470 77588 18508
rect 77756 18562 77812 18574
rect 77756 18510 77758 18562
rect 77810 18510 77812 18562
rect 76748 18452 76804 18462
rect 76748 18358 76804 18396
rect 77756 18452 77812 18510
rect 78092 18452 78148 18462
rect 77420 18340 77476 18350
rect 77308 17780 77364 17790
rect 76748 17668 76804 17678
rect 76748 16994 76804 17612
rect 77308 17666 77364 17724
rect 77308 17614 77310 17666
rect 77362 17614 77364 17666
rect 77308 17602 77364 17614
rect 77420 17554 77476 18284
rect 77756 17892 77812 18396
rect 77420 17502 77422 17554
rect 77474 17502 77476 17554
rect 77420 17332 77476 17502
rect 77420 17266 77476 17276
rect 77532 17836 77812 17892
rect 77868 18450 78148 18452
rect 77868 18398 78094 18450
rect 78146 18398 78148 18450
rect 77868 18396 78148 18398
rect 76748 16942 76750 16994
rect 76802 16942 76804 16994
rect 76748 16930 76804 16942
rect 77420 16882 77476 16894
rect 77420 16830 77422 16882
rect 77474 16830 77476 16882
rect 77084 16770 77140 16782
rect 77084 16718 77086 16770
rect 77138 16718 77140 16770
rect 76300 16098 76580 16100
rect 76300 16046 76302 16098
rect 76354 16046 76580 16098
rect 76300 16044 76580 16046
rect 76636 16660 76692 16670
rect 76300 16034 76356 16044
rect 76076 15934 76078 15986
rect 76130 15934 76132 15986
rect 76076 15922 76132 15934
rect 75404 15408 75460 15484
rect 76188 15540 76244 15550
rect 76188 15314 76244 15484
rect 76188 15262 76190 15314
rect 76242 15262 76244 15314
rect 76188 15250 76244 15262
rect 76636 15148 76692 16604
rect 77084 16100 77140 16718
rect 77420 16660 77476 16830
rect 77420 16594 77476 16604
rect 77420 16324 77476 16334
rect 77532 16324 77588 17836
rect 77644 17668 77700 17678
rect 77868 17668 77924 18396
rect 78092 18386 78148 18396
rect 77644 17666 77924 17668
rect 77644 17614 77646 17666
rect 77698 17614 77924 17666
rect 77644 17612 77924 17614
rect 77644 17602 77700 17612
rect 77980 17442 78036 17454
rect 77980 17390 77982 17442
rect 78034 17390 78036 17442
rect 77420 16322 77588 16324
rect 77420 16270 77422 16322
rect 77474 16270 77588 16322
rect 77420 16268 77588 16270
rect 77756 17332 77812 17342
rect 77420 16258 77476 16268
rect 77084 16034 77140 16044
rect 76748 15988 76804 15998
rect 76748 15316 76804 15932
rect 77308 15988 77364 15998
rect 77308 15894 77364 15932
rect 77420 15874 77476 15886
rect 77420 15822 77422 15874
rect 77474 15822 77476 15874
rect 77420 15540 77476 15822
rect 77420 15474 77476 15484
rect 76748 15250 76804 15260
rect 76860 15428 76916 15438
rect 76188 15092 76244 15102
rect 76636 15092 76804 15148
rect 74844 11454 74846 11506
rect 74898 11454 74900 11506
rect 74844 11442 74900 11454
rect 75180 13916 75348 13972
rect 76076 14418 76132 14430
rect 76076 14366 76078 14418
rect 76130 14366 76132 14418
rect 74956 11396 75012 11406
rect 74956 11302 75012 11340
rect 74732 11172 74788 11182
rect 74732 10836 74788 11116
rect 74732 10770 74788 10780
rect 74844 10612 74900 10622
rect 74844 10518 74900 10556
rect 74956 10500 75012 10510
rect 74956 10406 75012 10444
rect 74956 9940 75012 9950
rect 74620 9884 74956 9940
rect 74956 9808 75012 9884
rect 74620 9602 74676 9614
rect 74620 9550 74622 9602
rect 74674 9550 74676 9602
rect 74508 8930 74564 8942
rect 74508 8878 74510 8930
rect 74562 8878 74564 8930
rect 74508 8428 74564 8878
rect 73948 8372 74116 8428
rect 74396 8372 74564 8428
rect 74620 8428 74676 9550
rect 75180 9268 75236 13916
rect 75404 13860 75460 13870
rect 76076 13860 76132 14366
rect 75404 13858 75572 13860
rect 75404 13806 75406 13858
rect 75458 13806 75572 13858
rect 75404 13804 75572 13806
rect 75404 13794 75460 13804
rect 75292 13746 75348 13758
rect 75292 13694 75294 13746
rect 75346 13694 75348 13746
rect 75292 13412 75348 13694
rect 75404 13524 75460 13534
rect 75404 13430 75460 13468
rect 75292 13346 75348 13356
rect 75516 13188 75572 13804
rect 76076 13794 76132 13804
rect 76188 13634 76244 15036
rect 76188 13582 76190 13634
rect 76242 13582 76244 13634
rect 76188 13570 76244 13582
rect 76412 13636 76468 13646
rect 75516 13122 75572 13132
rect 76300 13412 76356 13422
rect 76076 12964 76132 12974
rect 76076 12870 76132 12908
rect 76300 12962 76356 13356
rect 76412 13186 76468 13580
rect 76748 13412 76804 15092
rect 76860 13746 76916 15372
rect 77532 15428 77588 15438
rect 77532 15334 77588 15372
rect 77420 15314 77476 15326
rect 77420 15262 77422 15314
rect 77474 15262 77476 15314
rect 77420 15148 77476 15262
rect 76860 13694 76862 13746
rect 76914 13694 76916 13746
rect 76860 13682 76916 13694
rect 77308 15092 77476 15148
rect 77532 15092 77588 15102
rect 76972 13636 77028 13646
rect 77308 13636 77364 15092
rect 77532 15090 77700 15092
rect 77532 15038 77534 15090
rect 77586 15038 77700 15090
rect 77532 15036 77700 15038
rect 77532 15026 77588 15036
rect 77420 14756 77476 14766
rect 77420 14662 77476 14700
rect 77532 14532 77588 14542
rect 77644 14532 77700 15036
rect 77756 14756 77812 17276
rect 77980 16660 78036 17390
rect 77980 16210 78036 16604
rect 77980 16158 77982 16210
rect 78034 16158 78036 16210
rect 77980 16146 78036 16158
rect 78092 15540 78148 15550
rect 78092 15446 78148 15484
rect 78204 14980 78260 31724
rect 78492 31388 78756 31398
rect 78548 31332 78596 31388
rect 78652 31332 78700 31388
rect 78492 31322 78756 31332
rect 78492 29820 78756 29830
rect 78548 29764 78596 29820
rect 78652 29764 78700 29820
rect 78492 29754 78756 29764
rect 78316 28532 78372 28542
rect 78316 26516 78372 28476
rect 78492 28252 78756 28262
rect 78548 28196 78596 28252
rect 78652 28196 78700 28252
rect 78492 28186 78756 28196
rect 78492 26684 78756 26694
rect 78548 26628 78596 26684
rect 78652 26628 78700 26684
rect 78492 26618 78756 26628
rect 78316 26450 78372 26460
rect 78492 25116 78756 25126
rect 78548 25060 78596 25116
rect 78652 25060 78700 25116
rect 78492 25050 78756 25060
rect 78492 23548 78756 23558
rect 78548 23492 78596 23548
rect 78652 23492 78700 23548
rect 78492 23482 78756 23492
rect 77756 14690 77812 14700
rect 77868 14924 78260 14980
rect 78316 23268 78372 23278
rect 77532 14530 77700 14532
rect 77532 14478 77534 14530
rect 77586 14478 77700 14530
rect 77532 14476 77700 14478
rect 77532 14466 77588 14476
rect 77028 13580 77364 13636
rect 77420 14306 77476 14318
rect 77420 14254 77422 14306
rect 77474 14254 77476 14306
rect 76972 13504 77028 13580
rect 77420 13524 77476 14254
rect 77420 13458 77476 13468
rect 76748 13356 77140 13412
rect 76412 13134 76414 13186
rect 76466 13134 76468 13186
rect 76412 13122 76468 13134
rect 76300 12910 76302 12962
rect 76354 12910 76356 12962
rect 76300 12292 76356 12910
rect 76748 12292 76804 12302
rect 76300 12236 76692 12292
rect 76188 12180 76244 12190
rect 76188 12086 76244 12124
rect 75516 12066 75572 12078
rect 75516 12014 75518 12066
rect 75570 12014 75572 12066
rect 75516 11508 75572 12014
rect 75516 11442 75572 11452
rect 76188 11956 76244 11966
rect 75628 11396 75684 11406
rect 75628 10500 75684 11340
rect 75852 11394 75908 11406
rect 75852 11342 75854 11394
rect 75906 11342 75908 11394
rect 75852 11172 75908 11342
rect 75852 11106 75908 11116
rect 75740 10724 75796 10734
rect 75740 10630 75796 10668
rect 75628 10434 75684 10444
rect 75516 9604 75572 9614
rect 75180 9202 75236 9212
rect 75292 9602 75572 9604
rect 75292 9550 75518 9602
rect 75570 9550 75572 9602
rect 75292 9548 75572 9550
rect 74956 9044 75012 9054
rect 74620 8372 74900 8428
rect 73388 8194 73444 8204
rect 73612 8260 73668 8270
rect 73612 8166 73668 8204
rect 73276 7812 73332 7822
rect 73276 7698 73332 7756
rect 73276 7646 73278 7698
rect 73330 7646 73332 7698
rect 73276 7634 73332 7646
rect 73836 7362 73892 7374
rect 73836 7310 73838 7362
rect 73890 7310 73892 7362
rect 73836 7250 73892 7310
rect 73836 7198 73838 7250
rect 73890 7198 73892 7250
rect 73164 6692 73220 6702
rect 73164 6132 73220 6636
rect 73612 6466 73668 6478
rect 73612 6414 73614 6466
rect 73666 6414 73668 6466
rect 73612 6356 73668 6414
rect 73612 6290 73668 6300
rect 73276 6132 73332 6142
rect 73164 6130 73332 6132
rect 73164 6078 73278 6130
rect 73330 6078 73332 6130
rect 73164 6076 73332 6078
rect 73276 6066 73332 6076
rect 73052 5852 73220 5908
rect 72492 5346 72548 5852
rect 72604 5796 72660 5806
rect 72604 5702 72660 5740
rect 72492 5294 72494 5346
rect 72546 5294 72548 5346
rect 72492 5282 72548 5294
rect 72044 4114 72212 4116
rect 72044 4062 72046 4114
rect 72098 4062 72212 4114
rect 72044 4060 72212 4062
rect 72380 4900 72436 4910
rect 72380 4340 72436 4844
rect 73052 4898 73108 4910
rect 73052 4846 73054 4898
rect 73106 4846 73108 4898
rect 73052 4788 73108 4846
rect 73052 4722 73108 4732
rect 72604 4564 72660 4574
rect 72604 4470 72660 4508
rect 72044 4050 72100 4060
rect 72380 3666 72436 4284
rect 72380 3614 72382 3666
rect 72434 3614 72436 3666
rect 72380 3602 72436 3614
rect 71932 3266 71988 3276
rect 73164 3330 73220 5852
rect 73500 5684 73556 5694
rect 73388 5236 73444 5246
rect 73276 4564 73332 4574
rect 73276 4470 73332 4508
rect 73388 3556 73444 5180
rect 73500 5234 73556 5628
rect 73836 5572 73892 7198
rect 73948 6244 74004 8372
rect 74172 8036 74228 8046
rect 74172 8034 74340 8036
rect 74172 7982 74174 8034
rect 74226 7982 74340 8034
rect 74172 7980 74340 7982
rect 74172 7970 74228 7980
rect 74172 7362 74228 7374
rect 74172 7310 74174 7362
rect 74226 7310 74228 7362
rect 74172 7250 74228 7310
rect 74172 7198 74174 7250
rect 74226 7198 74228 7250
rect 74172 7186 74228 7198
rect 74284 6804 74340 7980
rect 74060 6468 74116 6478
rect 74060 6374 74116 6412
rect 73948 6188 74116 6244
rect 73836 5506 73892 5516
rect 73500 5182 73502 5234
rect 73554 5182 73556 5234
rect 73500 5170 73556 5182
rect 73948 5124 74004 5134
rect 73948 5030 74004 5068
rect 74060 4562 74116 6188
rect 74284 6130 74340 6748
rect 74284 6078 74286 6130
rect 74338 6078 74340 6130
rect 74060 4510 74062 4562
rect 74114 4510 74116 4562
rect 74060 4498 74116 4510
rect 74172 5906 74228 5918
rect 74172 5854 74174 5906
rect 74226 5854 74228 5906
rect 74172 5012 74228 5854
rect 74284 5348 74340 6078
rect 74284 5282 74340 5292
rect 74396 5124 74452 8372
rect 74620 8260 74676 8270
rect 74620 8166 74676 8204
rect 74732 8036 74788 8046
rect 74732 7942 74788 7980
rect 74732 7362 74788 7374
rect 74732 7310 74734 7362
rect 74786 7310 74788 7362
rect 74620 6468 74676 6478
rect 74508 6132 74564 6142
rect 74508 6038 74564 6076
rect 74172 4116 74228 4956
rect 74284 5068 74452 5124
rect 74284 4340 74340 5068
rect 74396 4900 74452 4910
rect 74396 4806 74452 4844
rect 74620 4564 74676 6412
rect 74732 5012 74788 7310
rect 74732 4946 74788 4956
rect 74620 4498 74676 4508
rect 74396 4340 74452 4350
rect 74284 4338 74452 4340
rect 74284 4286 74398 4338
rect 74450 4286 74452 4338
rect 74284 4284 74452 4286
rect 74172 4050 74228 4060
rect 73164 3278 73166 3330
rect 73218 3278 73220 3330
rect 73164 3266 73220 3278
rect 73276 3554 73444 3556
rect 73276 3502 73390 3554
rect 73442 3502 73444 3554
rect 73276 3500 73444 3502
rect 73276 980 73332 3500
rect 73388 3490 73444 3500
rect 72940 924 73332 980
rect 72940 800 72996 924
rect 15708 700 16324 756
rect 17584 0 17696 800
rect 19712 0 19824 800
rect 21840 0 21952 800
rect 23968 0 24080 800
rect 26096 0 26208 800
rect 28224 0 28336 800
rect 30352 0 30464 800
rect 32480 0 32592 800
rect 34608 0 34720 800
rect 36736 0 36848 800
rect 38864 0 38976 800
rect 40992 0 41104 800
rect 43120 0 43232 800
rect 45248 0 45360 800
rect 47376 0 47488 800
rect 49504 0 49616 800
rect 51632 0 51744 800
rect 53760 0 53872 800
rect 55888 0 56000 800
rect 58016 0 58128 800
rect 60144 0 60256 800
rect 62272 0 62384 800
rect 64400 0 64512 800
rect 66528 0 66640 800
rect 68656 0 68768 800
rect 70784 0 70896 800
rect 72912 0 73024 800
rect 74396 756 74452 4284
rect 74844 3892 74900 8372
rect 74956 8258 75012 8988
rect 74956 8206 74958 8258
rect 75010 8206 75012 8258
rect 74956 8194 75012 8206
rect 75292 8148 75348 9548
rect 75516 9538 75572 9548
rect 75852 9602 75908 9614
rect 75852 9550 75854 9602
rect 75906 9550 75908 9602
rect 75852 9380 75908 9550
rect 75852 9314 75908 9324
rect 75964 9268 76020 9278
rect 75628 9156 75684 9166
rect 75516 8932 75572 8942
rect 75516 8838 75572 8876
rect 75404 8372 75460 8382
rect 75404 8278 75460 8316
rect 75516 8260 75572 8270
rect 75516 8166 75572 8204
rect 75292 8082 75348 8092
rect 75628 8036 75684 9100
rect 75964 9042 76020 9212
rect 75964 8990 75966 9042
rect 76018 8990 76020 9042
rect 75964 8978 76020 8990
rect 75516 7980 75684 8036
rect 75964 8258 76020 8270
rect 75964 8206 75966 8258
rect 76018 8206 76020 8258
rect 75964 8036 76020 8206
rect 75516 7698 75572 7980
rect 75516 7646 75518 7698
rect 75570 7646 75572 7698
rect 75516 7634 75572 7646
rect 75292 7586 75348 7598
rect 75292 7534 75294 7586
rect 75346 7534 75348 7586
rect 75180 7474 75236 7486
rect 75180 7422 75182 7474
rect 75234 7422 75236 7474
rect 75068 6578 75124 6590
rect 75068 6526 75070 6578
rect 75122 6526 75124 6578
rect 75068 6468 75124 6526
rect 75068 6402 75124 6412
rect 75068 5796 75124 5806
rect 75180 5796 75236 7422
rect 75292 6692 75348 7534
rect 75292 5906 75348 6636
rect 75964 6018 76020 7980
rect 76076 6804 76132 6814
rect 76076 6690 76132 6748
rect 76076 6638 76078 6690
rect 76130 6638 76132 6690
rect 76076 6626 76132 6638
rect 75964 5966 75966 6018
rect 76018 5966 76020 6018
rect 75964 5954 76020 5966
rect 75292 5854 75294 5906
rect 75346 5854 75348 5906
rect 75292 5842 75348 5854
rect 75124 5740 75236 5796
rect 75068 5702 75124 5740
rect 75516 5348 75572 5358
rect 76188 5348 76244 11900
rect 76524 11508 76580 11518
rect 76524 11414 76580 11452
rect 76412 10724 76468 10734
rect 76412 10610 76468 10668
rect 76412 10558 76414 10610
rect 76466 10558 76468 10610
rect 76300 10500 76356 10510
rect 76300 10406 76356 10444
rect 76412 9938 76468 10558
rect 76524 10612 76580 10622
rect 76524 10050 76580 10556
rect 76524 9998 76526 10050
rect 76578 9998 76580 10050
rect 76524 9986 76580 9998
rect 76412 9886 76414 9938
rect 76466 9886 76468 9938
rect 76412 9874 76468 9886
rect 76636 8372 76692 12236
rect 76748 12198 76804 12236
rect 76972 11284 77028 11294
rect 76748 10610 76804 10622
rect 76748 10558 76750 10610
rect 76802 10558 76804 10610
rect 76748 9380 76804 10558
rect 76748 9314 76804 9324
rect 76860 9156 76916 9166
rect 76860 9062 76916 9100
rect 76748 9044 76804 9054
rect 76748 8950 76804 8988
rect 76636 8306 76692 8316
rect 76860 8260 76916 8270
rect 76300 8148 76356 8158
rect 76300 7474 76356 8092
rect 76860 7476 76916 8204
rect 76972 7586 77028 11228
rect 77084 9266 77140 13356
rect 77308 13188 77364 13198
rect 77308 13094 77364 13132
rect 77868 13074 77924 14924
rect 78316 14420 78372 23212
rect 78492 21980 78756 21990
rect 78548 21924 78596 21980
rect 78652 21924 78700 21980
rect 78492 21914 78756 21924
rect 78492 20412 78756 20422
rect 78548 20356 78596 20412
rect 78652 20356 78700 20412
rect 78492 20346 78756 20356
rect 78492 18844 78756 18854
rect 78548 18788 78596 18844
rect 78652 18788 78700 18844
rect 78492 18778 78756 18788
rect 78876 17444 78932 34188
rect 79100 28084 79156 28094
rect 78988 26964 79044 26974
rect 78988 20132 79044 26908
rect 78988 20066 79044 20076
rect 78876 17378 78932 17388
rect 78492 17276 78756 17286
rect 78548 17220 78596 17276
rect 78652 17220 78700 17276
rect 78492 17210 78756 17220
rect 78492 15708 78756 15718
rect 78548 15652 78596 15708
rect 78652 15652 78700 15708
rect 78492 15642 78756 15652
rect 77868 13022 77870 13074
rect 77922 13022 77924 13074
rect 77420 12964 77476 12974
rect 77420 12850 77476 12908
rect 77420 12798 77422 12850
rect 77474 12798 77476 12850
rect 77196 12178 77252 12190
rect 77196 12126 77198 12178
rect 77250 12126 77252 12178
rect 77196 11284 77252 12126
rect 77420 11506 77476 12798
rect 77868 12180 77924 13022
rect 77868 12114 77924 12124
rect 78092 14364 78372 14420
rect 77420 11454 77422 11506
rect 77474 11454 77476 11506
rect 77420 11442 77476 11454
rect 77532 12066 77588 12078
rect 77532 12014 77534 12066
rect 77586 12014 77588 12066
rect 77532 11508 77588 12014
rect 77196 11218 77252 11228
rect 77308 11284 77364 11294
rect 77532 11284 77588 11452
rect 77756 11394 77812 11406
rect 77756 11342 77758 11394
rect 77810 11342 77812 11394
rect 77308 11282 77588 11284
rect 77308 11230 77310 11282
rect 77362 11230 77588 11282
rect 77308 11228 77588 11230
rect 77644 11284 77700 11294
rect 77308 11218 77364 11228
rect 77644 11190 77700 11228
rect 77532 10724 77588 10734
rect 77532 9602 77588 10668
rect 77532 9550 77534 9602
rect 77586 9550 77588 9602
rect 77532 9380 77588 9550
rect 77532 9314 77588 9324
rect 77644 10050 77700 10062
rect 77644 9998 77646 10050
rect 77698 9998 77700 10050
rect 77084 9214 77086 9266
rect 77138 9214 77140 9266
rect 77084 9202 77140 9214
rect 77420 9268 77476 9278
rect 77420 9174 77476 9212
rect 77308 8372 77364 8382
rect 77308 8258 77364 8316
rect 77308 8206 77310 8258
rect 77362 8206 77364 8258
rect 77308 8148 77364 8206
rect 77532 8260 77588 8270
rect 77532 8166 77588 8204
rect 77308 8082 77364 8092
rect 76972 7534 76974 7586
rect 77026 7534 77028 7586
rect 76972 7522 77028 7534
rect 77532 7586 77588 7598
rect 77532 7534 77534 7586
rect 77586 7534 77588 7586
rect 76300 7422 76302 7474
rect 76354 7422 76356 7474
rect 76300 7410 76356 7422
rect 76524 7474 76916 7476
rect 76524 7422 76862 7474
rect 76914 7422 76916 7474
rect 76524 7420 76916 7422
rect 76524 6018 76580 7420
rect 76860 7410 76916 7420
rect 77532 6804 77588 7534
rect 77532 6738 77588 6748
rect 77420 6692 77476 6702
rect 77420 6598 77476 6636
rect 76524 5966 76526 6018
rect 76578 5966 76580 6018
rect 76524 5954 76580 5966
rect 77308 6580 77364 6590
rect 76972 5908 77028 5918
rect 75516 5124 75572 5292
rect 76076 5292 76244 5348
rect 76300 5348 76356 5358
rect 75516 4992 75572 5068
rect 75628 5234 75684 5246
rect 75628 5182 75630 5234
rect 75682 5182 75684 5234
rect 75628 5012 75684 5182
rect 75628 4946 75684 4956
rect 75516 4226 75572 4238
rect 75516 4174 75518 4226
rect 75570 4174 75572 4226
rect 75516 4004 75572 4174
rect 76076 4116 76132 5292
rect 76300 5254 76356 5292
rect 76972 5348 77028 5852
rect 77308 5794 77364 6524
rect 77532 6466 77588 6478
rect 77532 6414 77534 6466
rect 77586 6414 77588 6466
rect 77532 5908 77588 6414
rect 77532 5842 77588 5852
rect 77308 5742 77310 5794
rect 77362 5742 77364 5794
rect 77308 5730 77364 5742
rect 77644 5684 77700 9998
rect 77756 8372 77812 11342
rect 78092 10948 78148 14364
rect 79100 14308 79156 28028
rect 77868 10892 78148 10948
rect 78204 14252 79156 14308
rect 77868 10050 77924 10892
rect 77980 10724 78036 10734
rect 77980 10630 78036 10668
rect 78092 10612 78148 10622
rect 78092 10518 78148 10556
rect 77980 10388 78036 10398
rect 77980 10294 78036 10332
rect 77868 9998 77870 10050
rect 77922 9998 77924 10050
rect 77868 9940 77924 9998
rect 77980 9940 78036 9950
rect 77868 9938 78036 9940
rect 77868 9886 77982 9938
rect 78034 9886 78036 9938
rect 77868 9884 78036 9886
rect 77980 9874 78036 9884
rect 77868 8930 77924 8942
rect 77868 8878 77870 8930
rect 77922 8878 77924 8930
rect 77868 8596 77924 8878
rect 77868 8530 77924 8540
rect 78204 8428 78260 14252
rect 78492 14140 78756 14150
rect 78548 14084 78596 14140
rect 78652 14084 78700 14140
rect 78492 14074 78756 14084
rect 78492 12572 78756 12582
rect 78548 12516 78596 12572
rect 78652 12516 78700 12572
rect 78492 12506 78756 12516
rect 78492 11004 78756 11014
rect 78548 10948 78596 11004
rect 78652 10948 78700 11004
rect 78492 10938 78756 10948
rect 77868 8372 77924 8382
rect 77756 8370 77924 8372
rect 77756 8318 77870 8370
rect 77922 8318 77924 8370
rect 77756 8316 77924 8318
rect 77868 8306 77924 8316
rect 77980 8372 78260 8428
rect 78316 9940 78372 9950
rect 77868 7588 77924 7598
rect 77980 7588 78036 8372
rect 77868 7586 78036 7588
rect 77868 7534 77870 7586
rect 77922 7534 78036 7586
rect 77868 7532 78036 7534
rect 77868 7522 77924 7532
rect 77756 6466 77812 6478
rect 77756 6414 77758 6466
rect 77810 6414 77812 6466
rect 77756 6132 77812 6414
rect 77756 6066 77812 6076
rect 77980 6130 78036 7532
rect 77980 6078 77982 6130
rect 78034 6078 78036 6130
rect 77980 6066 78036 6078
rect 76972 5282 77028 5292
rect 77532 5628 77700 5684
rect 77196 5236 77252 5246
rect 77196 5142 77252 5180
rect 76748 4450 76804 4462
rect 76748 4398 76750 4450
rect 76802 4398 76804 4450
rect 76188 4340 76244 4350
rect 76748 4340 76804 4398
rect 77084 4452 77140 4462
rect 77532 4452 77588 5628
rect 77644 5122 77700 5134
rect 77644 5070 77646 5122
rect 77698 5070 77700 5122
rect 77644 5012 77700 5070
rect 78092 5124 78148 5134
rect 78092 5030 78148 5068
rect 77644 4946 77700 4956
rect 77084 4450 77588 4452
rect 77084 4398 77086 4450
rect 77138 4398 77588 4450
rect 77084 4396 77588 4398
rect 77644 4450 77700 4462
rect 77644 4398 77646 4450
rect 77698 4398 77700 4450
rect 77084 4386 77140 4396
rect 76188 4338 76804 4340
rect 76188 4286 76190 4338
rect 76242 4286 76804 4338
rect 76188 4284 76804 4286
rect 76188 4274 76244 4284
rect 76076 4060 76356 4116
rect 75516 3938 75572 3948
rect 74844 3826 74900 3836
rect 74844 3666 74900 3678
rect 74844 3614 74846 3666
rect 74898 3614 74900 3666
rect 74844 1540 74900 3614
rect 76300 3666 76356 4060
rect 76300 3614 76302 3666
rect 76354 3614 76356 3666
rect 76300 3602 76356 3614
rect 76748 3892 76804 3902
rect 75516 3556 75572 3566
rect 75516 3462 75572 3500
rect 76748 3554 76804 3836
rect 76748 3502 76750 3554
rect 76802 3502 76804 3554
rect 76748 3490 76804 3502
rect 77196 3892 77252 3902
rect 74844 1474 74900 1484
rect 74844 924 75124 980
rect 74844 756 74900 924
rect 75068 800 75124 924
rect 77196 800 77252 3836
rect 77308 3668 77364 3678
rect 77308 3574 77364 3612
rect 77644 3556 77700 4398
rect 77980 4452 78036 4462
rect 78316 4452 78372 9884
rect 78492 9436 78756 9446
rect 78548 9380 78596 9436
rect 78652 9380 78700 9436
rect 78492 9370 78756 9380
rect 78492 7868 78756 7878
rect 78548 7812 78596 7868
rect 78652 7812 78700 7868
rect 78492 7802 78756 7812
rect 78492 6300 78756 6310
rect 78548 6244 78596 6300
rect 78652 6244 78700 6300
rect 78492 6234 78756 6244
rect 78492 4732 78756 4742
rect 78548 4676 78596 4732
rect 78652 4676 78700 4732
rect 78492 4666 78756 4676
rect 77980 4450 78372 4452
rect 77980 4398 77982 4450
rect 78034 4398 78372 4450
rect 77980 4396 78372 4398
rect 77980 4386 78036 4396
rect 77644 3490 77700 3500
rect 77756 3444 77812 3454
rect 77756 3350 77812 3388
rect 78492 3164 78756 3174
rect 78548 3108 78596 3164
rect 78652 3108 78700 3164
rect 78492 3098 78756 3108
rect 74396 700 74900 756
rect 75040 0 75152 800
rect 77168 0 77280 800
<< via2 >>
rect 2156 38444 2212 38500
rect 1932 35980 1988 36036
rect 2492 37660 2548 37716
rect 2268 37436 2324 37492
rect 1932 33516 1988 33572
rect 1596 31164 1652 31220
rect 1484 29708 1540 29764
rect 1372 25676 1428 25732
rect 1372 7532 1428 7588
rect 1484 5068 1540 5124
rect 1932 31052 1988 31108
rect 1932 28588 1988 28644
rect 1932 26178 1988 26180
rect 1932 26126 1934 26178
rect 1934 26126 1986 26178
rect 1986 26126 1988 26178
rect 1932 26124 1988 26126
rect 1932 23660 1988 23716
rect 2044 21756 2100 21812
rect 2156 21644 2212 21700
rect 1932 21196 1988 21252
rect 2380 29986 2436 29988
rect 2380 29934 2382 29986
rect 2382 29934 2434 29986
rect 2434 29934 2436 29986
rect 2380 29932 2436 29934
rect 5068 37100 5124 37156
rect 3164 36482 3220 36484
rect 3164 36430 3166 36482
rect 3166 36430 3218 36482
rect 3218 36430 3220 36482
rect 3164 36428 3220 36430
rect 4956 35868 5012 35924
rect 3052 35756 3108 35812
rect 3612 35810 3668 35812
rect 3612 35758 3614 35810
rect 3614 35758 3666 35810
rect 3666 35758 3668 35810
rect 3612 35756 3668 35758
rect 3948 35532 4004 35588
rect 3052 35308 3108 35364
rect 4844 35810 4900 35812
rect 4844 35758 4846 35810
rect 4846 35758 4898 35810
rect 4898 35758 4900 35810
rect 4844 35756 4900 35758
rect 4508 35308 4564 35364
rect 7084 36988 7140 37044
rect 6076 36428 6132 36484
rect 5292 36316 5348 36372
rect 5628 35868 5684 35924
rect 5292 35756 5348 35812
rect 4844 35532 4900 35588
rect 3948 34972 4004 35028
rect 4396 35026 4452 35028
rect 4396 34974 4398 35026
rect 4398 34974 4450 35026
rect 4450 34974 4452 35026
rect 4396 34972 4452 34974
rect 3052 34636 3108 34692
rect 3612 34690 3668 34692
rect 3612 34638 3614 34690
rect 3614 34638 3666 34690
rect 3666 34638 3668 34690
rect 3612 34636 3668 34638
rect 3724 33516 3780 33572
rect 3164 33404 3220 33460
rect 3612 33458 3668 33460
rect 3612 33406 3614 33458
rect 3614 33406 3666 33458
rect 3666 33406 3668 33458
rect 3612 33404 3668 33406
rect 3052 31612 3108 31668
rect 3500 31666 3556 31668
rect 3500 31614 3502 31666
rect 3502 31614 3554 31666
rect 3554 31614 3556 31666
rect 3500 31612 3556 31614
rect 4172 31500 4228 31556
rect 4508 30994 4564 30996
rect 4508 30942 4510 30994
rect 4510 30942 4562 30994
rect 4562 30942 4564 30994
rect 4508 30940 4564 30942
rect 9996 37548 10052 37604
rect 10872 36874 10928 36876
rect 10872 36822 10874 36874
rect 10874 36822 10926 36874
rect 10926 36822 10928 36874
rect 10872 36820 10928 36822
rect 10976 36874 11032 36876
rect 10976 36822 10978 36874
rect 10978 36822 11030 36874
rect 11030 36822 11032 36874
rect 10976 36820 11032 36822
rect 11080 36874 11136 36876
rect 11080 36822 11082 36874
rect 11082 36822 11134 36874
rect 11134 36822 11136 36874
rect 11080 36820 11136 36822
rect 15484 37212 15540 37268
rect 9996 36316 10052 36372
rect 8092 36092 8148 36148
rect 8540 36092 8596 36148
rect 7084 34972 7140 35028
rect 11900 35756 11956 35812
rect 11004 35698 11060 35700
rect 11004 35646 11006 35698
rect 11006 35646 11058 35698
rect 11058 35646 11060 35698
rect 11004 35644 11060 35646
rect 12012 35644 12068 35700
rect 8988 34860 9044 34916
rect 9772 34636 9828 34692
rect 6748 32732 6804 32788
rect 8764 33852 8820 33908
rect 7644 33068 7700 33124
rect 7420 32786 7476 32788
rect 7420 32734 7422 32786
rect 7422 32734 7474 32786
rect 7474 32734 7476 32786
rect 7420 32732 7476 32734
rect 7308 32674 7364 32676
rect 7308 32622 7310 32674
rect 7310 32622 7362 32674
rect 7362 32622 7364 32674
rect 7308 32620 7364 32622
rect 8988 33292 9044 33348
rect 8316 32844 8372 32900
rect 8204 32786 8260 32788
rect 8204 32734 8206 32786
rect 8206 32734 8258 32786
rect 8258 32734 8260 32786
rect 8204 32732 8260 32734
rect 8092 32674 8148 32676
rect 8092 32622 8094 32674
rect 8094 32622 8146 32674
rect 8146 32622 8148 32674
rect 8092 32620 8148 32622
rect 7196 32396 7252 32452
rect 7644 32508 7700 32564
rect 8316 32620 8372 32676
rect 10872 35306 10928 35308
rect 10872 35254 10874 35306
rect 10874 35254 10926 35306
rect 10926 35254 10928 35306
rect 10872 35252 10928 35254
rect 10976 35306 11032 35308
rect 10976 35254 10978 35306
rect 10978 35254 11030 35306
rect 11030 35254 11032 35306
rect 10976 35252 11032 35254
rect 11080 35306 11136 35308
rect 11080 35254 11082 35306
rect 11082 35254 11134 35306
rect 11134 35254 11136 35306
rect 11080 35252 11136 35254
rect 12236 35698 12292 35700
rect 12236 35646 12238 35698
rect 12238 35646 12290 35698
rect 12290 35646 12292 35698
rect 12236 35644 12292 35646
rect 12124 35196 12180 35252
rect 12012 35084 12068 35140
rect 11340 34914 11396 34916
rect 11340 34862 11342 34914
rect 11342 34862 11394 34914
rect 11394 34862 11396 34914
rect 11340 34860 11396 34862
rect 10444 34524 10500 34580
rect 11676 34188 11732 34244
rect 13692 36482 13748 36484
rect 13692 36430 13694 36482
rect 13694 36430 13746 36482
rect 13746 36430 13748 36482
rect 13692 36428 13748 36430
rect 12908 35698 12964 35700
rect 12908 35646 12910 35698
rect 12910 35646 12962 35698
rect 12962 35646 12964 35698
rect 12908 35644 12964 35646
rect 13244 34972 13300 35028
rect 13020 34860 13076 34916
rect 12908 34802 12964 34804
rect 12908 34750 12910 34802
rect 12910 34750 12962 34802
rect 12962 34750 12964 34802
rect 12908 34748 12964 34750
rect 10872 33738 10928 33740
rect 10872 33686 10874 33738
rect 10874 33686 10926 33738
rect 10926 33686 10928 33738
rect 10872 33684 10928 33686
rect 10976 33738 11032 33740
rect 10976 33686 10978 33738
rect 10978 33686 11030 33738
rect 11030 33686 11032 33738
rect 10976 33684 11032 33686
rect 11080 33738 11136 33740
rect 11080 33686 11082 33738
rect 11082 33686 11134 33738
rect 11134 33686 11136 33738
rect 11080 33684 11136 33686
rect 9660 33346 9716 33348
rect 9660 33294 9662 33346
rect 9662 33294 9714 33346
rect 9714 33294 9716 33346
rect 9660 33292 9716 33294
rect 10332 33346 10388 33348
rect 10332 33294 10334 33346
rect 10334 33294 10386 33346
rect 10386 33294 10388 33346
rect 10332 33292 10388 33294
rect 11452 33292 11508 33348
rect 9436 33122 9492 33124
rect 9436 33070 9438 33122
rect 9438 33070 9490 33122
rect 9490 33070 9492 33122
rect 9436 33068 9492 33070
rect 4956 31890 5012 31892
rect 4956 31838 4958 31890
rect 4958 31838 5010 31890
rect 5010 31838 5012 31890
rect 4956 31836 5012 31838
rect 5628 31836 5684 31892
rect 6188 31666 6244 31668
rect 6188 31614 6190 31666
rect 6190 31614 6242 31666
rect 6242 31614 6244 31666
rect 6188 31612 6244 31614
rect 6076 31554 6132 31556
rect 6076 31502 6078 31554
rect 6078 31502 6130 31554
rect 6130 31502 6132 31554
rect 6076 31500 6132 31502
rect 4732 31388 4788 31444
rect 6300 31388 6356 31444
rect 5964 31276 6020 31332
rect 2940 23660 2996 23716
rect 2492 22540 2548 22596
rect 2828 22540 2884 22596
rect 2716 21810 2772 21812
rect 2716 21758 2718 21810
rect 2718 21758 2770 21810
rect 2770 21758 2772 21810
rect 2716 21756 2772 21758
rect 2604 21698 2660 21700
rect 2604 21646 2606 21698
rect 2606 21646 2658 21698
rect 2658 21646 2660 21698
rect 2604 21644 2660 21646
rect 1820 20018 1876 20020
rect 1820 19966 1822 20018
rect 1822 19966 1874 20018
rect 1874 19966 1876 20018
rect 1820 19964 1876 19966
rect 1932 18732 1988 18788
rect 1932 18562 1988 18564
rect 1932 18510 1934 18562
rect 1934 18510 1986 18562
rect 1986 18510 1988 18562
rect 1932 18508 1988 18510
rect 2380 20018 2436 20020
rect 2380 19966 2382 20018
rect 2382 19966 2434 20018
rect 2434 19966 2436 20018
rect 2380 19964 2436 19966
rect 2380 18674 2436 18676
rect 2380 18622 2382 18674
rect 2382 18622 2434 18674
rect 2434 18622 2436 18674
rect 2380 18620 2436 18622
rect 2156 17388 2212 17444
rect 1932 13804 1988 13860
rect 3164 29932 3220 29988
rect 4172 29426 4228 29428
rect 4172 29374 4174 29426
rect 4174 29374 4226 29426
rect 4226 29374 4228 29426
rect 4172 29372 4228 29374
rect 4620 29538 4676 29540
rect 4620 29486 4622 29538
rect 4622 29486 4674 29538
rect 4674 29486 4676 29538
rect 4620 29484 4676 29486
rect 3612 28812 3668 28868
rect 3164 28530 3220 28532
rect 3164 28478 3166 28530
rect 3166 28478 3218 28530
rect 3218 28478 3220 28530
rect 3164 28476 3220 28478
rect 3612 28476 3668 28532
rect 3388 28364 3444 28420
rect 3164 27804 3220 27860
rect 4172 27804 4228 27860
rect 4284 27692 4340 27748
rect 4844 29372 4900 29428
rect 5404 29820 5460 29876
rect 4844 28418 4900 28420
rect 4844 28366 4846 28418
rect 4846 28366 4898 28418
rect 4898 28366 4900 28418
rect 4844 28364 4900 28366
rect 5068 28700 5124 28756
rect 6636 30044 6692 30100
rect 6972 30994 7028 30996
rect 6972 30942 6974 30994
rect 6974 30942 7026 30994
rect 7026 30942 7028 30994
rect 6972 30940 7028 30942
rect 8540 32396 8596 32452
rect 8204 31106 8260 31108
rect 8204 31054 8206 31106
rect 8206 31054 8258 31106
rect 8258 31054 8260 31106
rect 8204 31052 8260 31054
rect 6412 29596 6468 29652
rect 6860 30044 6916 30100
rect 6972 29484 7028 29540
rect 5628 28028 5684 28084
rect 5516 27858 5572 27860
rect 5516 27806 5518 27858
rect 5518 27806 5570 27858
rect 5570 27806 5572 27858
rect 5516 27804 5572 27806
rect 4620 27692 4676 27748
rect 4956 27692 5012 27748
rect 4508 27132 4564 27188
rect 3724 27074 3780 27076
rect 3724 27022 3726 27074
rect 3726 27022 3778 27074
rect 3778 27022 3780 27074
rect 3724 27020 3780 27022
rect 3164 26236 3220 26292
rect 3612 25900 3668 25956
rect 3276 25618 3332 25620
rect 3276 25566 3278 25618
rect 3278 25566 3330 25618
rect 3330 25566 3332 25618
rect 3276 25564 3332 25566
rect 3612 25564 3668 25620
rect 4396 27020 4452 27076
rect 6524 28364 6580 28420
rect 5740 27692 5796 27748
rect 5852 27186 5908 27188
rect 5852 27134 5854 27186
rect 5854 27134 5906 27186
rect 5906 27134 5908 27186
rect 5852 27132 5908 27134
rect 5740 27074 5796 27076
rect 5740 27022 5742 27074
rect 5742 27022 5794 27074
rect 5794 27022 5796 27074
rect 5740 27020 5796 27022
rect 6076 27074 6132 27076
rect 6076 27022 6078 27074
rect 6078 27022 6130 27074
rect 6130 27022 6132 27074
rect 6076 27020 6132 27022
rect 6636 27692 6692 27748
rect 5292 26290 5348 26292
rect 5292 26238 5294 26290
rect 5294 26238 5346 26290
rect 5346 26238 5348 26290
rect 5292 26236 5348 26238
rect 4620 25900 4676 25956
rect 5516 25564 5572 25620
rect 4396 24892 4452 24948
rect 3164 23772 3220 23828
rect 3612 23826 3668 23828
rect 3612 23774 3614 23826
rect 3614 23774 3666 23826
rect 3666 23774 3668 23826
rect 3612 23772 3668 23774
rect 3836 23714 3892 23716
rect 3836 23662 3838 23714
rect 3838 23662 3890 23714
rect 3890 23662 3892 23714
rect 3836 23660 3892 23662
rect 4396 23436 4452 23492
rect 4732 23436 4788 23492
rect 3388 23042 3444 23044
rect 3388 22990 3390 23042
rect 3390 22990 3442 23042
rect 3442 22990 3444 23042
rect 3388 22988 3444 22990
rect 3052 22482 3108 22484
rect 3052 22430 3054 22482
rect 3054 22430 3106 22482
rect 3106 22430 3108 22482
rect 3052 22428 3108 22430
rect 3388 22428 3444 22484
rect 3052 20860 3108 20916
rect 3164 20972 3220 21028
rect 3052 19068 3108 19124
rect 2716 18620 2772 18676
rect 2604 17388 2660 17444
rect 2492 16268 2548 16324
rect 4620 22930 4676 22932
rect 4620 22878 4622 22930
rect 4622 22878 4674 22930
rect 4674 22878 4676 22930
rect 4620 22876 4676 22878
rect 4508 22540 4564 22596
rect 3948 21644 4004 21700
rect 4732 21644 4788 21700
rect 3500 20076 3556 20132
rect 3164 18562 3220 18564
rect 3164 18510 3166 18562
rect 3166 18510 3218 18562
rect 3218 18510 3220 18562
rect 3164 18508 3220 18510
rect 3388 19964 3444 20020
rect 3052 16828 3108 16884
rect 2380 15260 2436 15316
rect 2716 14588 2772 14644
rect 2604 13746 2660 13748
rect 2604 13694 2606 13746
rect 2606 13694 2658 13746
rect 2658 13694 2660 13746
rect 2604 13692 2660 13694
rect 2380 13244 2436 13300
rect 2604 13356 2660 13412
rect 2044 11676 2100 11732
rect 1932 11340 1988 11396
rect 2604 10722 2660 10724
rect 2604 10670 2606 10722
rect 2606 10670 2658 10722
rect 2658 10670 2660 10722
rect 2604 10668 2660 10670
rect 1932 10332 1988 10388
rect 2828 13244 2884 13300
rect 3052 15314 3108 15316
rect 3052 15262 3054 15314
rect 3054 15262 3106 15314
rect 3106 15262 3108 15314
rect 3052 15260 3108 15262
rect 3724 20018 3780 20020
rect 3724 19966 3726 20018
rect 3726 19966 3778 20018
rect 3778 19966 3780 20018
rect 3724 19964 3780 19966
rect 3612 19906 3668 19908
rect 3612 19854 3614 19906
rect 3614 19854 3666 19906
rect 3666 19854 3668 19906
rect 3612 19852 3668 19854
rect 3612 19122 3668 19124
rect 3612 19070 3614 19122
rect 3614 19070 3666 19122
rect 3666 19070 3668 19122
rect 3612 19068 3668 19070
rect 3612 16882 3668 16884
rect 3612 16830 3614 16882
rect 3614 16830 3666 16882
rect 3666 16830 3668 16882
rect 3612 16828 3668 16830
rect 3612 15036 3668 15092
rect 4620 20130 4676 20132
rect 4620 20078 4622 20130
rect 4622 20078 4674 20130
rect 4674 20078 4676 20130
rect 4620 20076 4676 20078
rect 3948 19292 4004 19348
rect 3836 18674 3892 18676
rect 3836 18622 3838 18674
rect 3838 18622 3890 18674
rect 3890 18622 3892 18674
rect 3836 18620 3892 18622
rect 4620 19292 4676 19348
rect 3948 17890 4004 17892
rect 3948 17838 3950 17890
rect 3950 17838 4002 17890
rect 4002 17838 4004 17890
rect 3948 17836 4004 17838
rect 4060 17388 4116 17444
rect 5292 25116 5348 25172
rect 5068 23042 5124 23044
rect 5068 22990 5070 23042
rect 5070 22990 5122 23042
rect 5122 22990 5124 23042
rect 5068 22988 5124 22990
rect 5628 23436 5684 23492
rect 5292 21756 5348 21812
rect 5516 21810 5572 21812
rect 5516 21758 5518 21810
rect 5518 21758 5570 21810
rect 5570 21758 5572 21810
rect 5516 21756 5572 21758
rect 5404 21698 5460 21700
rect 5404 21646 5406 21698
rect 5406 21646 5458 21698
rect 5458 21646 5460 21698
rect 5404 21644 5460 21646
rect 5852 23324 5908 23380
rect 4844 20412 4900 20468
rect 4956 20690 5012 20692
rect 4956 20638 4958 20690
rect 4958 20638 5010 20690
rect 5010 20638 5012 20690
rect 4956 20636 5012 20638
rect 4844 19852 4900 19908
rect 5068 20018 5124 20020
rect 5068 19966 5070 20018
rect 5070 19966 5122 20018
rect 5122 19966 5124 20018
rect 5068 19964 5124 19966
rect 4956 19458 5012 19460
rect 4956 19406 4958 19458
rect 4958 19406 5010 19458
rect 5010 19406 5012 19458
rect 4956 19404 5012 19406
rect 4844 19180 4900 19236
rect 5404 18450 5460 18452
rect 5404 18398 5406 18450
rect 5406 18398 5458 18450
rect 5458 18398 5460 18450
rect 5404 18396 5460 18398
rect 4956 17836 5012 17892
rect 4956 17442 5012 17444
rect 4956 17390 4958 17442
rect 4958 17390 5010 17442
rect 5010 17390 5012 17442
rect 4956 17388 5012 17390
rect 4396 16828 4452 16884
rect 3836 16770 3892 16772
rect 3836 16718 3838 16770
rect 3838 16718 3890 16770
rect 3890 16718 3892 16770
rect 3836 16716 3892 16718
rect 4060 16156 4116 16212
rect 3948 15314 4004 15316
rect 3948 15262 3950 15314
rect 3950 15262 4002 15314
rect 4002 15262 4004 15314
rect 3948 15260 4004 15262
rect 3388 14252 3444 14308
rect 3612 14476 3668 14532
rect 3164 13916 3220 13972
rect 3724 14306 3780 14308
rect 3724 14254 3726 14306
rect 3726 14254 3778 14306
rect 3778 14254 3780 14306
rect 3724 14252 3780 14254
rect 3836 14140 3892 14196
rect 3948 14364 4004 14420
rect 3836 13916 3892 13972
rect 3388 13746 3444 13748
rect 3388 13694 3390 13746
rect 3390 13694 3442 13746
rect 3442 13694 3444 13746
rect 3388 13692 3444 13694
rect 3500 13580 3556 13636
rect 3164 11676 3220 11732
rect 2828 11452 2884 11508
rect 3276 11506 3332 11508
rect 3276 11454 3278 11506
rect 3278 11454 3330 11506
rect 3330 11454 3332 11506
rect 3276 11452 3332 11454
rect 2492 9772 2548 9828
rect 1932 9602 1988 9604
rect 1932 9550 1934 9602
rect 1934 9550 1986 9602
rect 1986 9550 1988 9602
rect 1932 9548 1988 9550
rect 1932 8930 1988 8932
rect 1932 8878 1934 8930
rect 1934 8878 1986 8930
rect 1986 8878 1988 8930
rect 1932 8876 1988 8878
rect 2156 8370 2212 8372
rect 2156 8318 2158 8370
rect 2158 8318 2210 8370
rect 2210 8318 2212 8370
rect 2156 8316 2212 8318
rect 1820 7868 1876 7924
rect 3164 8034 3220 8036
rect 3164 7982 3166 8034
rect 3166 7982 3218 8034
rect 3218 7982 3220 8034
rect 3164 7980 3220 7982
rect 2492 7868 2548 7924
rect 3500 10386 3556 10388
rect 3500 10334 3502 10386
rect 3502 10334 3554 10386
rect 3554 10334 3556 10386
rect 3500 10332 3556 10334
rect 4508 16770 4564 16772
rect 4508 16718 4510 16770
rect 4510 16718 4562 16770
rect 4562 16718 4564 16770
rect 4508 16716 4564 16718
rect 4172 12796 4228 12852
rect 5292 16882 5348 16884
rect 5292 16830 5294 16882
rect 5294 16830 5346 16882
rect 5346 16830 5348 16882
rect 5292 16828 5348 16830
rect 4844 16770 4900 16772
rect 4844 16718 4846 16770
rect 4846 16718 4898 16770
rect 4898 16718 4900 16770
rect 4844 16716 4900 16718
rect 5628 20412 5684 20468
rect 6412 23042 6468 23044
rect 6412 22990 6414 23042
rect 6414 22990 6466 23042
rect 6466 22990 6468 23042
rect 6412 22988 6468 22990
rect 6188 22482 6244 22484
rect 6188 22430 6190 22482
rect 6190 22430 6242 22482
rect 6242 22430 6244 22482
rect 6188 22428 6244 22430
rect 6860 26124 6916 26180
rect 7308 28642 7364 28644
rect 7308 28590 7310 28642
rect 7310 28590 7362 28642
rect 7362 28590 7364 28642
rect 7308 28588 7364 28590
rect 7756 28642 7812 28644
rect 7756 28590 7758 28642
rect 7758 28590 7810 28642
rect 7810 28590 7812 28642
rect 7756 28588 7812 28590
rect 7980 28588 8036 28644
rect 7084 27746 7140 27748
rect 7084 27694 7086 27746
rect 7086 27694 7138 27746
rect 7138 27694 7140 27746
rect 7084 27692 7140 27694
rect 7084 26850 7140 26852
rect 7084 26798 7086 26850
rect 7086 26798 7138 26850
rect 7138 26798 7140 26850
rect 7084 26796 7140 26798
rect 9884 32732 9940 32788
rect 8988 32396 9044 32452
rect 10108 32620 10164 32676
rect 8764 31724 8820 31780
rect 8652 31052 8708 31108
rect 8652 30380 8708 30436
rect 9324 31778 9380 31780
rect 9324 31726 9326 31778
rect 9326 31726 9378 31778
rect 9378 31726 9380 31778
rect 9324 31724 9380 31726
rect 8988 30882 9044 30884
rect 8988 30830 8990 30882
rect 8990 30830 9042 30882
rect 9042 30830 9044 30882
rect 8988 30828 9044 30830
rect 9436 30380 9492 30436
rect 10872 32170 10928 32172
rect 10872 32118 10874 32170
rect 10874 32118 10926 32170
rect 10926 32118 10928 32170
rect 10872 32116 10928 32118
rect 10976 32170 11032 32172
rect 10976 32118 10978 32170
rect 10978 32118 11030 32170
rect 11030 32118 11032 32170
rect 10976 32116 11032 32118
rect 11080 32170 11136 32172
rect 11080 32118 11082 32170
rect 11082 32118 11134 32170
rect 11134 32118 11136 32170
rect 11080 32116 11136 32118
rect 12012 33346 12068 33348
rect 12012 33294 12014 33346
rect 12014 33294 12066 33346
rect 12066 33294 12068 33346
rect 12012 33292 12068 33294
rect 12348 33068 12404 33124
rect 13580 34972 13636 35028
rect 15484 36482 15540 36484
rect 15484 36430 15486 36482
rect 15486 36430 15538 36482
rect 15538 36430 15540 36482
rect 15484 36428 15540 36430
rect 15596 36316 15652 36372
rect 14364 36204 14420 36260
rect 15036 35810 15092 35812
rect 15036 35758 15038 35810
rect 15038 35758 15090 35810
rect 15090 35758 15092 35810
rect 15036 35756 15092 35758
rect 16380 36258 16436 36260
rect 16380 36206 16382 36258
rect 16382 36206 16434 36258
rect 16434 36206 16436 36258
rect 16380 36204 16436 36206
rect 15596 35756 15652 35812
rect 15148 35586 15204 35588
rect 15148 35534 15150 35586
rect 15150 35534 15202 35586
rect 15202 35534 15204 35586
rect 15148 35532 15204 35534
rect 13692 34748 13748 34804
rect 13916 35196 13972 35252
rect 14140 35026 14196 35028
rect 14140 34974 14142 35026
rect 14142 34974 14194 35026
rect 14194 34974 14196 35026
rect 14140 34972 14196 34974
rect 15036 35196 15092 35252
rect 14924 34972 14980 35028
rect 14364 34914 14420 34916
rect 14364 34862 14366 34914
rect 14366 34862 14418 34914
rect 14418 34862 14420 34914
rect 14364 34860 14420 34862
rect 13468 34242 13524 34244
rect 13468 34190 13470 34242
rect 13470 34190 13522 34242
rect 13522 34190 13524 34242
rect 13468 34188 13524 34190
rect 13692 33628 13748 33684
rect 14700 34188 14756 34244
rect 14364 33906 14420 33908
rect 14364 33854 14366 33906
rect 14366 33854 14418 33906
rect 14418 33854 14420 33906
rect 14364 33852 14420 33854
rect 14812 33852 14868 33908
rect 14364 33628 14420 33684
rect 13804 33292 13860 33348
rect 13132 33180 13188 33236
rect 13692 33234 13748 33236
rect 13692 33182 13694 33234
rect 13694 33182 13746 33234
rect 13746 33182 13748 33234
rect 13692 33180 13748 33182
rect 10444 31724 10500 31780
rect 10332 30882 10388 30884
rect 10332 30830 10334 30882
rect 10334 30830 10386 30882
rect 10386 30830 10388 30882
rect 10332 30828 10388 30830
rect 10668 30492 10724 30548
rect 10872 30602 10928 30604
rect 10872 30550 10874 30602
rect 10874 30550 10926 30602
rect 10926 30550 10928 30602
rect 10872 30548 10928 30550
rect 10976 30602 11032 30604
rect 10976 30550 10978 30602
rect 10978 30550 11030 30602
rect 11030 30550 11032 30602
rect 10976 30548 11032 30550
rect 11080 30602 11136 30604
rect 11080 30550 11082 30602
rect 11082 30550 11134 30602
rect 11134 30550 11136 30602
rect 11080 30548 11136 30550
rect 9884 30380 9940 30436
rect 8876 30044 8932 30100
rect 9548 30098 9604 30100
rect 9548 30046 9550 30098
rect 9550 30046 9602 30098
rect 9602 30046 9604 30098
rect 9548 30044 9604 30046
rect 15260 34524 15316 34580
rect 15148 33628 15204 33684
rect 18844 37324 18900 37380
rect 16492 35756 16548 35812
rect 16604 36092 16660 36148
rect 16380 35698 16436 35700
rect 16380 35646 16382 35698
rect 16382 35646 16434 35698
rect 16434 35646 16436 35698
rect 16380 35644 16436 35646
rect 16044 35586 16100 35588
rect 16044 35534 16046 35586
rect 16046 35534 16098 35586
rect 16098 35534 16100 35586
rect 16044 35532 16100 35534
rect 16380 34914 16436 34916
rect 16380 34862 16382 34914
rect 16382 34862 16434 34914
rect 16434 34862 16436 34914
rect 16380 34860 16436 34862
rect 15820 34802 15876 34804
rect 15820 34750 15822 34802
rect 15822 34750 15874 34802
rect 15874 34750 15876 34802
rect 15820 34748 15876 34750
rect 15260 32620 15316 32676
rect 13020 32562 13076 32564
rect 13020 32510 13022 32562
rect 13022 32510 13074 32562
rect 13074 32510 13076 32562
rect 13020 32508 13076 32510
rect 14028 32562 14084 32564
rect 14028 32510 14030 32562
rect 14030 32510 14082 32562
rect 14082 32510 14084 32562
rect 14028 32508 14084 32510
rect 14252 32508 14308 32564
rect 13244 32396 13300 32452
rect 14140 32450 14196 32452
rect 14140 32398 14142 32450
rect 14142 32398 14194 32450
rect 14194 32398 14196 32450
rect 14140 32396 14196 32398
rect 12796 31164 12852 31220
rect 13468 31218 13524 31220
rect 13468 31166 13470 31218
rect 13470 31166 13522 31218
rect 13522 31166 13524 31218
rect 13468 31164 13524 31166
rect 11900 30380 11956 30436
rect 12460 30940 12516 30996
rect 10332 30268 10388 30324
rect 10668 30268 10724 30324
rect 10556 30210 10612 30212
rect 10556 30158 10558 30210
rect 10558 30158 10610 30210
rect 10610 30158 10612 30210
rect 10556 30156 10612 30158
rect 10444 30098 10500 30100
rect 10444 30046 10446 30098
rect 10446 30046 10498 30098
rect 10498 30046 10500 30098
rect 10444 30044 10500 30046
rect 11564 30322 11620 30324
rect 11564 30270 11566 30322
rect 11566 30270 11618 30322
rect 11618 30270 11620 30322
rect 11564 30268 11620 30270
rect 11788 30210 11844 30212
rect 11788 30158 11790 30210
rect 11790 30158 11842 30210
rect 11842 30158 11844 30210
rect 11788 30156 11844 30158
rect 14140 31778 14196 31780
rect 14140 31726 14142 31778
rect 14142 31726 14194 31778
rect 14194 31726 14196 31778
rect 14140 31724 14196 31726
rect 13804 30994 13860 30996
rect 13804 30942 13806 30994
rect 13806 30942 13858 30994
rect 13858 30942 13860 30994
rect 13804 30940 13860 30942
rect 13692 30380 13748 30436
rect 12908 29820 12964 29876
rect 11004 29596 11060 29652
rect 12124 29650 12180 29652
rect 12124 29598 12126 29650
rect 12126 29598 12178 29650
rect 12178 29598 12180 29650
rect 12124 29596 12180 29598
rect 11452 29426 11508 29428
rect 11452 29374 11454 29426
rect 11454 29374 11506 29426
rect 11506 29374 11508 29426
rect 11452 29372 11508 29374
rect 12348 29372 12404 29428
rect 11340 29314 11396 29316
rect 11340 29262 11342 29314
rect 11342 29262 11394 29314
rect 11394 29262 11396 29314
rect 11340 29260 11396 29262
rect 12124 29260 12180 29316
rect 10872 29034 10928 29036
rect 10872 28982 10874 29034
rect 10874 28982 10926 29034
rect 10926 28982 10928 29034
rect 10872 28980 10928 28982
rect 10976 29034 11032 29036
rect 10976 28982 10978 29034
rect 10978 28982 11030 29034
rect 11030 28982 11032 29034
rect 10976 28980 11032 28982
rect 11080 29034 11136 29036
rect 11080 28982 11082 29034
rect 11082 28982 11134 29034
rect 11134 28982 11136 29034
rect 11080 28980 11136 28982
rect 9884 28588 9940 28644
rect 8764 27244 8820 27300
rect 8316 26908 8372 26964
rect 8652 26962 8708 26964
rect 8652 26910 8654 26962
rect 8654 26910 8706 26962
rect 8706 26910 8708 26962
rect 8652 26908 8708 26910
rect 8204 26850 8260 26852
rect 8204 26798 8206 26850
rect 8206 26798 8258 26850
rect 8258 26798 8260 26850
rect 8204 26796 8260 26798
rect 7420 26402 7476 26404
rect 7420 26350 7422 26402
rect 7422 26350 7474 26402
rect 7474 26350 7476 26402
rect 7420 26348 7476 26350
rect 7084 26124 7140 26180
rect 7308 26124 7364 26180
rect 9212 27132 9268 27188
rect 9548 27186 9604 27188
rect 9548 27134 9550 27186
rect 9550 27134 9602 27186
rect 9602 27134 9604 27186
rect 9548 27132 9604 27134
rect 8876 26796 8932 26852
rect 9548 26684 9604 26740
rect 7980 26402 8036 26404
rect 7980 26350 7982 26402
rect 7982 26350 8034 26402
rect 8034 26350 8036 26402
rect 7980 26348 8036 26350
rect 8876 26402 8932 26404
rect 8876 26350 8878 26402
rect 8878 26350 8930 26402
rect 8930 26350 8932 26402
rect 8876 26348 8932 26350
rect 7644 25900 7700 25956
rect 7756 26236 7812 26292
rect 7420 25564 7476 25620
rect 8876 26012 8932 26068
rect 7084 24722 7140 24724
rect 7084 24670 7086 24722
rect 7086 24670 7138 24722
rect 7138 24670 7140 24722
rect 7084 24668 7140 24670
rect 7420 24332 7476 24388
rect 7644 24162 7700 24164
rect 7644 24110 7646 24162
rect 7646 24110 7698 24162
rect 7698 24110 7700 24162
rect 7644 24108 7700 24110
rect 8092 24108 8148 24164
rect 6972 23154 7028 23156
rect 6972 23102 6974 23154
rect 6974 23102 7026 23154
rect 7026 23102 7028 23154
rect 6972 23100 7028 23102
rect 7084 22988 7140 23044
rect 6748 22428 6804 22484
rect 6972 21698 7028 21700
rect 6972 21646 6974 21698
rect 6974 21646 7026 21698
rect 7026 21646 7028 21698
rect 6972 21644 7028 21646
rect 7196 21698 7252 21700
rect 7196 21646 7198 21698
rect 7198 21646 7250 21698
rect 7250 21646 7252 21698
rect 7196 21644 7252 21646
rect 6636 21586 6692 21588
rect 6636 21534 6638 21586
rect 6638 21534 6690 21586
rect 6690 21534 6692 21586
rect 6636 21532 6692 21534
rect 7868 23938 7924 23940
rect 7868 23886 7870 23938
rect 7870 23886 7922 23938
rect 7922 23886 7924 23938
rect 7868 23884 7924 23886
rect 8428 23884 8484 23940
rect 9660 26012 9716 26068
rect 9660 24722 9716 24724
rect 9660 24670 9662 24722
rect 9662 24670 9714 24722
rect 9714 24670 9716 24722
rect 9660 24668 9716 24670
rect 9212 23714 9268 23716
rect 9212 23662 9214 23714
rect 9214 23662 9266 23714
rect 9266 23662 9268 23714
rect 9212 23660 9268 23662
rect 8764 23548 8820 23604
rect 8204 23154 8260 23156
rect 8204 23102 8206 23154
rect 8206 23102 8258 23154
rect 8258 23102 8260 23154
rect 8204 23100 8260 23102
rect 7756 23042 7812 23044
rect 7756 22990 7758 23042
rect 7758 22990 7810 23042
rect 7810 22990 7812 23042
rect 7756 22988 7812 22990
rect 7644 21756 7700 21812
rect 8540 22482 8596 22484
rect 8540 22430 8542 22482
rect 8542 22430 8594 22482
rect 8594 22430 8596 22482
rect 8540 22428 8596 22430
rect 8092 22204 8148 22260
rect 8204 21698 8260 21700
rect 8204 21646 8206 21698
rect 8206 21646 8258 21698
rect 8258 21646 8260 21698
rect 8204 21644 8260 21646
rect 8540 21644 8596 21700
rect 7308 21586 7364 21588
rect 7308 21534 7310 21586
rect 7310 21534 7362 21586
rect 7362 21534 7364 21586
rect 7308 21532 7364 21534
rect 6524 20914 6580 20916
rect 6524 20862 6526 20914
rect 6526 20862 6578 20914
rect 6578 20862 6580 20914
rect 6524 20860 6580 20862
rect 7196 20802 7252 20804
rect 7196 20750 7198 20802
rect 7198 20750 7250 20802
rect 7250 20750 7252 20802
rect 7196 20748 7252 20750
rect 6076 20690 6132 20692
rect 6076 20638 6078 20690
rect 6078 20638 6130 20690
rect 6130 20638 6132 20690
rect 6076 20636 6132 20638
rect 5964 19404 6020 19460
rect 6076 19234 6132 19236
rect 6076 19182 6078 19234
rect 6078 19182 6130 19234
rect 6130 19182 6132 19234
rect 6076 19180 6132 19182
rect 5740 17836 5796 17892
rect 6524 18396 6580 18452
rect 6748 19740 6804 19796
rect 6972 17666 7028 17668
rect 6972 17614 6974 17666
rect 6974 17614 7026 17666
rect 7026 17614 7028 17666
rect 6972 17612 7028 17614
rect 6972 16716 7028 16772
rect 6188 16210 6244 16212
rect 6188 16158 6190 16210
rect 6190 16158 6242 16210
rect 6242 16158 6244 16210
rect 6188 16156 6244 16158
rect 6636 16098 6692 16100
rect 6636 16046 6638 16098
rect 6638 16046 6690 16098
rect 6690 16046 6692 16098
rect 6636 16044 6692 16046
rect 4844 15260 4900 15316
rect 4508 15202 4564 15204
rect 4508 15150 4510 15202
rect 4510 15150 4562 15202
rect 4562 15150 4564 15202
rect 4508 15148 4564 15150
rect 4620 14530 4676 14532
rect 4620 14478 4622 14530
rect 4622 14478 4674 14530
rect 4674 14478 4676 14530
rect 4620 14476 4676 14478
rect 5404 15314 5460 15316
rect 5404 15262 5406 15314
rect 5406 15262 5458 15314
rect 5458 15262 5460 15314
rect 5404 15260 5460 15262
rect 4956 15036 5012 15092
rect 4508 13970 4564 13972
rect 4508 13918 4510 13970
rect 4510 13918 4562 13970
rect 4562 13918 4564 13970
rect 4508 13916 4564 13918
rect 4844 13746 4900 13748
rect 4844 13694 4846 13746
rect 4846 13694 4898 13746
rect 4898 13694 4900 13746
rect 4844 13692 4900 13694
rect 4732 13580 4788 13636
rect 5628 15036 5684 15092
rect 5516 14476 5572 14532
rect 6076 14306 6132 14308
rect 6076 14254 6078 14306
rect 6078 14254 6130 14306
rect 6130 14254 6132 14306
rect 6076 14252 6132 14254
rect 5516 13692 5572 13748
rect 5292 13634 5348 13636
rect 5292 13582 5294 13634
rect 5294 13582 5346 13634
rect 5346 13582 5348 13634
rect 5292 13580 5348 13582
rect 4956 13468 5012 13524
rect 4620 13356 4676 13412
rect 4844 12850 4900 12852
rect 4844 12798 4846 12850
rect 4846 12798 4898 12850
rect 4898 12798 4900 12850
rect 4844 12796 4900 12798
rect 4396 11676 4452 11732
rect 4172 11394 4228 11396
rect 4172 11342 4174 11394
rect 4174 11342 4226 11394
rect 4226 11342 4228 11394
rect 4172 11340 4228 11342
rect 4956 12236 5012 12292
rect 4620 11170 4676 11172
rect 4620 11118 4622 11170
rect 4622 11118 4674 11170
rect 4674 11118 4676 11170
rect 4620 11116 4676 11118
rect 4396 10610 4452 10612
rect 4396 10558 4398 10610
rect 4398 10558 4450 10610
rect 4450 10558 4452 10610
rect 4396 10556 4452 10558
rect 4732 10108 4788 10164
rect 3276 7868 3332 7924
rect 4508 9602 4564 9604
rect 4508 9550 4510 9602
rect 4510 9550 4562 9602
rect 4562 9550 4564 9602
rect 4508 9548 4564 9550
rect 4956 9884 5012 9940
rect 6076 13580 6132 13636
rect 5516 9772 5572 9828
rect 5628 13468 5684 13524
rect 5852 12290 5908 12292
rect 5852 12238 5854 12290
rect 5854 12238 5906 12290
rect 5906 12238 5908 12290
rect 5852 12236 5908 12238
rect 6636 13692 6692 13748
rect 7084 14418 7140 14420
rect 7084 14366 7086 14418
rect 7086 14366 7138 14418
rect 7138 14366 7140 14418
rect 7084 14364 7140 14366
rect 7196 14306 7252 14308
rect 7196 14254 7198 14306
rect 7198 14254 7250 14306
rect 7250 14254 7252 14306
rect 7196 14252 7252 14254
rect 6636 13244 6692 13300
rect 6188 11900 6244 11956
rect 5740 11340 5796 11396
rect 5852 11452 5908 11508
rect 6076 10610 6132 10612
rect 6076 10558 6078 10610
rect 6078 10558 6130 10610
rect 6130 10558 6132 10610
rect 6076 10556 6132 10558
rect 5740 10332 5796 10388
rect 6412 9996 6468 10052
rect 5852 9602 5908 9604
rect 5852 9550 5854 9602
rect 5854 9550 5906 9602
rect 5906 9550 5908 9602
rect 5852 9548 5908 9550
rect 4508 9100 4564 9156
rect 5740 9154 5796 9156
rect 5740 9102 5742 9154
rect 5742 9102 5794 9154
rect 5794 9102 5796 9154
rect 5740 9100 5796 9102
rect 3836 8316 3892 8372
rect 4284 9042 4340 9044
rect 4284 8990 4286 9042
rect 4286 8990 4338 9042
rect 4338 8990 4340 9042
rect 4284 8988 4340 8990
rect 5516 9042 5572 9044
rect 5516 8990 5518 9042
rect 5518 8990 5570 9042
rect 5570 8990 5572 9042
rect 5516 8988 5572 8990
rect 4620 8258 4676 8260
rect 4620 8206 4622 8258
rect 4622 8206 4674 8258
rect 4674 8206 4676 8258
rect 4620 8204 4676 8206
rect 4956 8540 5012 8596
rect 5404 8652 5460 8708
rect 3724 7980 3780 8036
rect 2492 7532 2548 7588
rect 1932 6412 1988 6468
rect 2716 7586 2772 7588
rect 2716 7534 2718 7586
rect 2718 7534 2770 7586
rect 2770 7534 2772 7586
rect 2716 7532 2772 7534
rect 3612 7420 3668 7476
rect 3500 6300 3556 6356
rect 4732 7644 4788 7700
rect 4172 7532 4228 7588
rect 4508 7474 4564 7476
rect 4508 7422 4510 7474
rect 4510 7422 4562 7474
rect 4562 7422 4564 7474
rect 4508 7420 4564 7422
rect 4620 7362 4676 7364
rect 4620 7310 4622 7362
rect 4622 7310 4674 7362
rect 4674 7310 4676 7362
rect 4620 7308 4676 7310
rect 3724 6466 3780 6468
rect 3724 6414 3726 6466
rect 3726 6414 3778 6466
rect 3778 6414 3780 6466
rect 3724 6412 3780 6414
rect 5068 6412 5124 6468
rect 5852 8146 5908 8148
rect 5852 8094 5854 8146
rect 5854 8094 5906 8146
rect 5906 8094 5908 8146
rect 5852 8092 5908 8094
rect 6412 9602 6468 9604
rect 6412 9550 6414 9602
rect 6414 9550 6466 9602
rect 6466 9550 6468 9602
rect 6412 9548 6468 9550
rect 7644 20914 7700 20916
rect 7644 20862 7646 20914
rect 7646 20862 7698 20914
rect 7698 20862 7700 20914
rect 7644 20860 7700 20862
rect 8204 20802 8260 20804
rect 8204 20750 8206 20802
rect 8206 20750 8258 20802
rect 8258 20750 8260 20802
rect 8204 20748 8260 20750
rect 8316 20076 8372 20132
rect 8988 22652 9044 22708
rect 8876 21756 8932 21812
rect 8764 21532 8820 21588
rect 8764 20860 8820 20916
rect 10108 27298 10164 27300
rect 10108 27246 10110 27298
rect 10110 27246 10162 27298
rect 10162 27246 10164 27298
rect 10108 27244 10164 27246
rect 10332 28364 10388 28420
rect 9996 27020 10052 27076
rect 9996 26572 10052 26628
rect 10556 27804 10612 27860
rect 11004 27580 11060 27636
rect 10872 27466 10928 27468
rect 10872 27414 10874 27466
rect 10874 27414 10926 27466
rect 10926 27414 10928 27466
rect 10872 27412 10928 27414
rect 10976 27466 11032 27468
rect 10976 27414 10978 27466
rect 10978 27414 11030 27466
rect 11030 27414 11032 27466
rect 10976 27412 11032 27414
rect 11080 27466 11136 27468
rect 11080 27414 11082 27466
rect 11082 27414 11134 27466
rect 11134 27414 11136 27466
rect 11080 27412 11136 27414
rect 10668 26962 10724 26964
rect 10668 26910 10670 26962
rect 10670 26910 10722 26962
rect 10722 26910 10724 26962
rect 10668 26908 10724 26910
rect 11676 26962 11732 26964
rect 11676 26910 11678 26962
rect 11678 26910 11730 26962
rect 11730 26910 11732 26962
rect 11676 26908 11732 26910
rect 9884 25228 9940 25284
rect 9996 25116 10052 25172
rect 11564 26684 11620 26740
rect 12012 26684 12068 26740
rect 12012 26402 12068 26404
rect 12012 26350 12014 26402
rect 12014 26350 12066 26402
rect 12066 26350 12068 26402
rect 12012 26348 12068 26350
rect 11004 26290 11060 26292
rect 11004 26238 11006 26290
rect 11006 26238 11058 26290
rect 11058 26238 11060 26290
rect 11004 26236 11060 26238
rect 10872 25898 10928 25900
rect 10872 25846 10874 25898
rect 10874 25846 10926 25898
rect 10926 25846 10928 25898
rect 10872 25844 10928 25846
rect 10976 25898 11032 25900
rect 10976 25846 10978 25898
rect 10978 25846 11030 25898
rect 11030 25846 11032 25898
rect 10976 25844 11032 25846
rect 11080 25898 11136 25900
rect 11080 25846 11082 25898
rect 11082 25846 11134 25898
rect 11134 25846 11136 25898
rect 11080 25844 11136 25846
rect 10780 25004 10836 25060
rect 10108 24162 10164 24164
rect 10108 24110 10110 24162
rect 10110 24110 10162 24162
rect 10162 24110 10164 24162
rect 10108 24108 10164 24110
rect 11676 26236 11732 26292
rect 12460 29260 12516 29316
rect 12908 29314 12964 29316
rect 12908 29262 12910 29314
rect 12910 29262 12962 29314
rect 12962 29262 12964 29314
rect 12908 29260 12964 29262
rect 12572 28364 12628 28420
rect 13244 28476 13300 28532
rect 13356 28364 13412 28420
rect 14812 31724 14868 31780
rect 13916 29820 13972 29876
rect 13804 28530 13860 28532
rect 13804 28478 13806 28530
rect 13806 28478 13858 28530
rect 13858 28478 13860 28530
rect 13804 28476 13860 28478
rect 14364 31276 14420 31332
rect 14700 31218 14756 31220
rect 14700 31166 14702 31218
rect 14702 31166 14754 31218
rect 14754 31166 14756 31218
rect 14700 31164 14756 31166
rect 15708 31666 15764 31668
rect 15708 31614 15710 31666
rect 15710 31614 15762 31666
rect 15762 31614 15764 31666
rect 15708 31612 15764 31614
rect 14924 31276 14980 31332
rect 15596 31164 15652 31220
rect 14924 30940 14980 30996
rect 14812 29820 14868 29876
rect 12124 25452 12180 25508
rect 12348 27692 12404 27748
rect 11900 25116 11956 25172
rect 12124 25004 12180 25060
rect 11228 24668 11284 24724
rect 11564 24556 11620 24612
rect 10872 24330 10928 24332
rect 10872 24278 10874 24330
rect 10874 24278 10926 24330
rect 10926 24278 10928 24330
rect 10872 24276 10928 24278
rect 10976 24330 11032 24332
rect 10976 24278 10978 24330
rect 10978 24278 11030 24330
rect 11030 24278 11032 24330
rect 10976 24276 11032 24278
rect 11080 24330 11136 24332
rect 11080 24278 11082 24330
rect 11082 24278 11134 24330
rect 11134 24278 11136 24330
rect 11080 24276 11136 24278
rect 11004 23884 11060 23940
rect 10556 23772 10612 23828
rect 9996 23660 10052 23716
rect 9660 23548 9716 23604
rect 9324 22876 9380 22932
rect 9772 22652 9828 22708
rect 9436 22482 9492 22484
rect 9436 22430 9438 22482
rect 9438 22430 9490 22482
rect 9490 22430 9492 22482
rect 9436 22428 9492 22430
rect 9772 22428 9828 22484
rect 9324 21868 9380 21924
rect 9436 22204 9492 22260
rect 9212 20690 9268 20692
rect 9212 20638 9214 20690
rect 9214 20638 9266 20690
rect 9266 20638 9268 20690
rect 9212 20636 9268 20638
rect 9324 20860 9380 20916
rect 8540 19404 8596 19460
rect 8316 18732 8372 18788
rect 8876 19234 8932 19236
rect 8876 19182 8878 19234
rect 8878 19182 8930 19234
rect 8930 19182 8932 19234
rect 8876 19180 8932 19182
rect 7868 18338 7924 18340
rect 7868 18286 7870 18338
rect 7870 18286 7922 18338
rect 7922 18286 7924 18338
rect 7868 18284 7924 18286
rect 8876 18674 8932 18676
rect 8876 18622 8878 18674
rect 8878 18622 8930 18674
rect 8930 18622 8932 18674
rect 8876 18620 8932 18622
rect 10108 23100 10164 23156
rect 9996 22204 10052 22260
rect 9884 21756 9940 21812
rect 9884 21474 9940 21476
rect 9884 21422 9886 21474
rect 9886 21422 9938 21474
rect 9938 21422 9940 21474
rect 9884 21420 9940 21422
rect 11116 23548 11172 23604
rect 11228 23884 11284 23940
rect 10872 22762 10928 22764
rect 10872 22710 10874 22762
rect 10874 22710 10926 22762
rect 10926 22710 10928 22762
rect 10872 22708 10928 22710
rect 10976 22762 11032 22764
rect 10976 22710 10978 22762
rect 10978 22710 11030 22762
rect 11030 22710 11032 22762
rect 10976 22708 11032 22710
rect 11080 22762 11136 22764
rect 11080 22710 11082 22762
rect 11082 22710 11134 22762
rect 11134 22710 11136 22762
rect 11080 22708 11136 22710
rect 10872 21194 10928 21196
rect 10872 21142 10874 21194
rect 10874 21142 10926 21194
rect 10926 21142 10928 21194
rect 10872 21140 10928 21142
rect 10976 21194 11032 21196
rect 10976 21142 10978 21194
rect 10978 21142 11030 21194
rect 11030 21142 11032 21194
rect 10976 21140 11032 21142
rect 11080 21194 11136 21196
rect 11080 21142 11082 21194
rect 11082 21142 11134 21194
rect 11134 21142 11136 21194
rect 11080 21140 11136 21142
rect 10668 20802 10724 20804
rect 10668 20750 10670 20802
rect 10670 20750 10722 20802
rect 10722 20750 10724 20802
rect 10668 20748 10724 20750
rect 9884 20690 9940 20692
rect 9884 20638 9886 20690
rect 9886 20638 9938 20690
rect 9938 20638 9940 20690
rect 9884 20636 9940 20638
rect 10556 20690 10612 20692
rect 10556 20638 10558 20690
rect 10558 20638 10610 20690
rect 10610 20638 10612 20690
rect 10780 20972 10836 21028
rect 10556 20636 10612 20638
rect 9436 19458 9492 19460
rect 9436 19406 9438 19458
rect 9438 19406 9490 19458
rect 9490 19406 9492 19458
rect 9436 19404 9492 19406
rect 9660 19234 9716 19236
rect 9660 19182 9662 19234
rect 9662 19182 9714 19234
rect 9714 19182 9716 19234
rect 9660 19180 9716 19182
rect 9884 19404 9940 19460
rect 11340 23772 11396 23828
rect 12012 24834 12068 24836
rect 12012 24782 12014 24834
rect 12014 24782 12066 24834
rect 12066 24782 12068 24834
rect 12012 24780 12068 24782
rect 12012 24556 12068 24612
rect 11788 24050 11844 24052
rect 11788 23998 11790 24050
rect 11790 23998 11842 24050
rect 11842 23998 11844 24050
rect 11788 23996 11844 23998
rect 11676 23772 11732 23828
rect 11676 22540 11732 22596
rect 11564 20802 11620 20804
rect 11564 20750 11566 20802
rect 11566 20750 11618 20802
rect 11618 20750 11620 20802
rect 11564 20748 11620 20750
rect 11116 20636 11172 20692
rect 10780 20412 10836 20468
rect 10108 20130 10164 20132
rect 10108 20078 10110 20130
rect 10110 20078 10162 20130
rect 10162 20078 10164 20130
rect 10108 20076 10164 20078
rect 9884 18674 9940 18676
rect 9884 18622 9886 18674
rect 9886 18622 9938 18674
rect 9938 18622 9940 18674
rect 9884 18620 9940 18622
rect 8764 17836 8820 17892
rect 8988 18284 9044 18340
rect 7980 17778 8036 17780
rect 7980 17726 7982 17778
rect 7982 17726 8034 17778
rect 8034 17726 8036 17778
rect 7980 17724 8036 17726
rect 7420 16156 7476 16212
rect 7756 16044 7812 16100
rect 7756 13634 7812 13636
rect 7756 13582 7758 13634
rect 7758 13582 7810 13634
rect 7810 13582 7812 13634
rect 7756 13580 7812 13582
rect 8428 17724 8484 17780
rect 8876 17666 8932 17668
rect 8876 17614 8878 17666
rect 8878 17614 8930 17666
rect 8930 17614 8932 17666
rect 8876 17612 8932 17614
rect 8540 17554 8596 17556
rect 8540 17502 8542 17554
rect 8542 17502 8594 17554
rect 8594 17502 8596 17554
rect 8540 17500 8596 17502
rect 9548 18396 9604 18452
rect 9772 18172 9828 18228
rect 10108 18284 10164 18340
rect 9660 17836 9716 17892
rect 10220 18396 10276 18452
rect 10556 18620 10612 18676
rect 10444 18172 10500 18228
rect 10220 17612 10276 17668
rect 8988 15820 9044 15876
rect 9212 15932 9268 15988
rect 7980 15148 8036 15204
rect 8540 15148 8596 15204
rect 9996 15986 10052 15988
rect 9996 15934 9998 15986
rect 9998 15934 10050 15986
rect 10050 15934 10052 15986
rect 9996 15932 10052 15934
rect 9884 15874 9940 15876
rect 9884 15822 9886 15874
rect 9886 15822 9938 15874
rect 9938 15822 9940 15874
rect 9884 15820 9940 15822
rect 10444 15874 10500 15876
rect 10444 15822 10446 15874
rect 10446 15822 10498 15874
rect 10498 15822 10500 15874
rect 10444 15820 10500 15822
rect 9660 15372 9716 15428
rect 9660 15202 9716 15204
rect 9660 15150 9662 15202
rect 9662 15150 9714 15202
rect 9714 15150 9716 15202
rect 9660 15148 9716 15150
rect 8092 14364 8148 14420
rect 8764 14530 8820 14532
rect 8764 14478 8766 14530
rect 8766 14478 8818 14530
rect 8818 14478 8820 14530
rect 8764 14476 8820 14478
rect 8652 14364 8708 14420
rect 8204 13746 8260 13748
rect 8204 13694 8206 13746
rect 8206 13694 8258 13746
rect 8258 13694 8260 13746
rect 8204 13692 8260 13694
rect 7868 13132 7924 13188
rect 9436 14700 9492 14756
rect 9324 14418 9380 14420
rect 9324 14366 9326 14418
rect 9326 14366 9378 14418
rect 9378 14366 9380 14418
rect 9324 14364 9380 14366
rect 9548 14306 9604 14308
rect 9548 14254 9550 14306
rect 9550 14254 9602 14306
rect 9602 14254 9604 14306
rect 9548 14252 9604 14254
rect 9884 14252 9940 14308
rect 9884 13692 9940 13748
rect 9772 13580 9828 13636
rect 10444 13804 10500 13860
rect 10220 13580 10276 13636
rect 7196 12684 7252 12740
rect 7756 12738 7812 12740
rect 7756 12686 7758 12738
rect 7758 12686 7810 12738
rect 7810 12686 7812 12738
rect 7756 12684 7812 12686
rect 6860 9548 6916 9604
rect 6524 9100 6580 9156
rect 5964 7868 6020 7924
rect 6188 7868 6244 7924
rect 6748 9042 6804 9044
rect 6748 8990 6750 9042
rect 6750 8990 6802 9042
rect 6802 8990 6804 9042
rect 6748 8988 6804 8990
rect 6412 7586 6468 7588
rect 6412 7534 6414 7586
rect 6414 7534 6466 7586
rect 6466 7534 6468 7586
rect 6412 7532 6468 7534
rect 5740 7474 5796 7476
rect 5740 7422 5742 7474
rect 5742 7422 5794 7474
rect 5794 7422 5796 7474
rect 5740 7420 5796 7422
rect 4508 6300 4564 6356
rect 4732 6300 4788 6356
rect 1596 4396 1652 4452
rect 3836 5122 3892 5124
rect 3836 5070 3838 5122
rect 3838 5070 3890 5122
rect 3890 5070 3892 5122
rect 3836 5068 3892 5070
rect 4844 5122 4900 5124
rect 4844 5070 4846 5122
rect 4846 5070 4898 5122
rect 4898 5070 4900 5122
rect 4844 5068 4900 5070
rect 2940 4508 2996 4564
rect 3052 4844 3108 4900
rect 3612 4898 3668 4900
rect 3612 4846 3614 4898
rect 3614 4846 3666 4898
rect 3666 4846 3668 4898
rect 3612 4844 3668 4846
rect 6076 6300 6132 6356
rect 5628 5964 5684 6020
rect 5404 5906 5460 5908
rect 5404 5854 5406 5906
rect 5406 5854 5458 5906
rect 5458 5854 5460 5906
rect 5404 5852 5460 5854
rect 5068 4732 5124 4788
rect 3612 4562 3668 4564
rect 3612 4510 3614 4562
rect 3614 4510 3666 4562
rect 3666 4510 3668 4562
rect 3612 4508 3668 4510
rect 3948 4450 4004 4452
rect 3948 4398 3950 4450
rect 3950 4398 4002 4450
rect 4002 4398 4004 4450
rect 3948 4396 4004 4398
rect 4508 4450 4564 4452
rect 4508 4398 4510 4450
rect 4510 4398 4562 4450
rect 4562 4398 4564 4450
rect 4508 4396 4564 4398
rect 1932 3948 1988 4004
rect 4956 3666 5012 3668
rect 4956 3614 4958 3666
rect 4958 3614 5010 3666
rect 5010 3614 5012 3666
rect 4956 3612 5012 3614
rect 2156 3554 2212 3556
rect 2156 3502 2158 3554
rect 2158 3502 2210 3554
rect 2210 3502 2212 3554
rect 2156 3500 2212 3502
rect 2716 3500 2772 3556
rect 1820 1484 1876 1540
rect 5628 3554 5684 3556
rect 5628 3502 5630 3554
rect 5630 3502 5682 3554
rect 5682 3502 5684 3554
rect 5628 3500 5684 3502
rect 2828 3442 2884 3444
rect 2828 3390 2830 3442
rect 2830 3390 2882 3442
rect 2882 3390 2884 3442
rect 2828 3388 2884 3390
rect 6748 5964 6804 6020
rect 6636 5292 6692 5348
rect 7084 9772 7140 9828
rect 7084 8988 7140 9044
rect 8540 12684 8596 12740
rect 8876 12460 8932 12516
rect 8092 12236 8148 12292
rect 7532 11900 7588 11956
rect 7420 10108 7476 10164
rect 7196 9212 7252 9268
rect 7196 8370 7252 8372
rect 7196 8318 7198 8370
rect 7198 8318 7250 8370
rect 7250 8318 7252 8370
rect 7196 8316 7252 8318
rect 7420 6018 7476 6020
rect 7420 5966 7422 6018
rect 7422 5966 7474 6018
rect 7474 5966 7476 6018
rect 7420 5964 7476 5966
rect 6860 4396 6916 4452
rect 7196 3500 7252 3556
rect 6748 3442 6804 3444
rect 6748 3390 6750 3442
rect 6750 3390 6802 3442
rect 6802 3390 6804 3442
rect 6748 3388 6804 3390
rect 6972 3388 7028 3444
rect 6524 2828 6580 2884
rect 7868 10722 7924 10724
rect 7868 10670 7870 10722
rect 7870 10670 7922 10722
rect 7922 10670 7924 10722
rect 7868 10668 7924 10670
rect 7980 10556 8036 10612
rect 7644 10050 7700 10052
rect 7644 9998 7646 10050
rect 7646 9998 7698 10050
rect 7698 9998 7700 10050
rect 7644 9996 7700 9998
rect 7868 9938 7924 9940
rect 7868 9886 7870 9938
rect 7870 9886 7922 9938
rect 7922 9886 7924 9938
rect 7868 9884 7924 9886
rect 7980 9772 8036 9828
rect 8876 11676 8932 11732
rect 8764 11394 8820 11396
rect 8764 11342 8766 11394
rect 8766 11342 8818 11394
rect 8818 11342 8820 11394
rect 8764 11340 8820 11342
rect 8988 12178 9044 12180
rect 8988 12126 8990 12178
rect 8990 12126 9042 12178
rect 9042 12126 9044 12178
rect 8988 12124 9044 12126
rect 9884 12012 9940 12068
rect 8876 11116 8932 11172
rect 8652 10722 8708 10724
rect 8652 10670 8654 10722
rect 8654 10670 8706 10722
rect 8706 10670 8708 10722
rect 8652 10668 8708 10670
rect 8652 10108 8708 10164
rect 8204 9938 8260 9940
rect 8204 9886 8206 9938
rect 8206 9886 8258 9938
rect 8258 9886 8260 9938
rect 8204 9884 8260 9886
rect 8204 8428 8260 8484
rect 7756 8370 7812 8372
rect 7756 8318 7758 8370
rect 7758 8318 7810 8370
rect 7810 8318 7812 8370
rect 7756 8316 7812 8318
rect 7868 8204 7924 8260
rect 8988 10108 9044 10164
rect 8876 9826 8932 9828
rect 8876 9774 8878 9826
rect 8878 9774 8930 9826
rect 8930 9774 8932 9826
rect 8876 9772 8932 9774
rect 8876 9266 8932 9268
rect 8876 9214 8878 9266
rect 8878 9214 8930 9266
rect 8930 9214 8932 9266
rect 8876 9212 8932 9214
rect 8316 8204 8372 8260
rect 8204 8034 8260 8036
rect 8204 7982 8206 8034
rect 8206 7982 8258 8034
rect 8258 7982 8260 8034
rect 8204 7980 8260 7982
rect 8540 8988 8596 9044
rect 7644 5234 7700 5236
rect 7644 5182 7646 5234
rect 7646 5182 7698 5234
rect 7698 5182 7700 5234
rect 7644 5180 7700 5182
rect 9772 9212 9828 9268
rect 8652 8316 8708 8372
rect 8876 8316 8932 8372
rect 10108 12124 10164 12180
rect 9996 11676 10052 11732
rect 10872 19626 10928 19628
rect 10872 19574 10874 19626
rect 10874 19574 10926 19626
rect 10926 19574 10928 19626
rect 10872 19572 10928 19574
rect 10976 19626 11032 19628
rect 10976 19574 10978 19626
rect 10978 19574 11030 19626
rect 11030 19574 11032 19626
rect 10976 19572 11032 19574
rect 11080 19626 11136 19628
rect 11080 19574 11082 19626
rect 11082 19574 11134 19626
rect 11134 19574 11136 19626
rect 11080 19572 11136 19574
rect 11452 18508 11508 18564
rect 11340 18338 11396 18340
rect 11340 18286 11342 18338
rect 11342 18286 11394 18338
rect 11394 18286 11396 18338
rect 11340 18284 11396 18286
rect 10872 18058 10928 18060
rect 10872 18006 10874 18058
rect 10874 18006 10926 18058
rect 10926 18006 10928 18058
rect 10872 18004 10928 18006
rect 10976 18058 11032 18060
rect 10976 18006 10978 18058
rect 10978 18006 11030 18058
rect 11030 18006 11032 18058
rect 10976 18004 11032 18006
rect 11080 18058 11136 18060
rect 11080 18006 11082 18058
rect 11082 18006 11134 18058
rect 11134 18006 11136 18058
rect 11080 18004 11136 18006
rect 10872 16490 10928 16492
rect 10872 16438 10874 16490
rect 10874 16438 10926 16490
rect 10926 16438 10928 16490
rect 10872 16436 10928 16438
rect 10976 16490 11032 16492
rect 10976 16438 10978 16490
rect 10978 16438 11030 16490
rect 11030 16438 11032 16490
rect 10976 16436 11032 16438
rect 11080 16490 11136 16492
rect 11080 16438 11082 16490
rect 11082 16438 11134 16490
rect 11134 16438 11136 16490
rect 11080 16436 11136 16438
rect 11564 18396 11620 18452
rect 11676 17836 11732 17892
rect 11788 17554 11844 17556
rect 11788 17502 11790 17554
rect 11790 17502 11842 17554
rect 11842 17502 11844 17554
rect 11788 17500 11844 17502
rect 12124 23996 12180 24052
rect 12236 24220 12292 24276
rect 12124 22540 12180 22596
rect 13244 27692 13300 27748
rect 12908 26908 12964 26964
rect 12796 26796 12852 26852
rect 12908 26514 12964 26516
rect 12908 26462 12910 26514
rect 12910 26462 12962 26514
rect 12962 26462 12964 26514
rect 12908 26460 12964 26462
rect 12460 26348 12516 26404
rect 12460 26178 12516 26180
rect 12460 26126 12462 26178
rect 12462 26126 12514 26178
rect 12514 26126 12516 26178
rect 12460 26124 12516 26126
rect 12572 25116 12628 25172
rect 12908 25116 12964 25172
rect 12460 24892 12516 24948
rect 13580 27858 13636 27860
rect 13580 27806 13582 27858
rect 13582 27806 13634 27858
rect 13634 27806 13636 27858
rect 13580 27804 13636 27806
rect 13692 26962 13748 26964
rect 13692 26910 13694 26962
rect 13694 26910 13746 26962
rect 13746 26910 13748 26962
rect 13692 26908 13748 26910
rect 14028 28140 14084 28196
rect 14588 28140 14644 28196
rect 15484 29932 15540 29988
rect 16156 31612 16212 31668
rect 17276 35644 17332 35700
rect 17948 36316 18004 36372
rect 17836 35810 17892 35812
rect 17836 35758 17838 35810
rect 17838 35758 17890 35810
rect 17890 35758 17892 35810
rect 17836 35756 17892 35758
rect 18060 35644 18116 35700
rect 18508 36316 18564 36372
rect 17724 34972 17780 35028
rect 16828 34300 16884 34356
rect 16940 34242 16996 34244
rect 16940 34190 16942 34242
rect 16942 34190 16994 34242
rect 16994 34190 16996 34242
rect 16940 34188 16996 34190
rect 18172 34690 18228 34692
rect 18172 34638 18174 34690
rect 18174 34638 18226 34690
rect 18226 34638 18228 34690
rect 18172 34636 18228 34638
rect 17836 34354 17892 34356
rect 17836 34302 17838 34354
rect 17838 34302 17890 34354
rect 17890 34302 17892 34354
rect 17836 34300 17892 34302
rect 21868 36540 21924 36596
rect 18844 36204 18900 36260
rect 19628 35644 19684 35700
rect 18732 35084 18788 35140
rect 19964 35698 20020 35700
rect 19964 35646 19966 35698
rect 19966 35646 20018 35698
rect 20018 35646 20020 35698
rect 19964 35644 20020 35646
rect 19740 35138 19796 35140
rect 19740 35086 19742 35138
rect 19742 35086 19794 35138
rect 19794 35086 19796 35138
rect 19740 35084 19796 35086
rect 20076 35138 20132 35140
rect 20076 35086 20078 35138
rect 20078 35086 20130 35138
rect 20130 35086 20132 35138
rect 20076 35084 20132 35086
rect 20532 36090 20588 36092
rect 20532 36038 20534 36090
rect 20534 36038 20586 36090
rect 20586 36038 20588 36090
rect 20532 36036 20588 36038
rect 20636 36090 20692 36092
rect 20636 36038 20638 36090
rect 20638 36038 20690 36090
rect 20690 36038 20692 36090
rect 20636 36036 20692 36038
rect 20740 36090 20796 36092
rect 20740 36038 20742 36090
rect 20742 36038 20794 36090
rect 20794 36038 20796 36090
rect 20740 36036 20796 36038
rect 21532 35196 21588 35252
rect 20412 34972 20468 35028
rect 22764 36540 22820 36596
rect 24892 37772 24948 37828
rect 24892 36540 24948 36596
rect 24556 36482 24612 36484
rect 24556 36430 24558 36482
rect 24558 36430 24610 36482
rect 24610 36430 24612 36482
rect 24556 36428 24612 36430
rect 23884 36316 23940 36372
rect 23212 35868 23268 35924
rect 19740 34860 19796 34916
rect 20524 34914 20580 34916
rect 20524 34862 20526 34914
rect 20526 34862 20578 34914
rect 20578 34862 20580 34914
rect 20524 34860 20580 34862
rect 18620 34802 18676 34804
rect 18620 34750 18622 34802
rect 18622 34750 18674 34802
rect 18674 34750 18676 34802
rect 18620 34748 18676 34750
rect 20532 34522 20588 34524
rect 20532 34470 20534 34522
rect 20534 34470 20586 34522
rect 20586 34470 20588 34522
rect 20532 34468 20588 34470
rect 20636 34522 20692 34524
rect 20636 34470 20638 34522
rect 20638 34470 20690 34522
rect 20690 34470 20692 34522
rect 20636 34468 20692 34470
rect 20740 34522 20796 34524
rect 20740 34470 20742 34522
rect 20742 34470 20794 34522
rect 20794 34470 20796 34522
rect 20740 34468 20796 34470
rect 18172 33852 18228 33908
rect 17948 33740 18004 33796
rect 17276 33628 17332 33684
rect 17612 33628 17668 33684
rect 16604 31164 16660 31220
rect 21196 34188 21252 34244
rect 22428 35698 22484 35700
rect 22428 35646 22430 35698
rect 22430 35646 22482 35698
rect 22482 35646 22484 35698
rect 22428 35644 22484 35646
rect 22988 35532 23044 35588
rect 22652 35196 22708 35252
rect 23100 35084 23156 35140
rect 20188 33852 20244 33908
rect 21980 33852 22036 33908
rect 20188 33628 20244 33684
rect 22988 33852 23044 33908
rect 22764 33628 22820 33684
rect 19964 33122 20020 33124
rect 19964 33070 19966 33122
rect 19966 33070 20018 33122
rect 20018 33070 20020 33122
rect 19964 33068 20020 33070
rect 19068 32562 19124 32564
rect 19068 32510 19070 32562
rect 19070 32510 19122 32562
rect 19122 32510 19124 32562
rect 19068 32508 19124 32510
rect 17052 31276 17108 31332
rect 20532 32954 20588 32956
rect 20532 32902 20534 32954
rect 20534 32902 20586 32954
rect 20586 32902 20588 32954
rect 20532 32900 20588 32902
rect 20636 32954 20692 32956
rect 20636 32902 20638 32954
rect 20638 32902 20690 32954
rect 20690 32902 20692 32954
rect 20636 32900 20692 32902
rect 20740 32954 20796 32956
rect 20740 32902 20742 32954
rect 20742 32902 20794 32954
rect 20794 32902 20796 32954
rect 20740 32900 20796 32902
rect 22652 32674 22708 32676
rect 22652 32622 22654 32674
rect 22654 32622 22706 32674
rect 22706 32622 22708 32674
rect 22652 32620 22708 32622
rect 20300 32508 20356 32564
rect 20188 31388 20244 31444
rect 20636 31778 20692 31780
rect 20636 31726 20638 31778
rect 20638 31726 20690 31778
rect 20690 31726 20692 31778
rect 20636 31724 20692 31726
rect 21756 31778 21812 31780
rect 21756 31726 21758 31778
rect 21758 31726 21810 31778
rect 21810 31726 21812 31778
rect 21756 31724 21812 31726
rect 20860 31612 20916 31668
rect 20532 31386 20588 31388
rect 20532 31334 20534 31386
rect 20534 31334 20586 31386
rect 20586 31334 20588 31386
rect 20532 31332 20588 31334
rect 20636 31386 20692 31388
rect 20636 31334 20638 31386
rect 20638 31334 20690 31386
rect 20690 31334 20692 31386
rect 20636 31332 20692 31334
rect 20740 31386 20796 31388
rect 20740 31334 20742 31386
rect 20742 31334 20794 31386
rect 20794 31334 20796 31386
rect 20740 31332 20796 31334
rect 16716 30882 16772 30884
rect 16716 30830 16718 30882
rect 16718 30830 16770 30882
rect 16770 30830 16772 30882
rect 16716 30828 16772 30830
rect 17612 30882 17668 30884
rect 17612 30830 17614 30882
rect 17614 30830 17666 30882
rect 17666 30830 17668 30882
rect 17612 30828 17668 30830
rect 18732 30994 18788 30996
rect 18732 30942 18734 30994
rect 18734 30942 18786 30994
rect 18786 30942 18788 30994
rect 18732 30940 18788 30942
rect 19180 30604 19236 30660
rect 17612 30380 17668 30436
rect 18732 30380 18788 30436
rect 16044 29596 16100 29652
rect 16380 29650 16436 29652
rect 16380 29598 16382 29650
rect 16382 29598 16434 29650
rect 16434 29598 16436 29650
rect 16380 29596 16436 29598
rect 17164 29596 17220 29652
rect 15372 29036 15428 29092
rect 15484 28924 15540 28980
rect 15372 28642 15428 28644
rect 15372 28590 15374 28642
rect 15374 28590 15426 28642
rect 15426 28590 15428 28642
rect 15372 28588 15428 28590
rect 14924 27970 14980 27972
rect 14924 27918 14926 27970
rect 14926 27918 14978 27970
rect 14978 27918 14980 27970
rect 14924 27916 14980 27918
rect 14140 27804 14196 27860
rect 14028 27580 14084 27636
rect 14252 27244 14308 27300
rect 13804 26572 13860 26628
rect 13580 26514 13636 26516
rect 13580 26462 13582 26514
rect 13582 26462 13634 26514
rect 13634 26462 13636 26514
rect 13580 26460 13636 26462
rect 13356 26348 13412 26404
rect 13692 26402 13748 26404
rect 13692 26350 13694 26402
rect 13694 26350 13746 26402
rect 13746 26350 13748 26402
rect 13692 26348 13748 26350
rect 13916 26290 13972 26292
rect 13916 26238 13918 26290
rect 13918 26238 13970 26290
rect 13970 26238 13972 26290
rect 13916 26236 13972 26238
rect 13244 24892 13300 24948
rect 15036 27858 15092 27860
rect 15036 27806 15038 27858
rect 15038 27806 15090 27858
rect 15090 27806 15092 27858
rect 15036 27804 15092 27806
rect 15260 27916 15316 27972
rect 14364 26962 14420 26964
rect 14364 26910 14366 26962
rect 14366 26910 14418 26962
rect 14418 26910 14420 26962
rect 14364 26908 14420 26910
rect 14140 26124 14196 26180
rect 15148 26962 15204 26964
rect 15148 26910 15150 26962
rect 15150 26910 15202 26962
rect 15202 26910 15204 26962
rect 15148 26908 15204 26910
rect 15596 27244 15652 27300
rect 14700 26124 14756 26180
rect 14588 25900 14644 25956
rect 13020 24722 13076 24724
rect 13020 24670 13022 24722
rect 13022 24670 13074 24722
rect 13074 24670 13076 24722
rect 13020 24668 13076 24670
rect 12908 23884 12964 23940
rect 13692 24722 13748 24724
rect 13692 24670 13694 24722
rect 13694 24670 13746 24722
rect 13746 24670 13748 24722
rect 13692 24668 13748 24670
rect 14364 24722 14420 24724
rect 14364 24670 14366 24722
rect 14366 24670 14418 24722
rect 14418 24670 14420 24722
rect 14364 24668 14420 24670
rect 14028 23938 14084 23940
rect 14028 23886 14030 23938
rect 14030 23886 14082 23938
rect 14082 23886 14084 23938
rect 14028 23884 14084 23886
rect 14812 25900 14868 25956
rect 14924 24556 14980 24612
rect 13468 23154 13524 23156
rect 13468 23102 13470 23154
rect 13470 23102 13522 23154
rect 13522 23102 13524 23154
rect 13468 23100 13524 23102
rect 13916 23100 13972 23156
rect 12684 22764 12740 22820
rect 12572 22594 12628 22596
rect 12572 22542 12574 22594
rect 12574 22542 12626 22594
rect 12626 22542 12628 22594
rect 12572 22540 12628 22542
rect 12012 20524 12068 20580
rect 12348 18172 12404 18228
rect 11340 16098 11396 16100
rect 11340 16046 11342 16098
rect 11342 16046 11394 16098
rect 11394 16046 11396 16098
rect 11340 16044 11396 16046
rect 11228 15874 11284 15876
rect 11228 15822 11230 15874
rect 11230 15822 11282 15874
rect 11282 15822 11284 15874
rect 11228 15820 11284 15822
rect 12460 17890 12516 17892
rect 12460 17838 12462 17890
rect 12462 17838 12514 17890
rect 12514 17838 12516 17890
rect 12460 17836 12516 17838
rect 12572 17554 12628 17556
rect 12572 17502 12574 17554
rect 12574 17502 12626 17554
rect 12626 17502 12628 17554
rect 12572 17500 12628 17502
rect 12460 17442 12516 17444
rect 12460 17390 12462 17442
rect 12462 17390 12514 17442
rect 12514 17390 12516 17442
rect 12460 17388 12516 17390
rect 12348 16940 12404 16996
rect 13356 22652 13412 22708
rect 12908 22316 12964 22372
rect 12796 22258 12852 22260
rect 12796 22206 12798 22258
rect 12798 22206 12850 22258
rect 12850 22206 12852 22258
rect 12796 22204 12852 22206
rect 13804 22482 13860 22484
rect 13804 22430 13806 22482
rect 13806 22430 13858 22482
rect 13858 22430 13860 22482
rect 13804 22428 13860 22430
rect 13692 22370 13748 22372
rect 13692 22318 13694 22370
rect 13694 22318 13746 22370
rect 13746 22318 13748 22370
rect 13692 22316 13748 22318
rect 13916 22092 13972 22148
rect 13356 20860 13412 20916
rect 13020 20524 13076 20580
rect 13020 20076 13076 20132
rect 12796 17388 12852 17444
rect 12124 15932 12180 15988
rect 11900 15820 11956 15876
rect 11004 15372 11060 15428
rect 11228 15202 11284 15204
rect 11228 15150 11230 15202
rect 11230 15150 11282 15202
rect 11282 15150 11284 15202
rect 11228 15148 11284 15150
rect 10872 14922 10928 14924
rect 10872 14870 10874 14922
rect 10874 14870 10926 14922
rect 10926 14870 10928 14922
rect 10872 14868 10928 14870
rect 10976 14922 11032 14924
rect 10976 14870 10978 14922
rect 10978 14870 11030 14922
rect 11030 14870 11032 14922
rect 10976 14868 11032 14870
rect 11080 14922 11136 14924
rect 11080 14870 11082 14922
rect 11082 14870 11134 14922
rect 11134 14870 11136 14922
rect 11080 14868 11136 14870
rect 11452 13746 11508 13748
rect 11452 13694 11454 13746
rect 11454 13694 11506 13746
rect 11506 13694 11508 13746
rect 11452 13692 11508 13694
rect 12348 15874 12404 15876
rect 12348 15822 12350 15874
rect 12350 15822 12402 15874
rect 12402 15822 12404 15874
rect 12348 15820 12404 15822
rect 12348 15148 12404 15204
rect 12572 15986 12628 15988
rect 12572 15934 12574 15986
rect 12574 15934 12626 15986
rect 12626 15934 12628 15986
rect 12572 15932 12628 15934
rect 12684 15596 12740 15652
rect 12908 15820 12964 15876
rect 12684 15426 12740 15428
rect 12684 15374 12686 15426
rect 12686 15374 12738 15426
rect 12738 15374 12740 15426
rect 12684 15372 12740 15374
rect 12460 14700 12516 14756
rect 14028 20636 14084 20692
rect 13916 20578 13972 20580
rect 13916 20526 13918 20578
rect 13918 20526 13970 20578
rect 13970 20526 13972 20578
rect 13916 20524 13972 20526
rect 13916 19906 13972 19908
rect 13916 19854 13918 19906
rect 13918 19854 13970 19906
rect 13970 19854 13972 19906
rect 13916 19852 13972 19854
rect 13804 19404 13860 19460
rect 13244 18562 13300 18564
rect 13244 18510 13246 18562
rect 13246 18510 13298 18562
rect 13298 18510 13300 18562
rect 13244 18508 13300 18510
rect 13468 18338 13524 18340
rect 13468 18286 13470 18338
rect 13470 18286 13522 18338
rect 13522 18286 13524 18338
rect 13468 18284 13524 18286
rect 15260 26460 15316 26516
rect 15148 26348 15204 26404
rect 15260 26124 15316 26180
rect 16492 27580 16548 27636
rect 16492 27132 16548 27188
rect 17052 27132 17108 27188
rect 15148 25618 15204 25620
rect 15148 25566 15150 25618
rect 15150 25566 15202 25618
rect 15202 25566 15204 25618
rect 15148 25564 15204 25566
rect 14812 22540 14868 22596
rect 14924 22258 14980 22260
rect 14924 22206 14926 22258
rect 14926 22206 14978 22258
rect 14978 22206 14980 22258
rect 14924 22204 14980 22206
rect 16156 26962 16212 26964
rect 16156 26910 16158 26962
rect 16158 26910 16210 26962
rect 16210 26910 16212 26962
rect 16156 26908 16212 26910
rect 15932 26460 15988 26516
rect 16156 26348 16212 26404
rect 16044 26236 16100 26292
rect 15708 25900 15764 25956
rect 16156 25564 16212 25620
rect 15932 25228 15988 25284
rect 15820 24722 15876 24724
rect 15820 24670 15822 24722
rect 15822 24670 15874 24722
rect 15874 24670 15876 24722
rect 15820 24668 15876 24670
rect 16044 24556 16100 24612
rect 15932 24444 15988 24500
rect 15372 21420 15428 21476
rect 14252 20076 14308 20132
rect 14140 20018 14196 20020
rect 14140 19966 14142 20018
rect 14142 19966 14194 20018
rect 14194 19966 14196 20018
rect 14140 19964 14196 19966
rect 15036 19964 15092 20020
rect 14252 19516 14308 19572
rect 14700 19404 14756 19460
rect 15036 19292 15092 19348
rect 15148 19852 15204 19908
rect 15148 18732 15204 18788
rect 14252 18620 14308 18676
rect 14364 17612 14420 17668
rect 13804 17442 13860 17444
rect 13804 17390 13806 17442
rect 13806 17390 13858 17442
rect 13858 17390 13860 17442
rect 13804 17388 13860 17390
rect 13468 17106 13524 17108
rect 13468 17054 13470 17106
rect 13470 17054 13522 17106
rect 13522 17054 13524 17106
rect 13468 17052 13524 17054
rect 13580 16994 13636 16996
rect 13580 16942 13582 16994
rect 13582 16942 13634 16994
rect 13634 16942 13636 16994
rect 13580 16940 13636 16942
rect 12236 14418 12292 14420
rect 12236 14366 12238 14418
rect 12238 14366 12290 14418
rect 12290 14366 12292 14418
rect 12236 14364 12292 14366
rect 12348 14306 12404 14308
rect 12348 14254 12350 14306
rect 12350 14254 12402 14306
rect 12402 14254 12404 14306
rect 12348 14252 12404 14254
rect 11900 13692 11956 13748
rect 12124 13804 12180 13860
rect 11676 13522 11732 13524
rect 11676 13470 11678 13522
rect 11678 13470 11730 13522
rect 11730 13470 11732 13522
rect 11676 13468 11732 13470
rect 10872 13354 10928 13356
rect 10872 13302 10874 13354
rect 10874 13302 10926 13354
rect 10926 13302 10928 13354
rect 10872 13300 10928 13302
rect 10976 13354 11032 13356
rect 10976 13302 10978 13354
rect 10978 13302 11030 13354
rect 11030 13302 11032 13354
rect 10976 13300 11032 13302
rect 11080 13354 11136 13356
rect 11080 13302 11082 13354
rect 11082 13302 11134 13354
rect 11134 13302 11136 13354
rect 11080 13300 11136 13302
rect 11788 12290 11844 12292
rect 11788 12238 11790 12290
rect 11790 12238 11842 12290
rect 11842 12238 11844 12290
rect 11788 12236 11844 12238
rect 10780 11954 10836 11956
rect 10780 11902 10782 11954
rect 10782 11902 10834 11954
rect 10834 11902 10836 11954
rect 10780 11900 10836 11902
rect 10872 11786 10928 11788
rect 10872 11734 10874 11786
rect 10874 11734 10926 11786
rect 10926 11734 10928 11786
rect 10872 11732 10928 11734
rect 10976 11786 11032 11788
rect 10976 11734 10978 11786
rect 10978 11734 11030 11786
rect 11030 11734 11032 11786
rect 10976 11732 11032 11734
rect 11080 11786 11136 11788
rect 11080 11734 11082 11786
rect 11082 11734 11134 11786
rect 11134 11734 11136 11786
rect 11080 11732 11136 11734
rect 12908 13692 12964 13748
rect 12348 13074 12404 13076
rect 12348 13022 12350 13074
rect 12350 13022 12402 13074
rect 12402 13022 12404 13074
rect 12348 13020 12404 13022
rect 12348 12796 12404 12852
rect 13020 12796 13076 12852
rect 12460 12290 12516 12292
rect 12460 12238 12462 12290
rect 12462 12238 12514 12290
rect 12514 12238 12516 12290
rect 12460 12236 12516 12238
rect 12796 12236 12852 12292
rect 12684 12178 12740 12180
rect 12684 12126 12686 12178
rect 12686 12126 12738 12178
rect 12738 12126 12740 12178
rect 12684 12124 12740 12126
rect 12908 11900 12964 11956
rect 10220 10108 10276 10164
rect 11228 10610 11284 10612
rect 11228 10558 11230 10610
rect 11230 10558 11282 10610
rect 11282 10558 11284 10610
rect 11228 10556 11284 10558
rect 10872 10218 10928 10220
rect 10872 10166 10874 10218
rect 10874 10166 10926 10218
rect 10926 10166 10928 10218
rect 10872 10164 10928 10166
rect 10976 10218 11032 10220
rect 10976 10166 10978 10218
rect 10978 10166 11030 10218
rect 11030 10166 11032 10218
rect 10976 10164 11032 10166
rect 11080 10218 11136 10220
rect 11080 10166 11082 10218
rect 11082 10166 11134 10218
rect 11134 10166 11136 10218
rect 11080 10164 11136 10166
rect 10444 9884 10500 9940
rect 11004 9884 11060 9940
rect 10556 9436 10612 9492
rect 9884 8652 9940 8708
rect 10444 8988 10500 9044
rect 10444 8540 10500 8596
rect 9660 8316 9716 8372
rect 8652 6636 8708 6692
rect 8540 6076 8596 6132
rect 8652 6412 8708 6468
rect 8428 5964 8484 6020
rect 8652 5906 8708 5908
rect 8652 5854 8654 5906
rect 8654 5854 8706 5906
rect 8706 5854 8708 5906
rect 8652 5852 8708 5854
rect 8652 5346 8708 5348
rect 8652 5294 8654 5346
rect 8654 5294 8706 5346
rect 8706 5294 8708 5346
rect 8652 5292 8708 5294
rect 9772 8258 9828 8260
rect 9772 8206 9774 8258
rect 9774 8206 9826 8258
rect 9826 8206 9828 8258
rect 9772 8204 9828 8206
rect 9324 8092 9380 8148
rect 9996 8034 10052 8036
rect 9996 7982 9998 8034
rect 9998 7982 10050 8034
rect 10050 7982 10052 8034
rect 9996 7980 10052 7982
rect 10108 7868 10164 7924
rect 10892 9100 10948 9156
rect 10872 8650 10928 8652
rect 10872 8598 10874 8650
rect 10874 8598 10926 8650
rect 10926 8598 10928 8650
rect 10872 8596 10928 8598
rect 10976 8650 11032 8652
rect 10976 8598 10978 8650
rect 10978 8598 11030 8650
rect 11030 8598 11032 8650
rect 10976 8596 11032 8598
rect 11080 8650 11136 8652
rect 11080 8598 11082 8650
rect 11082 8598 11134 8650
rect 11134 8598 11136 8650
rect 11080 8596 11136 8598
rect 10668 8034 10724 8036
rect 10668 7982 10670 8034
rect 10670 7982 10722 8034
rect 10722 7982 10724 8034
rect 10668 7980 10724 7982
rect 10668 7756 10724 7812
rect 10892 7868 10948 7924
rect 9324 6860 9380 6916
rect 9772 7586 9828 7588
rect 9772 7534 9774 7586
rect 9774 7534 9826 7586
rect 9826 7534 9828 7586
rect 9772 7532 9828 7534
rect 9660 6748 9716 6804
rect 9324 6690 9380 6692
rect 9324 6638 9326 6690
rect 9326 6638 9378 6690
rect 9378 6638 9380 6690
rect 9324 6636 9380 6638
rect 9436 6524 9492 6580
rect 8876 6076 8932 6132
rect 9436 5964 9492 6020
rect 8988 5794 9044 5796
rect 8988 5742 8990 5794
rect 8990 5742 9042 5794
rect 9042 5742 9044 5794
rect 8988 5740 9044 5742
rect 8764 5180 8820 5236
rect 9548 6076 9604 6132
rect 8652 4338 8708 4340
rect 8652 4286 8654 4338
rect 8654 4286 8706 4338
rect 8706 4286 8708 4338
rect 8652 4284 8708 4286
rect 9100 4226 9156 4228
rect 9100 4174 9102 4226
rect 9102 4174 9154 4226
rect 9154 4174 9156 4226
rect 9100 4172 9156 4174
rect 8204 3442 8260 3444
rect 8204 3390 8206 3442
rect 8206 3390 8258 3442
rect 8258 3390 8260 3442
rect 8204 3388 8260 3390
rect 9100 3388 9156 3444
rect 7532 3276 7588 3332
rect 9884 6524 9940 6580
rect 10872 7082 10928 7084
rect 10872 7030 10874 7082
rect 10874 7030 10926 7082
rect 10926 7030 10928 7082
rect 10872 7028 10928 7030
rect 10976 7082 11032 7084
rect 10976 7030 10978 7082
rect 10978 7030 11030 7082
rect 11030 7030 11032 7082
rect 10976 7028 11032 7030
rect 11080 7082 11136 7084
rect 11080 7030 11082 7082
rect 11082 7030 11134 7082
rect 11134 7030 11136 7082
rect 11080 7028 11136 7030
rect 9996 6748 10052 6804
rect 10220 6636 10276 6692
rect 10108 6466 10164 6468
rect 10108 6414 10110 6466
rect 10110 6414 10162 6466
rect 10162 6414 10164 6466
rect 10108 6412 10164 6414
rect 9996 6188 10052 6244
rect 9884 6076 9940 6132
rect 9772 5292 9828 5348
rect 10444 6690 10500 6692
rect 10444 6638 10446 6690
rect 10446 6638 10498 6690
rect 10498 6638 10500 6690
rect 10444 6636 10500 6638
rect 10892 6690 10948 6692
rect 10892 6638 10894 6690
rect 10894 6638 10946 6690
rect 10946 6638 10948 6690
rect 10892 6636 10948 6638
rect 10332 6466 10388 6468
rect 10332 6414 10334 6466
rect 10334 6414 10386 6466
rect 10386 6414 10388 6466
rect 10332 6412 10388 6414
rect 11340 6466 11396 6468
rect 11340 6414 11342 6466
rect 11342 6414 11394 6466
rect 11394 6414 11396 6466
rect 11340 6412 11396 6414
rect 11116 6188 11172 6244
rect 10444 6130 10500 6132
rect 10444 6078 10446 6130
rect 10446 6078 10498 6130
rect 10498 6078 10500 6130
rect 10444 6076 10500 6078
rect 10332 5964 10388 6020
rect 9996 5794 10052 5796
rect 9996 5742 9998 5794
rect 9998 5742 10050 5794
rect 10050 5742 10052 5794
rect 9996 5740 10052 5742
rect 9660 3612 9716 3668
rect 9996 5068 10052 5124
rect 10872 5514 10928 5516
rect 10872 5462 10874 5514
rect 10874 5462 10926 5514
rect 10926 5462 10928 5514
rect 10872 5460 10928 5462
rect 10976 5514 11032 5516
rect 10976 5462 10978 5514
rect 10978 5462 11030 5514
rect 11030 5462 11032 5514
rect 10976 5460 11032 5462
rect 11080 5514 11136 5516
rect 11080 5462 11082 5514
rect 11082 5462 11134 5514
rect 11134 5462 11136 5514
rect 11080 5460 11136 5462
rect 10332 5068 10388 5124
rect 10668 5122 10724 5124
rect 10668 5070 10670 5122
rect 10670 5070 10722 5122
rect 10722 5070 10724 5122
rect 10668 5068 10724 5070
rect 9996 3500 10052 3556
rect 13916 16156 13972 16212
rect 13580 15874 13636 15876
rect 13580 15822 13582 15874
rect 13582 15822 13634 15874
rect 13634 15822 13636 15874
rect 13580 15820 13636 15822
rect 13580 15596 13636 15652
rect 13804 15148 13860 15204
rect 14476 17388 14532 17444
rect 14588 18060 14644 18116
rect 15820 18562 15876 18564
rect 15820 18510 15822 18562
rect 15822 18510 15874 18562
rect 15874 18510 15876 18562
rect 15820 18508 15876 18510
rect 15372 18172 15428 18228
rect 15260 18060 15316 18116
rect 14812 17442 14868 17444
rect 14812 17390 14814 17442
rect 14814 17390 14866 17442
rect 14866 17390 14868 17442
rect 14812 17388 14868 17390
rect 14588 17106 14644 17108
rect 14588 17054 14590 17106
rect 14590 17054 14642 17106
rect 14642 17054 14644 17106
rect 14588 17052 14644 17054
rect 14812 16940 14868 16996
rect 14364 16210 14420 16212
rect 14364 16158 14366 16210
rect 14366 16158 14418 16210
rect 14418 16158 14420 16210
rect 14364 16156 14420 16158
rect 17052 26684 17108 26740
rect 16828 26402 16884 26404
rect 16828 26350 16830 26402
rect 16830 26350 16882 26402
rect 16882 26350 16884 26402
rect 16828 26348 16884 26350
rect 17052 26290 17108 26292
rect 17052 26238 17054 26290
rect 17054 26238 17106 26290
rect 17106 26238 17108 26290
rect 17052 26236 17108 26238
rect 18284 29538 18340 29540
rect 18284 29486 18286 29538
rect 18286 29486 18338 29538
rect 18338 29486 18340 29538
rect 18284 29484 18340 29486
rect 17836 28754 17892 28756
rect 17836 28702 17838 28754
rect 17838 28702 17890 28754
rect 17890 28702 17892 28754
rect 17836 28700 17892 28702
rect 18620 28588 18676 28644
rect 17388 28530 17444 28532
rect 17388 28478 17390 28530
rect 17390 28478 17442 28530
rect 17442 28478 17444 28530
rect 17388 28476 17444 28478
rect 17612 28364 17668 28420
rect 17164 26124 17220 26180
rect 17500 27074 17556 27076
rect 17500 27022 17502 27074
rect 17502 27022 17554 27074
rect 17554 27022 17556 27074
rect 17500 27020 17556 27022
rect 17500 26348 17556 26404
rect 16268 24780 16324 24836
rect 15932 17724 15988 17780
rect 17948 28364 18004 28420
rect 18284 28364 18340 28420
rect 17948 27634 18004 27636
rect 17948 27582 17950 27634
rect 17950 27582 18002 27634
rect 18002 27582 18004 27634
rect 17948 27580 18004 27582
rect 18060 26684 18116 26740
rect 18172 26850 18228 26852
rect 18172 26798 18174 26850
rect 18174 26798 18226 26850
rect 18226 26798 18228 26850
rect 18172 26796 18228 26798
rect 18172 26348 18228 26404
rect 18844 29484 18900 29540
rect 19964 30994 20020 30996
rect 19964 30942 19966 30994
rect 19966 30942 20018 30994
rect 20018 30942 20020 30994
rect 19964 30940 20020 30942
rect 19740 30604 19796 30660
rect 20532 29818 20588 29820
rect 20532 29766 20534 29818
rect 20534 29766 20586 29818
rect 20586 29766 20588 29818
rect 20532 29764 20588 29766
rect 20636 29818 20692 29820
rect 20636 29766 20638 29818
rect 20638 29766 20690 29818
rect 20690 29766 20692 29818
rect 20636 29764 20692 29766
rect 20740 29818 20796 29820
rect 20740 29766 20742 29818
rect 20742 29766 20794 29818
rect 20794 29766 20796 29818
rect 20740 29764 20796 29766
rect 21980 31612 22036 31668
rect 22988 29986 23044 29988
rect 22988 29934 22990 29986
rect 22990 29934 23042 29986
rect 23042 29934 23044 29986
rect 22988 29932 23044 29934
rect 21308 29372 21364 29428
rect 18956 28700 19012 28756
rect 19180 28588 19236 28644
rect 19068 28476 19124 28532
rect 19068 27074 19124 27076
rect 19068 27022 19070 27074
rect 19070 27022 19122 27074
rect 19122 27022 19124 27074
rect 19068 27020 19124 27022
rect 22428 29426 22484 29428
rect 22428 29374 22430 29426
rect 22430 29374 22482 29426
rect 22482 29374 22484 29426
rect 22428 29372 22484 29374
rect 23100 29426 23156 29428
rect 23100 29374 23102 29426
rect 23102 29374 23154 29426
rect 23154 29374 23156 29426
rect 23100 29372 23156 29374
rect 21532 29314 21588 29316
rect 21532 29262 21534 29314
rect 21534 29262 21586 29314
rect 21586 29262 21588 29314
rect 21532 29260 21588 29262
rect 22204 29314 22260 29316
rect 22204 29262 22206 29314
rect 22206 29262 22258 29314
rect 22258 29262 22260 29314
rect 22204 29260 22260 29262
rect 22876 29260 22932 29316
rect 21756 29148 21812 29204
rect 20188 28364 20244 28420
rect 20532 28250 20588 28252
rect 20532 28198 20534 28250
rect 20534 28198 20586 28250
rect 20586 28198 20588 28250
rect 20532 28196 20588 28198
rect 20636 28250 20692 28252
rect 20636 28198 20638 28250
rect 20638 28198 20690 28250
rect 20690 28198 20692 28250
rect 20636 28196 20692 28198
rect 20740 28250 20796 28252
rect 20740 28198 20742 28250
rect 20742 28198 20794 28250
rect 20794 28198 20796 28250
rect 20740 28196 20796 28198
rect 21196 28252 21252 28308
rect 20076 26908 20132 26964
rect 18508 26348 18564 26404
rect 17948 26236 18004 26292
rect 18284 26124 18340 26180
rect 18396 25506 18452 25508
rect 18396 25454 18398 25506
rect 18398 25454 18450 25506
rect 18450 25454 18452 25506
rect 18396 25452 18452 25454
rect 17612 24220 17668 24276
rect 18844 26796 18900 26852
rect 18956 26684 19012 26740
rect 20412 26908 20468 26964
rect 19628 26850 19684 26852
rect 19628 26798 19630 26850
rect 19630 26798 19682 26850
rect 19682 26798 19684 26850
rect 19628 26796 19684 26798
rect 19516 26290 19572 26292
rect 19516 26238 19518 26290
rect 19518 26238 19570 26290
rect 19570 26238 19572 26290
rect 19516 26236 19572 26238
rect 19292 25618 19348 25620
rect 19292 25566 19294 25618
rect 19294 25566 19346 25618
rect 19346 25566 19348 25618
rect 19292 25564 19348 25566
rect 19852 26348 19908 26404
rect 20188 26236 20244 26292
rect 17276 23436 17332 23492
rect 15260 16716 15316 16772
rect 15372 17276 15428 17332
rect 15148 16268 15204 16324
rect 14588 15932 14644 15988
rect 14476 15538 14532 15540
rect 14476 15486 14478 15538
rect 14478 15486 14530 15538
rect 14530 15486 14532 15538
rect 14476 15484 14532 15486
rect 14252 15260 14308 15316
rect 13356 13020 13412 13076
rect 13468 14364 13524 14420
rect 14364 14418 14420 14420
rect 14364 14366 14366 14418
rect 14366 14366 14418 14418
rect 14418 14366 14420 14418
rect 14364 14364 14420 14366
rect 13804 13468 13860 13524
rect 13692 13020 13748 13076
rect 15148 15708 15204 15764
rect 15708 16716 15764 16772
rect 15708 16044 15764 16100
rect 15372 15484 15428 15540
rect 15932 15874 15988 15876
rect 15932 15822 15934 15874
rect 15934 15822 15986 15874
rect 15986 15822 15988 15874
rect 15932 15820 15988 15822
rect 14812 14812 14868 14868
rect 14588 14418 14644 14420
rect 14588 14366 14590 14418
rect 14590 14366 14642 14418
rect 14642 14366 14644 14418
rect 14588 14364 14644 14366
rect 14700 14252 14756 14308
rect 15596 14418 15652 14420
rect 15596 14366 15598 14418
rect 15598 14366 15650 14418
rect 15650 14366 15652 14418
rect 15596 14364 15652 14366
rect 15148 14306 15204 14308
rect 15148 14254 15150 14306
rect 15150 14254 15202 14306
rect 15202 14254 15204 14306
rect 15148 14252 15204 14254
rect 16156 21532 16212 21588
rect 16492 22258 16548 22260
rect 16492 22206 16494 22258
rect 16494 22206 16546 22258
rect 16546 22206 16548 22258
rect 16492 22204 16548 22206
rect 18060 23548 18116 23604
rect 18620 23938 18676 23940
rect 18620 23886 18622 23938
rect 18622 23886 18674 23938
rect 18674 23886 18676 23938
rect 18620 23884 18676 23886
rect 20300 25564 20356 25620
rect 20076 25228 20132 25284
rect 19516 24050 19572 24052
rect 19516 23998 19518 24050
rect 19518 23998 19570 24050
rect 19570 23998 19572 24050
rect 19516 23996 19572 23998
rect 19292 23884 19348 23940
rect 19852 24220 19908 24276
rect 18284 23436 18340 23492
rect 18060 23212 18116 23268
rect 19180 23436 19236 23492
rect 18284 22988 18340 23044
rect 17836 22876 17892 22932
rect 16716 21586 16772 21588
rect 16716 21534 16718 21586
rect 16718 21534 16770 21586
rect 16770 21534 16772 21586
rect 16716 21532 16772 21534
rect 16156 19516 16212 19572
rect 17724 20524 17780 20580
rect 17500 19964 17556 20020
rect 16940 19346 16996 19348
rect 16940 19294 16942 19346
rect 16942 19294 16994 19346
rect 16994 19294 16996 19346
rect 16940 19292 16996 19294
rect 16604 19180 16660 19236
rect 16268 18732 16324 18788
rect 16380 18620 16436 18676
rect 16492 18956 16548 19012
rect 16380 18396 16436 18452
rect 16156 16882 16212 16884
rect 16156 16830 16158 16882
rect 16158 16830 16210 16882
rect 16210 16830 16212 16882
rect 16156 16828 16212 16830
rect 16380 16828 16436 16884
rect 16268 16268 16324 16324
rect 17052 19234 17108 19236
rect 17052 19182 17054 19234
rect 17054 19182 17106 19234
rect 17106 19182 17108 19234
rect 17052 19180 17108 19182
rect 16940 18732 16996 18788
rect 16716 18396 16772 18452
rect 16828 18674 16884 18676
rect 16828 18622 16830 18674
rect 16830 18622 16882 18674
rect 16882 18622 16884 18674
rect 16828 18620 16884 18622
rect 17276 19346 17332 19348
rect 17276 19294 17278 19346
rect 17278 19294 17330 19346
rect 17330 19294 17332 19346
rect 17276 19292 17332 19294
rect 17164 18732 17220 18788
rect 17052 18396 17108 18452
rect 16940 18060 16996 18116
rect 16492 16156 16548 16212
rect 16716 16716 16772 16772
rect 17052 17106 17108 17108
rect 17052 17054 17054 17106
rect 17054 17054 17106 17106
rect 17106 17054 17108 17106
rect 17052 17052 17108 17054
rect 16940 16940 16996 16996
rect 19068 23266 19124 23268
rect 19068 23214 19070 23266
rect 19070 23214 19122 23266
rect 19122 23214 19124 23266
rect 19068 23212 19124 23214
rect 18508 22876 18564 22932
rect 19964 23212 20020 23268
rect 20748 26962 20804 26964
rect 20748 26910 20750 26962
rect 20750 26910 20802 26962
rect 20802 26910 20804 26962
rect 20748 26908 20804 26910
rect 20524 26796 20580 26852
rect 20532 26682 20588 26684
rect 20532 26630 20534 26682
rect 20534 26630 20586 26682
rect 20586 26630 20588 26682
rect 20532 26628 20588 26630
rect 20636 26682 20692 26684
rect 20636 26630 20638 26682
rect 20638 26630 20690 26682
rect 20690 26630 20692 26682
rect 20636 26628 20692 26630
rect 20740 26682 20796 26684
rect 20740 26630 20742 26682
rect 20742 26630 20794 26682
rect 20794 26630 20796 26682
rect 20740 26628 20796 26630
rect 20636 26402 20692 26404
rect 20636 26350 20638 26402
rect 20638 26350 20690 26402
rect 20690 26350 20692 26402
rect 20636 26348 20692 26350
rect 20524 25788 20580 25844
rect 20636 25564 20692 25620
rect 20524 25228 20580 25284
rect 20860 25228 20916 25284
rect 20532 25114 20588 25116
rect 20532 25062 20534 25114
rect 20534 25062 20586 25114
rect 20586 25062 20588 25114
rect 20532 25060 20588 25062
rect 20636 25114 20692 25116
rect 20636 25062 20638 25114
rect 20638 25062 20690 25114
rect 20690 25062 20692 25114
rect 20636 25060 20692 25062
rect 20740 25114 20796 25116
rect 20740 25062 20742 25114
rect 20742 25062 20794 25114
rect 20794 25062 20796 25114
rect 20740 25060 20796 25062
rect 20532 23546 20588 23548
rect 20188 23436 20244 23492
rect 20532 23494 20534 23546
rect 20534 23494 20586 23546
rect 20586 23494 20588 23546
rect 20532 23492 20588 23494
rect 20636 23546 20692 23548
rect 20636 23494 20638 23546
rect 20638 23494 20690 23546
rect 20690 23494 20692 23546
rect 20636 23492 20692 23494
rect 20740 23546 20796 23548
rect 20740 23494 20742 23546
rect 20742 23494 20794 23546
rect 20794 23494 20796 23546
rect 20740 23492 20796 23494
rect 21868 27858 21924 27860
rect 21868 27806 21870 27858
rect 21870 27806 21922 27858
rect 21922 27806 21924 27858
rect 21868 27804 21924 27806
rect 21420 26908 21476 26964
rect 23324 35698 23380 35700
rect 23324 35646 23326 35698
rect 23326 35646 23378 35698
rect 23378 35646 23380 35698
rect 23324 35644 23380 35646
rect 23660 35644 23716 35700
rect 23548 35084 23604 35140
rect 27804 36540 27860 36596
rect 25228 36428 25284 36484
rect 30192 36874 30248 36876
rect 30192 36822 30194 36874
rect 30194 36822 30246 36874
rect 30246 36822 30248 36874
rect 30192 36820 30248 36822
rect 30296 36874 30352 36876
rect 30296 36822 30298 36874
rect 30298 36822 30350 36874
rect 30350 36822 30352 36874
rect 30296 36820 30352 36822
rect 30400 36874 30456 36876
rect 30400 36822 30402 36874
rect 30402 36822 30454 36874
rect 30454 36822 30456 36874
rect 30400 36820 30456 36822
rect 33964 37884 34020 37940
rect 33964 36652 34020 36708
rect 33516 36594 33572 36596
rect 33516 36542 33518 36594
rect 33518 36542 33570 36594
rect 33570 36542 33572 36594
rect 33516 36540 33572 36542
rect 25788 36370 25844 36372
rect 25788 36318 25790 36370
rect 25790 36318 25842 36370
rect 25842 36318 25844 36370
rect 25788 36316 25844 36318
rect 27356 36316 27412 36372
rect 25340 34914 25396 34916
rect 25340 34862 25342 34914
rect 25342 34862 25394 34914
rect 25394 34862 25396 34914
rect 25340 34860 25396 34862
rect 25004 34690 25060 34692
rect 25004 34638 25006 34690
rect 25006 34638 25058 34690
rect 25058 34638 25060 34690
rect 25004 34636 25060 34638
rect 24780 34412 24836 34468
rect 23884 34130 23940 34132
rect 23884 34078 23886 34130
rect 23886 34078 23938 34130
rect 23938 34078 23940 34130
rect 23884 34076 23940 34078
rect 23324 33628 23380 33684
rect 23436 33852 23492 33908
rect 23884 33852 23940 33908
rect 24332 33628 24388 33684
rect 24108 32508 24164 32564
rect 23436 32450 23492 32452
rect 23436 32398 23438 32450
rect 23438 32398 23490 32450
rect 23490 32398 23492 32450
rect 23436 32396 23492 32398
rect 23996 32450 24052 32452
rect 23996 32398 23998 32450
rect 23998 32398 24050 32450
rect 24050 32398 24052 32450
rect 23996 32396 24052 32398
rect 23548 31500 23604 31556
rect 24556 31500 24612 31556
rect 24892 34242 24948 34244
rect 24892 34190 24894 34242
rect 24894 34190 24946 34242
rect 24946 34190 24948 34242
rect 24892 34188 24948 34190
rect 26124 36258 26180 36260
rect 26124 36206 26126 36258
rect 26126 36206 26178 36258
rect 26178 36206 26180 36258
rect 26124 36204 26180 36206
rect 26796 35922 26852 35924
rect 26796 35870 26798 35922
rect 26798 35870 26850 35922
rect 26850 35870 26852 35922
rect 26796 35868 26852 35870
rect 25900 35532 25956 35588
rect 26012 35756 26068 35812
rect 26460 35756 26516 35812
rect 27468 35922 27524 35924
rect 27468 35870 27470 35922
rect 27470 35870 27522 35922
rect 27522 35870 27524 35922
rect 27468 35868 27524 35870
rect 27468 35644 27524 35700
rect 26236 35586 26292 35588
rect 26236 35534 26238 35586
rect 26238 35534 26290 35586
rect 26290 35534 26292 35586
rect 26236 35532 26292 35534
rect 28588 36370 28644 36372
rect 28588 36318 28590 36370
rect 28590 36318 28642 36370
rect 28642 36318 28644 36370
rect 28588 36316 28644 36318
rect 30492 36316 30548 36372
rect 29596 36204 29652 36260
rect 28476 35922 28532 35924
rect 28476 35870 28478 35922
rect 28478 35870 28530 35922
rect 28530 35870 28532 35922
rect 28476 35868 28532 35870
rect 28588 35810 28644 35812
rect 28588 35758 28590 35810
rect 28590 35758 28642 35810
rect 28642 35758 28644 35810
rect 28588 35756 28644 35758
rect 28476 35698 28532 35700
rect 28476 35646 28478 35698
rect 28478 35646 28530 35698
rect 28530 35646 28532 35698
rect 28476 35644 28532 35646
rect 25452 34748 25508 34804
rect 25676 34690 25732 34692
rect 25676 34638 25678 34690
rect 25678 34638 25730 34690
rect 25730 34638 25732 34690
rect 25676 34636 25732 34638
rect 26012 34636 26068 34692
rect 26796 34914 26852 34916
rect 26796 34862 26798 34914
rect 26798 34862 26850 34914
rect 26850 34862 26852 34914
rect 26796 34860 26852 34862
rect 27132 34860 27188 34916
rect 26460 34188 26516 34244
rect 25900 34076 25956 34132
rect 26236 34130 26292 34132
rect 26236 34078 26238 34130
rect 26238 34078 26290 34130
rect 26290 34078 26292 34130
rect 26236 34076 26292 34078
rect 28364 34860 28420 34916
rect 27468 34354 27524 34356
rect 27468 34302 27470 34354
rect 27470 34302 27522 34354
rect 27522 34302 27524 34354
rect 27468 34300 27524 34302
rect 27244 34242 27300 34244
rect 27244 34190 27246 34242
rect 27246 34190 27298 34242
rect 27298 34190 27300 34242
rect 27244 34188 27300 34190
rect 26460 33852 26516 33908
rect 29820 35698 29876 35700
rect 29820 35646 29822 35698
rect 29822 35646 29874 35698
rect 29874 35646 29876 35698
rect 29820 35644 29876 35646
rect 30192 35306 30248 35308
rect 30192 35254 30194 35306
rect 30194 35254 30246 35306
rect 30246 35254 30248 35306
rect 30192 35252 30248 35254
rect 30296 35306 30352 35308
rect 30296 35254 30298 35306
rect 30298 35254 30350 35306
rect 30350 35254 30352 35306
rect 30296 35252 30352 35254
rect 30400 35306 30456 35308
rect 30400 35254 30402 35306
rect 30402 35254 30454 35306
rect 30454 35254 30456 35306
rect 30400 35252 30456 35254
rect 30268 35084 30324 35140
rect 28476 34802 28532 34804
rect 28476 34750 28478 34802
rect 28478 34750 28530 34802
rect 28530 34750 28532 34802
rect 28476 34748 28532 34750
rect 29596 34412 29652 34468
rect 31052 35084 31108 35140
rect 30380 34690 30436 34692
rect 30380 34638 30382 34690
rect 30382 34638 30434 34690
rect 30434 34638 30436 34690
rect 30380 34636 30436 34638
rect 30268 34300 30324 34356
rect 28700 33964 28756 34020
rect 28252 33346 28308 33348
rect 28252 33294 28254 33346
rect 28254 33294 28306 33346
rect 28306 33294 28308 33346
rect 28252 33292 28308 33294
rect 27020 33068 27076 33124
rect 24220 31164 24276 31220
rect 23436 29932 23492 29988
rect 23660 29426 23716 29428
rect 23660 29374 23662 29426
rect 23662 29374 23714 29426
rect 23714 29374 23716 29426
rect 23660 29372 23716 29374
rect 23548 29036 23604 29092
rect 24108 29932 24164 29988
rect 23996 29372 24052 29428
rect 25004 30268 25060 30324
rect 24220 29372 24276 29428
rect 24556 29314 24612 29316
rect 24556 29262 24558 29314
rect 24558 29262 24610 29314
rect 24610 29262 24612 29314
rect 24556 29260 24612 29262
rect 24780 28754 24836 28756
rect 24780 28702 24782 28754
rect 24782 28702 24834 28754
rect 24834 28702 24836 28754
rect 24780 28700 24836 28702
rect 23212 28476 23268 28532
rect 23772 28476 23828 28532
rect 22988 28028 23044 28084
rect 23660 28082 23716 28084
rect 23660 28030 23662 28082
rect 23662 28030 23714 28082
rect 23714 28030 23716 28082
rect 23660 28028 23716 28030
rect 22876 27858 22932 27860
rect 22876 27806 22878 27858
rect 22878 27806 22930 27858
rect 22930 27806 22932 27858
rect 22876 27804 22932 27806
rect 22652 27020 22708 27076
rect 22764 27468 22820 27524
rect 21532 26850 21588 26852
rect 21532 26798 21534 26850
rect 21534 26798 21586 26850
rect 21586 26798 21588 26850
rect 21532 26796 21588 26798
rect 21532 26348 21588 26404
rect 22764 26962 22820 26964
rect 22764 26910 22766 26962
rect 22766 26910 22818 26962
rect 22818 26910 22820 26962
rect 22764 26908 22820 26910
rect 22540 26796 22596 26852
rect 24444 28140 24500 28196
rect 24892 28364 24948 28420
rect 23772 27356 23828 27412
rect 23884 27132 23940 27188
rect 23212 27074 23268 27076
rect 23212 27022 23214 27074
rect 23214 27022 23266 27074
rect 23266 27022 23268 27074
rect 23212 27020 23268 27022
rect 23548 26908 23604 26964
rect 22988 26514 23044 26516
rect 22988 26462 22990 26514
rect 22990 26462 23042 26514
rect 23042 26462 23044 26514
rect 22988 26460 23044 26462
rect 21868 26348 21924 26404
rect 21756 25788 21812 25844
rect 22428 26178 22484 26180
rect 22428 26126 22430 26178
rect 22430 26126 22482 26178
rect 22482 26126 22484 26178
rect 22428 26124 22484 26126
rect 21980 25506 22036 25508
rect 21980 25454 21982 25506
rect 21982 25454 22034 25506
rect 22034 25454 22036 25506
rect 21980 25452 22036 25454
rect 21868 25394 21924 25396
rect 21868 25342 21870 25394
rect 21870 25342 21922 25394
rect 21922 25342 21924 25394
rect 21868 25340 21924 25342
rect 22092 25282 22148 25284
rect 22092 25230 22094 25282
rect 22094 25230 22146 25282
rect 22146 25230 22148 25282
rect 22092 25228 22148 25230
rect 22428 25228 22484 25284
rect 22652 25228 22708 25284
rect 22316 25004 22372 25060
rect 21868 24892 21924 24948
rect 21868 23884 21924 23940
rect 21868 23660 21924 23716
rect 19404 23154 19460 23156
rect 19404 23102 19406 23154
rect 19406 23102 19458 23154
rect 19458 23102 19460 23154
rect 19404 23100 19460 23102
rect 19180 22876 19236 22932
rect 20076 22258 20132 22260
rect 20076 22206 20078 22258
rect 20078 22206 20130 22258
rect 20130 22206 20132 22258
rect 20076 22204 20132 22206
rect 18172 21698 18228 21700
rect 18172 21646 18174 21698
rect 18174 21646 18226 21698
rect 18226 21646 18228 21698
rect 18172 21644 18228 21646
rect 17948 20802 18004 20804
rect 17948 20750 17950 20802
rect 17950 20750 18002 20802
rect 18002 20750 18004 20802
rect 17948 20748 18004 20750
rect 18284 20300 18340 20356
rect 19516 21586 19572 21588
rect 19516 21534 19518 21586
rect 19518 21534 19570 21586
rect 19570 21534 19572 21586
rect 19516 21532 19572 21534
rect 19964 21474 20020 21476
rect 19964 21422 19966 21474
rect 19966 21422 20018 21474
rect 20018 21422 20020 21474
rect 19964 21420 20020 21422
rect 20188 21308 20244 21364
rect 20636 23100 20692 23156
rect 20300 21644 20356 21700
rect 19964 20860 20020 20916
rect 19852 20748 19908 20804
rect 18396 20188 18452 20244
rect 18620 20636 18676 20692
rect 18172 19122 18228 19124
rect 18172 19070 18174 19122
rect 18174 19070 18226 19122
rect 18226 19070 18228 19122
rect 18172 19068 18228 19070
rect 18060 18674 18116 18676
rect 18060 18622 18062 18674
rect 18062 18622 18114 18674
rect 18114 18622 18116 18674
rect 18060 18620 18116 18622
rect 19628 20690 19684 20692
rect 19628 20638 19630 20690
rect 19630 20638 19682 20690
rect 19682 20638 19684 20690
rect 19628 20636 19684 20638
rect 18732 20578 18788 20580
rect 18732 20526 18734 20578
rect 18734 20526 18786 20578
rect 18786 20526 18788 20578
rect 18732 20524 18788 20526
rect 18844 19404 18900 19460
rect 18620 19068 18676 19124
rect 18508 18844 18564 18900
rect 19404 20188 19460 20244
rect 19180 20018 19236 20020
rect 19180 19966 19182 20018
rect 19182 19966 19234 20018
rect 19234 19966 19236 20018
rect 19180 19964 19236 19966
rect 19068 19404 19124 19460
rect 18732 18732 18788 18788
rect 16828 16828 16884 16884
rect 17836 18562 17892 18564
rect 17836 18510 17838 18562
rect 17838 18510 17890 18562
rect 17890 18510 17892 18562
rect 17836 18508 17892 18510
rect 18396 18450 18452 18452
rect 18396 18398 18398 18450
rect 18398 18398 18450 18450
rect 18450 18398 18452 18450
rect 18396 18396 18452 18398
rect 17724 17612 17780 17668
rect 18172 17836 18228 17892
rect 17612 17052 17668 17108
rect 18620 18562 18676 18564
rect 18620 18510 18622 18562
rect 18622 18510 18674 18562
rect 18674 18510 18676 18562
rect 18620 18508 18676 18510
rect 18508 17836 18564 17892
rect 18732 17724 18788 17780
rect 16716 15932 16772 15988
rect 16716 15484 16772 15540
rect 16268 15202 16324 15204
rect 16268 15150 16270 15202
rect 16270 15150 16322 15202
rect 16322 15150 16324 15202
rect 16268 15148 16324 15150
rect 16044 15036 16100 15092
rect 15260 13804 15316 13860
rect 14140 13468 14196 13524
rect 12908 10892 12964 10948
rect 13804 12178 13860 12180
rect 13804 12126 13806 12178
rect 13806 12126 13858 12178
rect 13858 12126 13860 12178
rect 13804 12124 13860 12126
rect 12796 10834 12852 10836
rect 12796 10782 12798 10834
rect 12798 10782 12850 10834
rect 12850 10782 12852 10834
rect 12796 10780 12852 10782
rect 12460 10722 12516 10724
rect 12460 10670 12462 10722
rect 12462 10670 12514 10722
rect 12514 10670 12516 10722
rect 12460 10668 12516 10670
rect 12012 10444 12068 10500
rect 12572 10444 12628 10500
rect 12684 10668 12740 10724
rect 11676 9826 11732 9828
rect 11676 9774 11678 9826
rect 11678 9774 11730 9826
rect 11730 9774 11732 9826
rect 11676 9772 11732 9774
rect 12572 9938 12628 9940
rect 12572 9886 12574 9938
rect 12574 9886 12626 9938
rect 12626 9886 12628 9938
rect 12572 9884 12628 9886
rect 12012 9154 12068 9156
rect 12012 9102 12014 9154
rect 12014 9102 12066 9154
rect 12066 9102 12068 9154
rect 12012 9100 12068 9102
rect 11900 9042 11956 9044
rect 11900 8990 11902 9042
rect 11902 8990 11954 9042
rect 11954 8990 11956 9042
rect 11900 8988 11956 8990
rect 12908 10444 12964 10500
rect 12908 9324 12964 9380
rect 12572 6690 12628 6692
rect 12572 6638 12574 6690
rect 12574 6638 12626 6690
rect 12626 6638 12628 6690
rect 12572 6636 12628 6638
rect 12908 6748 12964 6804
rect 12012 6466 12068 6468
rect 12012 6414 12014 6466
rect 12014 6414 12066 6466
rect 12066 6414 12068 6466
rect 12012 6412 12068 6414
rect 13244 10780 13300 10836
rect 13244 10220 13300 10276
rect 13468 10444 13524 10500
rect 14364 13074 14420 13076
rect 14364 13022 14366 13074
rect 14366 13022 14418 13074
rect 14418 13022 14420 13074
rect 14364 13020 14420 13022
rect 14476 12236 14532 12292
rect 14252 11394 14308 11396
rect 14252 11342 14254 11394
rect 14254 11342 14306 11394
rect 14306 11342 14308 11394
rect 14252 11340 14308 11342
rect 14364 10780 14420 10836
rect 14364 10444 14420 10500
rect 13692 10108 13748 10164
rect 13356 9884 13412 9940
rect 13804 9602 13860 9604
rect 13804 9550 13806 9602
rect 13806 9550 13858 9602
rect 13858 9550 13860 9602
rect 13804 9548 13860 9550
rect 14252 10220 14308 10276
rect 13580 9100 13636 9156
rect 13468 7644 13524 7700
rect 12684 6466 12740 6468
rect 12684 6414 12686 6466
rect 12686 6414 12738 6466
rect 12738 6414 12740 6466
rect 12684 6412 12740 6414
rect 13132 6748 13188 6804
rect 11452 4508 11508 4564
rect 11228 4284 11284 4340
rect 10556 3612 10612 3668
rect 11116 4226 11172 4228
rect 11116 4174 11118 4226
rect 11118 4174 11170 4226
rect 11170 4174 11172 4226
rect 11116 4172 11172 4174
rect 10332 3388 10388 3444
rect 9772 2604 9828 2660
rect 10872 3946 10928 3948
rect 10872 3894 10874 3946
rect 10874 3894 10926 3946
rect 10926 3894 10928 3946
rect 10872 3892 10928 3894
rect 10976 3946 11032 3948
rect 10976 3894 10978 3946
rect 10978 3894 11030 3946
rect 11030 3894 11032 3946
rect 10976 3892 11032 3894
rect 11080 3946 11136 3948
rect 11080 3894 11082 3946
rect 11082 3894 11134 3946
rect 11134 3894 11136 3946
rect 11080 3892 11136 3894
rect 10668 2380 10724 2436
rect 9548 1036 9604 1092
rect 11452 4060 11508 4116
rect 12124 5404 12180 5460
rect 12796 5180 12852 5236
rect 11564 3724 11620 3780
rect 11452 3612 11508 3668
rect 11676 3554 11732 3556
rect 11676 3502 11678 3554
rect 11678 3502 11730 3554
rect 11730 3502 11732 3554
rect 11676 3500 11732 3502
rect 13020 5516 13076 5572
rect 15708 13804 15764 13860
rect 16156 13916 16212 13972
rect 15708 13634 15764 13636
rect 15708 13582 15710 13634
rect 15710 13582 15762 13634
rect 15762 13582 15764 13634
rect 15708 13580 15764 13582
rect 15932 12908 15988 12964
rect 15372 11788 15428 11844
rect 15260 11394 15316 11396
rect 15260 11342 15262 11394
rect 15262 11342 15314 11394
rect 15314 11342 15316 11394
rect 15260 11340 15316 11342
rect 15148 11170 15204 11172
rect 15148 11118 15150 11170
rect 15150 11118 15202 11170
rect 15202 11118 15204 11170
rect 15148 11116 15204 11118
rect 14924 10834 14980 10836
rect 14924 10782 14926 10834
rect 14926 10782 14978 10834
rect 14978 10782 14980 10834
rect 14924 10780 14980 10782
rect 15148 10444 15204 10500
rect 14924 10332 14980 10388
rect 14700 10108 14756 10164
rect 14476 9548 14532 9604
rect 14588 9436 14644 9492
rect 14476 9324 14532 9380
rect 14252 7644 14308 7700
rect 13692 6802 13748 6804
rect 13692 6750 13694 6802
rect 13694 6750 13746 6802
rect 13746 6750 13748 6802
rect 13692 6748 13748 6750
rect 14252 6300 14308 6356
rect 13916 5516 13972 5572
rect 13468 5180 13524 5236
rect 14364 5516 14420 5572
rect 14252 5234 14308 5236
rect 14252 5182 14254 5234
rect 14254 5182 14306 5234
rect 14306 5182 14308 5234
rect 14252 5180 14308 5182
rect 14028 5068 14084 5124
rect 14028 4508 14084 4564
rect 12236 4338 12292 4340
rect 12236 4286 12238 4338
rect 12238 4286 12290 4338
rect 12290 4286 12292 4338
rect 12236 4284 12292 4286
rect 12124 4172 12180 4228
rect 13356 4226 13412 4228
rect 13356 4174 13358 4226
rect 13358 4174 13410 4226
rect 13410 4174 13412 4226
rect 13356 4172 13412 4174
rect 12012 4060 12068 4116
rect 13356 3724 13412 3780
rect 12908 3442 12964 3444
rect 12908 3390 12910 3442
rect 12910 3390 12962 3442
rect 12962 3390 12964 3442
rect 12908 3388 12964 3390
rect 11788 812 11844 868
rect 13580 3724 13636 3780
rect 14588 8204 14644 8260
rect 14588 7698 14644 7700
rect 14588 7646 14590 7698
rect 14590 7646 14642 7698
rect 14642 7646 14644 7698
rect 14588 7644 14644 7646
rect 15484 11340 15540 11396
rect 15484 10332 15540 10388
rect 15596 11228 15652 11284
rect 15372 10108 15428 10164
rect 15708 11170 15764 11172
rect 15708 11118 15710 11170
rect 15710 11118 15762 11170
rect 15762 11118 15764 11170
rect 15708 11116 15764 11118
rect 16156 12402 16212 12404
rect 16156 12350 16158 12402
rect 16158 12350 16210 12402
rect 16210 12350 16212 12402
rect 16156 12348 16212 12350
rect 16156 12124 16212 12180
rect 16828 13970 16884 13972
rect 16828 13918 16830 13970
rect 16830 13918 16882 13970
rect 16882 13918 16884 13970
rect 16828 13916 16884 13918
rect 16716 13580 16772 13636
rect 16716 13132 16772 13188
rect 18284 16882 18340 16884
rect 18284 16830 18286 16882
rect 18286 16830 18338 16882
rect 18338 16830 18340 16882
rect 18284 16828 18340 16830
rect 17164 16210 17220 16212
rect 17164 16158 17166 16210
rect 17166 16158 17218 16210
rect 17218 16158 17220 16210
rect 17164 16156 17220 16158
rect 17388 16156 17444 16212
rect 18172 16268 18228 16324
rect 18508 16716 18564 16772
rect 18732 16268 18788 16324
rect 18508 16156 18564 16212
rect 17948 15986 18004 15988
rect 17948 15934 17950 15986
rect 17950 15934 18002 15986
rect 18002 15934 18004 15986
rect 17948 15932 18004 15934
rect 17836 15874 17892 15876
rect 17836 15822 17838 15874
rect 17838 15822 17890 15874
rect 17890 15822 17892 15874
rect 17836 15820 17892 15822
rect 17836 15260 17892 15316
rect 17836 13746 17892 13748
rect 17836 13694 17838 13746
rect 17838 13694 17890 13746
rect 17890 13694 17892 13746
rect 17836 13692 17892 13694
rect 17724 13580 17780 13636
rect 16492 12178 16548 12180
rect 16492 12126 16494 12178
rect 16494 12126 16546 12178
rect 16546 12126 16548 12178
rect 16492 12124 16548 12126
rect 18060 15484 18116 15540
rect 18060 15148 18116 15204
rect 17724 12460 17780 12516
rect 17948 12796 18004 12852
rect 17052 12402 17108 12404
rect 17052 12350 17054 12402
rect 17054 12350 17106 12402
rect 17106 12350 17108 12402
rect 17052 12348 17108 12350
rect 16156 11340 16212 11396
rect 16716 11282 16772 11284
rect 16716 11230 16718 11282
rect 16718 11230 16770 11282
rect 16770 11230 16772 11282
rect 16716 11228 16772 11230
rect 17724 11282 17780 11284
rect 17724 11230 17726 11282
rect 17726 11230 17778 11282
rect 17778 11230 17780 11282
rect 17724 11228 17780 11230
rect 17276 11170 17332 11172
rect 17276 11118 17278 11170
rect 17278 11118 17330 11170
rect 17330 11118 17332 11170
rect 17276 11116 17332 11118
rect 15932 10834 15988 10836
rect 15932 10782 15934 10834
rect 15934 10782 15986 10834
rect 15986 10782 15988 10834
rect 15932 10780 15988 10782
rect 16604 10332 16660 10388
rect 15036 9938 15092 9940
rect 15036 9886 15038 9938
rect 15038 9886 15090 9938
rect 15090 9886 15092 9938
rect 15036 9884 15092 9886
rect 15148 9436 15204 9492
rect 15260 9548 15316 9604
rect 15932 9548 15988 9604
rect 14924 7644 14980 7700
rect 14924 7308 14980 7364
rect 15260 8258 15316 8260
rect 15260 8206 15262 8258
rect 15262 8206 15314 8258
rect 15314 8206 15316 8258
rect 15260 8204 15316 8206
rect 15820 8034 15876 8036
rect 15820 7982 15822 8034
rect 15822 7982 15874 8034
rect 15874 7982 15876 8034
rect 15820 7980 15876 7982
rect 15372 7698 15428 7700
rect 15372 7646 15374 7698
rect 15374 7646 15426 7698
rect 15426 7646 15428 7698
rect 15372 7644 15428 7646
rect 16268 9602 16324 9604
rect 16268 9550 16270 9602
rect 16270 9550 16322 9602
rect 16322 9550 16324 9602
rect 16268 9548 16324 9550
rect 16716 9436 16772 9492
rect 17052 9996 17108 10052
rect 17052 8988 17108 9044
rect 17836 11170 17892 11172
rect 17836 11118 17838 11170
rect 17838 11118 17890 11170
rect 17890 11118 17892 11170
rect 17836 11116 17892 11118
rect 19292 18508 19348 18564
rect 19180 17890 19236 17892
rect 19180 17838 19182 17890
rect 19182 17838 19234 17890
rect 19234 17838 19236 17890
rect 19180 17836 19236 17838
rect 19068 17724 19124 17780
rect 19292 17052 19348 17108
rect 18956 15932 19012 15988
rect 19068 16940 19124 16996
rect 18844 15484 18900 15540
rect 19516 20076 19572 20132
rect 19628 19346 19684 19348
rect 19628 19294 19630 19346
rect 19630 19294 19682 19346
rect 19682 19294 19684 19346
rect 19628 19292 19684 19294
rect 19740 19234 19796 19236
rect 19740 19182 19742 19234
rect 19742 19182 19794 19234
rect 19794 19182 19796 19234
rect 19740 19180 19796 19182
rect 19628 19010 19684 19012
rect 19628 18958 19630 19010
rect 19630 18958 19682 19010
rect 19682 18958 19684 19010
rect 19628 18956 19684 18958
rect 19516 18620 19572 18676
rect 19740 18732 19796 18788
rect 21084 22316 21140 22372
rect 21196 23212 21252 23268
rect 20532 21978 20588 21980
rect 20532 21926 20534 21978
rect 20534 21926 20586 21978
rect 20586 21926 20588 21978
rect 20532 21924 20588 21926
rect 20636 21978 20692 21980
rect 20636 21926 20638 21978
rect 20638 21926 20690 21978
rect 20690 21926 20692 21978
rect 20636 21924 20692 21926
rect 20740 21978 20796 21980
rect 20740 21926 20742 21978
rect 20742 21926 20794 21978
rect 20794 21926 20796 21978
rect 20740 21924 20796 21926
rect 20748 21420 20804 21476
rect 20636 21362 20692 21364
rect 20636 21310 20638 21362
rect 20638 21310 20690 21362
rect 20690 21310 20692 21362
rect 20636 21308 20692 21310
rect 21644 23212 21700 23268
rect 21308 23154 21364 23156
rect 21308 23102 21310 23154
rect 21310 23102 21362 23154
rect 21362 23102 21364 23154
rect 21308 23100 21364 23102
rect 21420 21698 21476 21700
rect 21420 21646 21422 21698
rect 21422 21646 21474 21698
rect 21474 21646 21476 21698
rect 21420 21644 21476 21646
rect 21532 21586 21588 21588
rect 21532 21534 21534 21586
rect 21534 21534 21586 21586
rect 21586 21534 21588 21586
rect 21532 21532 21588 21534
rect 21644 21420 21700 21476
rect 20412 20860 20468 20916
rect 20860 20690 20916 20692
rect 20860 20638 20862 20690
rect 20862 20638 20914 20690
rect 20914 20638 20916 20690
rect 20860 20636 20916 20638
rect 20532 20410 20588 20412
rect 20532 20358 20534 20410
rect 20534 20358 20586 20410
rect 20586 20358 20588 20410
rect 20532 20356 20588 20358
rect 20636 20410 20692 20412
rect 20636 20358 20638 20410
rect 20638 20358 20690 20410
rect 20690 20358 20692 20410
rect 20636 20356 20692 20358
rect 20740 20410 20796 20412
rect 20740 20358 20742 20410
rect 20742 20358 20794 20410
rect 20794 20358 20796 20410
rect 20740 20356 20796 20358
rect 20076 20188 20132 20244
rect 20860 20242 20916 20244
rect 20860 20190 20862 20242
rect 20862 20190 20914 20242
rect 20914 20190 20916 20242
rect 20860 20188 20916 20190
rect 21644 20412 21700 20468
rect 21868 21644 21924 21700
rect 21868 20914 21924 20916
rect 21868 20862 21870 20914
rect 21870 20862 21922 20914
rect 21922 20862 21924 20914
rect 21868 20860 21924 20862
rect 21756 20188 21812 20244
rect 21532 20076 21588 20132
rect 20972 19404 21028 19460
rect 21308 19404 21364 19460
rect 21532 19234 21588 19236
rect 21532 19182 21534 19234
rect 21534 19182 21586 19234
rect 21586 19182 21588 19234
rect 21532 19180 21588 19182
rect 20188 19122 20244 19124
rect 20188 19070 20190 19122
rect 20190 19070 20242 19122
rect 20242 19070 20244 19122
rect 20188 19068 20244 19070
rect 20860 19068 20916 19124
rect 19740 17948 19796 18004
rect 20412 18956 20468 19012
rect 20188 18620 20244 18676
rect 20076 18562 20132 18564
rect 20076 18510 20078 18562
rect 20078 18510 20130 18562
rect 20130 18510 20132 18562
rect 20076 18508 20132 18510
rect 19964 17724 20020 17780
rect 19628 17276 19684 17332
rect 19404 16716 19460 16772
rect 19852 16940 19908 16996
rect 19292 16604 19348 16660
rect 18732 15314 18788 15316
rect 18732 15262 18734 15314
rect 18734 15262 18786 15314
rect 18786 15262 18788 15314
rect 18732 15260 18788 15262
rect 18284 15148 18340 15204
rect 18956 13970 19012 13972
rect 18956 13918 18958 13970
rect 18958 13918 19010 13970
rect 19010 13918 19012 13970
rect 18956 13916 19012 13918
rect 19068 13746 19124 13748
rect 19068 13694 19070 13746
rect 19070 13694 19122 13746
rect 19122 13694 19124 13746
rect 19068 13692 19124 13694
rect 18172 13020 18228 13076
rect 18844 13020 18900 13076
rect 18396 12962 18452 12964
rect 18396 12910 18398 12962
rect 18398 12910 18450 12962
rect 18450 12910 18452 12962
rect 18396 12908 18452 12910
rect 18508 12850 18564 12852
rect 18508 12798 18510 12850
rect 18510 12798 18562 12850
rect 18562 12798 18564 12850
rect 18508 12796 18564 12798
rect 18732 12850 18788 12852
rect 18732 12798 18734 12850
rect 18734 12798 18786 12850
rect 18786 12798 18788 12850
rect 18732 12796 18788 12798
rect 18284 12402 18340 12404
rect 18284 12350 18286 12402
rect 18286 12350 18338 12402
rect 18338 12350 18340 12402
rect 18284 12348 18340 12350
rect 18172 12124 18228 12180
rect 18732 12124 18788 12180
rect 18620 11506 18676 11508
rect 18620 11454 18622 11506
rect 18622 11454 18674 11506
rect 18674 11454 18676 11506
rect 18620 11452 18676 11454
rect 18172 10722 18228 10724
rect 18172 10670 18174 10722
rect 18174 10670 18226 10722
rect 18226 10670 18228 10722
rect 18172 10668 18228 10670
rect 17164 10220 17220 10276
rect 15932 7644 15988 7700
rect 16156 8428 16212 8484
rect 18172 9996 18228 10052
rect 18396 9996 18452 10052
rect 17388 9884 17444 9940
rect 18732 10332 18788 10388
rect 19628 15986 19684 15988
rect 19628 15934 19630 15986
rect 19630 15934 19682 15986
rect 19682 15934 19684 15986
rect 19628 15932 19684 15934
rect 19404 15538 19460 15540
rect 19404 15486 19406 15538
rect 19406 15486 19458 15538
rect 19458 15486 19460 15538
rect 19404 15484 19460 15486
rect 19516 15314 19572 15316
rect 19516 15262 19518 15314
rect 19518 15262 19570 15314
rect 19570 15262 19572 15314
rect 19516 15260 19572 15262
rect 19740 15148 19796 15204
rect 23100 25004 23156 25060
rect 23548 25228 23604 25284
rect 22316 23714 22372 23716
rect 22316 23662 22318 23714
rect 22318 23662 22370 23714
rect 22370 23662 22372 23714
rect 22316 23660 22372 23662
rect 22092 21698 22148 21700
rect 22092 21646 22094 21698
rect 22094 21646 22146 21698
rect 22146 21646 22148 21698
rect 22092 21644 22148 21646
rect 22316 21420 22372 21476
rect 22092 20802 22148 20804
rect 22092 20750 22094 20802
rect 22094 20750 22146 20802
rect 22146 20750 22148 20802
rect 22092 20748 22148 20750
rect 23324 24780 23380 24836
rect 22988 24556 23044 24612
rect 23212 24556 23268 24612
rect 22876 23996 22932 24052
rect 22988 24108 23044 24164
rect 23100 23938 23156 23940
rect 23100 23886 23102 23938
rect 23102 23886 23154 23938
rect 23154 23886 23156 23938
rect 23100 23884 23156 23886
rect 22988 23714 23044 23716
rect 22988 23662 22990 23714
rect 22990 23662 23042 23714
rect 23042 23662 23044 23714
rect 22988 23660 23044 23662
rect 24332 27074 24388 27076
rect 24332 27022 24334 27074
rect 24334 27022 24386 27074
rect 24386 27022 24388 27074
rect 24332 27020 24388 27022
rect 24892 27804 24948 27860
rect 24556 26908 24612 26964
rect 24780 27132 24836 27188
rect 24780 26962 24836 26964
rect 24780 26910 24782 26962
rect 24782 26910 24834 26962
rect 24834 26910 24836 26962
rect 24780 26908 24836 26910
rect 24108 26178 24164 26180
rect 24108 26126 24110 26178
rect 24110 26126 24162 26178
rect 24162 26126 24164 26178
rect 24108 26124 24164 26126
rect 24892 25452 24948 25508
rect 24444 24834 24500 24836
rect 24444 24782 24446 24834
rect 24446 24782 24498 24834
rect 24498 24782 24500 24834
rect 24444 24780 24500 24782
rect 23996 24610 24052 24612
rect 23996 24558 23998 24610
rect 23998 24558 24050 24610
rect 24050 24558 24052 24610
rect 23996 24556 24052 24558
rect 24892 24780 24948 24836
rect 24444 24108 24500 24164
rect 23548 23660 23604 23716
rect 24444 23714 24500 23716
rect 24444 23662 24446 23714
rect 24446 23662 24498 23714
rect 24498 23662 24500 23714
rect 24444 23660 24500 23662
rect 23548 23042 23604 23044
rect 23548 22990 23550 23042
rect 23550 22990 23602 23042
rect 23602 22990 23604 23042
rect 23548 22988 23604 22990
rect 23660 21698 23716 21700
rect 23660 21646 23662 21698
rect 23662 21646 23714 21698
rect 23714 21646 23716 21698
rect 23660 21644 23716 21646
rect 23100 21474 23156 21476
rect 23100 21422 23102 21474
rect 23102 21422 23154 21474
rect 23154 21422 23156 21474
rect 23100 21420 23156 21422
rect 22988 20972 23044 21028
rect 23548 20972 23604 21028
rect 24892 23826 24948 23828
rect 24892 23774 24894 23826
rect 24894 23774 24946 23826
rect 24946 23774 24948 23826
rect 24892 23772 24948 23774
rect 24108 22988 24164 23044
rect 24444 21868 24500 21924
rect 23660 20748 23716 20804
rect 24220 20748 24276 20804
rect 22540 20188 22596 20244
rect 24556 20412 24612 20468
rect 24780 22258 24836 22260
rect 24780 22206 24782 22258
rect 24782 22206 24834 22258
rect 24834 22206 24836 22258
rect 24780 22204 24836 22206
rect 24780 20972 24836 21028
rect 24892 21586 24948 21588
rect 24892 21534 24894 21586
rect 24894 21534 24946 21586
rect 24946 21534 24948 21586
rect 24892 21532 24948 21534
rect 24668 20076 24724 20132
rect 22204 19740 22260 19796
rect 23548 19964 23604 20020
rect 22316 19404 22372 19460
rect 22652 19404 22708 19460
rect 22204 19180 22260 19236
rect 21980 19068 22036 19124
rect 24332 20018 24388 20020
rect 24332 19966 24334 20018
rect 24334 19966 24386 20018
rect 24386 19966 24388 20018
rect 24332 19964 24388 19966
rect 23436 19234 23492 19236
rect 23436 19182 23438 19234
rect 23438 19182 23490 19234
rect 23490 19182 23492 19234
rect 23436 19180 23492 19182
rect 22764 19068 22820 19124
rect 24108 19068 24164 19124
rect 20532 18842 20588 18844
rect 20532 18790 20534 18842
rect 20534 18790 20586 18842
rect 20586 18790 20588 18842
rect 20532 18788 20588 18790
rect 20636 18842 20692 18844
rect 20636 18790 20638 18842
rect 20638 18790 20690 18842
rect 20690 18790 20692 18842
rect 20636 18788 20692 18790
rect 20740 18842 20796 18844
rect 20740 18790 20742 18842
rect 20742 18790 20794 18842
rect 20794 18790 20796 18842
rect 20740 18788 20796 18790
rect 20412 17836 20468 17892
rect 20188 17276 20244 17332
rect 20532 17274 20588 17276
rect 20532 17222 20534 17274
rect 20534 17222 20586 17274
rect 20586 17222 20588 17274
rect 20532 17220 20588 17222
rect 20636 17274 20692 17276
rect 20636 17222 20638 17274
rect 20638 17222 20690 17274
rect 20690 17222 20692 17274
rect 20636 17220 20692 17222
rect 20740 17274 20796 17276
rect 20740 17222 20742 17274
rect 20742 17222 20794 17274
rect 20794 17222 20796 17274
rect 20740 17220 20796 17222
rect 20188 17106 20244 17108
rect 20188 17054 20190 17106
rect 20190 17054 20242 17106
rect 20242 17054 20244 17106
rect 20188 17052 20244 17054
rect 20412 16716 20468 16772
rect 20636 16770 20692 16772
rect 20636 16718 20638 16770
rect 20638 16718 20690 16770
rect 20690 16718 20692 16770
rect 20636 16716 20692 16718
rect 20300 15986 20356 15988
rect 20300 15934 20302 15986
rect 20302 15934 20354 15986
rect 20354 15934 20356 15986
rect 20300 15932 20356 15934
rect 20300 15148 20356 15204
rect 21196 18956 21252 19012
rect 21196 18620 21252 18676
rect 23436 18674 23492 18676
rect 23436 18622 23438 18674
rect 23438 18622 23490 18674
rect 23490 18622 23492 18674
rect 23436 18620 23492 18622
rect 24108 18620 24164 18676
rect 22204 18508 22260 18564
rect 20972 18284 21028 18340
rect 23548 18562 23604 18564
rect 23548 18510 23550 18562
rect 23550 18510 23602 18562
rect 23602 18510 23604 18562
rect 24780 19404 24836 19460
rect 23548 18508 23604 18510
rect 21868 18284 21924 18340
rect 21420 18172 21476 18228
rect 21868 16940 21924 16996
rect 21532 16882 21588 16884
rect 21532 16830 21534 16882
rect 21534 16830 21586 16882
rect 21586 16830 21588 16882
rect 21532 16828 21588 16830
rect 21980 16828 22036 16884
rect 23324 18284 23380 18340
rect 25116 29932 25172 29988
rect 26908 31164 26964 31220
rect 25340 30268 25396 30324
rect 26348 30940 26404 30996
rect 26012 30322 26068 30324
rect 26012 30270 26014 30322
rect 26014 30270 26066 30322
rect 26066 30270 26068 30322
rect 26012 30268 26068 30270
rect 26908 29708 26964 29764
rect 26908 29538 26964 29540
rect 26908 29486 26910 29538
rect 26910 29486 26962 29538
rect 26962 29486 26964 29538
rect 26908 29484 26964 29486
rect 25564 28700 25620 28756
rect 26348 29314 26404 29316
rect 26348 29262 26350 29314
rect 26350 29262 26402 29314
rect 26402 29262 26404 29314
rect 26348 29260 26404 29262
rect 27468 32562 27524 32564
rect 27468 32510 27470 32562
rect 27470 32510 27522 32562
rect 27522 32510 27524 32562
rect 27468 32508 27524 32510
rect 28476 33122 28532 33124
rect 28476 33070 28478 33122
rect 28478 33070 28530 33122
rect 28530 33070 28532 33122
rect 28476 33068 28532 33070
rect 27580 32284 27636 32340
rect 27244 30994 27300 30996
rect 27244 30942 27246 30994
rect 27246 30942 27298 30994
rect 27298 30942 27300 30994
rect 27244 30940 27300 30942
rect 27692 31500 27748 31556
rect 27804 31164 27860 31220
rect 25900 28530 25956 28532
rect 25900 28478 25902 28530
rect 25902 28478 25954 28530
rect 25954 28478 25956 28530
rect 25900 28476 25956 28478
rect 26796 28476 26852 28532
rect 25788 28418 25844 28420
rect 25788 28366 25790 28418
rect 25790 28366 25842 28418
rect 25842 28366 25844 28418
rect 25788 28364 25844 28366
rect 25228 28252 25284 28308
rect 26012 27804 26068 27860
rect 25564 27746 25620 27748
rect 25564 27694 25566 27746
rect 25566 27694 25618 27746
rect 25618 27694 25620 27746
rect 25564 27692 25620 27694
rect 25228 27074 25284 27076
rect 25228 27022 25230 27074
rect 25230 27022 25282 27074
rect 25282 27022 25284 27074
rect 25228 27020 25284 27022
rect 26572 27858 26628 27860
rect 26572 27806 26574 27858
rect 26574 27806 26626 27858
rect 26626 27806 26628 27858
rect 26572 27804 26628 27806
rect 26012 27020 26068 27076
rect 27020 28418 27076 28420
rect 27020 28366 27022 28418
rect 27022 28366 27074 28418
rect 27074 28366 27076 28418
rect 27020 28364 27076 28366
rect 26124 26908 26180 26964
rect 25564 26514 25620 26516
rect 25564 26462 25566 26514
rect 25566 26462 25618 26514
rect 25618 26462 25620 26514
rect 25564 26460 25620 26462
rect 25676 25900 25732 25956
rect 25676 25618 25732 25620
rect 25676 25566 25678 25618
rect 25678 25566 25730 25618
rect 25730 25566 25732 25618
rect 25676 25564 25732 25566
rect 25228 25340 25284 25396
rect 26236 25394 26292 25396
rect 26236 25342 26238 25394
rect 26238 25342 26290 25394
rect 26290 25342 26292 25394
rect 26236 25340 26292 25342
rect 26684 26962 26740 26964
rect 26684 26910 26686 26962
rect 26686 26910 26738 26962
rect 26738 26910 26740 26962
rect 26684 26908 26740 26910
rect 26908 26850 26964 26852
rect 26908 26798 26910 26850
rect 26910 26798 26962 26850
rect 26962 26798 26964 26850
rect 26908 26796 26964 26798
rect 26796 26572 26852 26628
rect 27356 29708 27412 29764
rect 27468 29484 27524 29540
rect 28588 29708 28644 29764
rect 27356 28924 27412 28980
rect 30192 33738 30248 33740
rect 30192 33686 30194 33738
rect 30194 33686 30246 33738
rect 30246 33686 30248 33738
rect 30192 33684 30248 33686
rect 30296 33738 30352 33740
rect 30296 33686 30298 33738
rect 30298 33686 30350 33738
rect 30350 33686 30352 33738
rect 30296 33684 30352 33686
rect 30400 33738 30456 33740
rect 30400 33686 30402 33738
rect 30402 33686 30454 33738
rect 30454 33686 30456 33738
rect 30400 33684 30456 33686
rect 30716 34412 30772 34468
rect 32060 35868 32116 35924
rect 32396 35756 32452 35812
rect 31500 34412 31556 34468
rect 32732 35868 32788 35924
rect 40236 37996 40292 38052
rect 35196 36540 35252 36596
rect 34972 36428 35028 36484
rect 34860 36316 34916 36372
rect 34860 35810 34916 35812
rect 34860 35758 34862 35810
rect 34862 35758 34914 35810
rect 34914 35758 34916 35810
rect 34860 35756 34916 35758
rect 32844 35698 32900 35700
rect 32844 35646 32846 35698
rect 32846 35646 32898 35698
rect 32898 35646 32900 35698
rect 32844 35644 32900 35646
rect 33628 35698 33684 35700
rect 33628 35646 33630 35698
rect 33630 35646 33682 35698
rect 33682 35646 33684 35698
rect 35644 36482 35700 36484
rect 35644 36430 35646 36482
rect 35646 36430 35698 36482
rect 35698 36430 35700 36482
rect 35644 36428 35700 36430
rect 35868 36482 35924 36484
rect 35868 36430 35870 36482
rect 35870 36430 35922 36482
rect 35922 36430 35924 36482
rect 35868 36428 35924 36430
rect 36092 36370 36148 36372
rect 36092 36318 36094 36370
rect 36094 36318 36146 36370
rect 36146 36318 36148 36370
rect 36092 36316 36148 36318
rect 34972 35868 35028 35924
rect 33628 35644 33684 35646
rect 34748 34914 34804 34916
rect 34748 34862 34750 34914
rect 34750 34862 34802 34914
rect 34802 34862 34804 34914
rect 34748 34860 34804 34862
rect 35532 35474 35588 35476
rect 35532 35422 35534 35474
rect 35534 35422 35586 35474
rect 35586 35422 35588 35474
rect 35532 35420 35588 35422
rect 35084 34748 35140 34804
rect 33852 34354 33908 34356
rect 33852 34302 33854 34354
rect 33854 34302 33906 34354
rect 33906 34302 33908 34354
rect 33852 34300 33908 34302
rect 32620 34188 32676 34244
rect 32060 34076 32116 34132
rect 31612 33906 31668 33908
rect 31612 33854 31614 33906
rect 31614 33854 31666 33906
rect 31666 33854 31668 33906
rect 31612 33852 31668 33854
rect 32844 34130 32900 34132
rect 32844 34078 32846 34130
rect 32846 34078 32898 34130
rect 32898 34078 32900 34130
rect 32844 34076 32900 34078
rect 29932 33292 29988 33348
rect 29820 33068 29876 33124
rect 31836 33068 31892 33124
rect 28924 32562 28980 32564
rect 28924 32510 28926 32562
rect 28926 32510 28978 32562
rect 28978 32510 28980 32562
rect 28924 32508 28980 32510
rect 29148 32338 29204 32340
rect 29148 32286 29150 32338
rect 29150 32286 29202 32338
rect 29202 32286 29204 32338
rect 29148 32284 29204 32286
rect 30192 32170 30248 32172
rect 30192 32118 30194 32170
rect 30194 32118 30246 32170
rect 30246 32118 30248 32170
rect 30192 32116 30248 32118
rect 30296 32170 30352 32172
rect 30296 32118 30298 32170
rect 30298 32118 30350 32170
rect 30350 32118 30352 32170
rect 30296 32116 30352 32118
rect 30400 32170 30456 32172
rect 30400 32118 30402 32170
rect 30402 32118 30454 32170
rect 30454 32118 30456 32170
rect 30400 32116 30456 32118
rect 31388 32450 31444 32452
rect 31388 32398 31390 32450
rect 31390 32398 31442 32450
rect 31442 32398 31444 32450
rect 31388 32396 31444 32398
rect 31164 31948 31220 32004
rect 31612 31948 31668 32004
rect 29596 30940 29652 30996
rect 30492 30994 30548 30996
rect 30492 30942 30494 30994
rect 30494 30942 30546 30994
rect 30546 30942 30548 30994
rect 30492 30940 30548 30942
rect 29372 30156 29428 30212
rect 28812 29986 28868 29988
rect 28812 29934 28814 29986
rect 28814 29934 28866 29986
rect 28866 29934 28868 29986
rect 28812 29932 28868 29934
rect 28812 29372 28868 29428
rect 28476 28642 28532 28644
rect 28476 28590 28478 28642
rect 28478 28590 28530 28642
rect 28530 28590 28532 28642
rect 28476 28588 28532 28590
rect 28140 28476 28196 28532
rect 27580 28364 27636 28420
rect 27356 27692 27412 27748
rect 27916 27916 27972 27972
rect 28028 28364 28084 28420
rect 27692 27692 27748 27748
rect 27020 26460 27076 26516
rect 26796 25564 26852 25620
rect 26684 25394 26740 25396
rect 26684 25342 26686 25394
rect 26686 25342 26738 25394
rect 26738 25342 26740 25394
rect 26684 25340 26740 25342
rect 26908 25900 26964 25956
rect 27356 25900 27412 25956
rect 27692 25900 27748 25956
rect 27580 25452 27636 25508
rect 26124 24834 26180 24836
rect 26124 24782 26126 24834
rect 26126 24782 26178 24834
rect 26178 24782 26180 24834
rect 26124 24780 26180 24782
rect 25676 24668 25732 24724
rect 25564 24610 25620 24612
rect 25564 24558 25566 24610
rect 25566 24558 25618 24610
rect 25618 24558 25620 24610
rect 25564 24556 25620 24558
rect 25452 23826 25508 23828
rect 25452 23774 25454 23826
rect 25454 23774 25506 23826
rect 25506 23774 25508 23826
rect 25452 23772 25508 23774
rect 26012 24050 26068 24052
rect 26012 23998 26014 24050
rect 26014 23998 26066 24050
rect 26066 23998 26068 24050
rect 26012 23996 26068 23998
rect 25676 23772 25732 23828
rect 25228 23212 25284 23268
rect 27132 25340 27188 25396
rect 26348 24722 26404 24724
rect 26348 24670 26350 24722
rect 26350 24670 26402 24722
rect 26402 24670 26404 24722
rect 26348 24668 26404 24670
rect 26572 24556 26628 24612
rect 25228 22258 25284 22260
rect 25228 22206 25230 22258
rect 25230 22206 25282 22258
rect 25282 22206 25284 22258
rect 25228 22204 25284 22206
rect 25900 23714 25956 23716
rect 25900 23662 25902 23714
rect 25902 23662 25954 23714
rect 25954 23662 25956 23714
rect 25900 23660 25956 23662
rect 25900 23266 25956 23268
rect 25900 23214 25902 23266
rect 25902 23214 25954 23266
rect 25954 23214 25956 23266
rect 25900 23212 25956 23214
rect 25676 21868 25732 21924
rect 26572 23436 26628 23492
rect 26572 23266 26628 23268
rect 26572 23214 26574 23266
rect 26574 23214 26626 23266
rect 26626 23214 26628 23266
rect 26572 23212 26628 23214
rect 26908 23714 26964 23716
rect 26908 23662 26910 23714
rect 26910 23662 26962 23714
rect 26962 23662 26964 23714
rect 26908 23660 26964 23662
rect 26348 22258 26404 22260
rect 26348 22206 26350 22258
rect 26350 22206 26402 22258
rect 26402 22206 26404 22258
rect 26348 22204 26404 22206
rect 26460 21868 26516 21924
rect 25116 20748 25172 20804
rect 25788 20972 25844 21028
rect 25564 20690 25620 20692
rect 25564 20638 25566 20690
rect 25566 20638 25618 20690
rect 25618 20638 25620 20690
rect 25564 20636 25620 20638
rect 25116 20578 25172 20580
rect 25116 20526 25118 20578
rect 25118 20526 25170 20578
rect 25170 20526 25172 20578
rect 25116 20524 25172 20526
rect 24892 18450 24948 18452
rect 24892 18398 24894 18450
rect 24894 18398 24946 18450
rect 24946 18398 24948 18450
rect 24892 18396 24948 18398
rect 25004 19234 25060 19236
rect 25004 19182 25006 19234
rect 25006 19182 25058 19234
rect 25058 19182 25060 19234
rect 25004 19180 25060 19182
rect 22764 18172 22820 18228
rect 22204 16940 22260 16996
rect 21644 16098 21700 16100
rect 21644 16046 21646 16098
rect 21646 16046 21698 16098
rect 21698 16046 21700 16098
rect 21644 16044 21700 16046
rect 20636 15874 20692 15876
rect 20636 15822 20638 15874
rect 20638 15822 20690 15874
rect 20690 15822 20692 15874
rect 20636 15820 20692 15822
rect 20532 15706 20588 15708
rect 20532 15654 20534 15706
rect 20534 15654 20586 15706
rect 20586 15654 20588 15706
rect 20532 15652 20588 15654
rect 20636 15706 20692 15708
rect 20636 15654 20638 15706
rect 20638 15654 20690 15706
rect 20690 15654 20692 15706
rect 20636 15652 20692 15654
rect 20740 15706 20796 15708
rect 20740 15654 20742 15706
rect 20742 15654 20794 15706
rect 20794 15654 20796 15706
rect 20740 15652 20796 15654
rect 21084 15484 21140 15540
rect 21084 15260 21140 15316
rect 21308 15314 21364 15316
rect 21308 15262 21310 15314
rect 21310 15262 21362 15314
rect 21362 15262 21364 15314
rect 21308 15260 21364 15262
rect 19740 13468 19796 13524
rect 19292 13020 19348 13076
rect 19404 12962 19460 12964
rect 19404 12910 19406 12962
rect 19406 12910 19458 12962
rect 19458 12910 19460 12962
rect 19404 12908 19460 12910
rect 19180 12796 19236 12852
rect 19292 12738 19348 12740
rect 19292 12686 19294 12738
rect 19294 12686 19346 12738
rect 19346 12686 19348 12738
rect 19292 12684 19348 12686
rect 20532 14138 20588 14140
rect 20532 14086 20534 14138
rect 20534 14086 20586 14138
rect 20586 14086 20588 14138
rect 20532 14084 20588 14086
rect 20636 14138 20692 14140
rect 20636 14086 20638 14138
rect 20638 14086 20690 14138
rect 20690 14086 20692 14138
rect 20636 14084 20692 14086
rect 20740 14138 20796 14140
rect 20740 14086 20742 14138
rect 20742 14086 20794 14138
rect 20794 14086 20796 14138
rect 20740 14084 20796 14086
rect 20972 13746 21028 13748
rect 20972 13694 20974 13746
rect 20974 13694 21026 13746
rect 21026 13694 21028 13746
rect 20972 13692 21028 13694
rect 20300 12850 20356 12852
rect 20300 12798 20302 12850
rect 20302 12798 20354 12850
rect 20354 12798 20356 12850
rect 20300 12796 20356 12798
rect 19964 12684 20020 12740
rect 19068 12402 19124 12404
rect 19068 12350 19070 12402
rect 19070 12350 19122 12402
rect 19122 12350 19124 12402
rect 19068 12348 19124 12350
rect 19292 12402 19348 12404
rect 19292 12350 19294 12402
rect 19294 12350 19346 12402
rect 19346 12350 19348 12402
rect 19292 12348 19348 12350
rect 18956 11900 19012 11956
rect 19964 12124 20020 12180
rect 19068 11228 19124 11284
rect 19068 10444 19124 10500
rect 19292 11564 19348 11620
rect 17276 9548 17332 9604
rect 17388 9436 17444 9492
rect 15820 7308 15876 7364
rect 15596 6690 15652 6692
rect 15596 6638 15598 6690
rect 15598 6638 15650 6690
rect 15650 6638 15652 6690
rect 15596 6636 15652 6638
rect 16044 6636 16100 6692
rect 14812 6412 14868 6468
rect 14700 5794 14756 5796
rect 14700 5742 14702 5794
rect 14702 5742 14754 5794
rect 14754 5742 14756 5794
rect 14700 5740 14756 5742
rect 14924 5516 14980 5572
rect 15036 5068 15092 5124
rect 16604 8258 16660 8260
rect 16604 8206 16606 8258
rect 16606 8206 16658 8258
rect 16658 8206 16660 8258
rect 16604 8204 16660 8206
rect 17164 8258 17220 8260
rect 17164 8206 17166 8258
rect 17166 8206 17218 8258
rect 17218 8206 17220 8258
rect 17164 8204 17220 8206
rect 16604 7644 16660 7700
rect 16268 6636 16324 6692
rect 16268 5180 16324 5236
rect 14924 4172 14980 4228
rect 14924 3500 14980 3556
rect 15036 3724 15092 3780
rect 15372 4060 15428 4116
rect 15036 3442 15092 3444
rect 15036 3390 15038 3442
rect 15038 3390 15090 3442
rect 15090 3390 15092 3442
rect 15036 3388 15092 3390
rect 15820 5068 15876 5124
rect 16492 5852 16548 5908
rect 16940 5516 16996 5572
rect 16380 5068 16436 5124
rect 16716 5180 16772 5236
rect 16380 4562 16436 4564
rect 16380 4510 16382 4562
rect 16382 4510 16434 4562
rect 16434 4510 16436 4562
rect 16380 4508 16436 4510
rect 15708 3554 15764 3556
rect 15708 3502 15710 3554
rect 15710 3502 15762 3554
rect 15762 3502 15764 3554
rect 15708 3500 15764 3502
rect 16268 3330 16324 3332
rect 16268 3278 16270 3330
rect 16270 3278 16322 3330
rect 16322 3278 16324 3330
rect 16268 3276 16324 3278
rect 14700 2156 14756 2212
rect 16604 5010 16660 5012
rect 16604 4958 16606 5010
rect 16606 4958 16658 5010
rect 16658 4958 16660 5010
rect 16604 4956 16660 4958
rect 16492 1260 16548 1316
rect 17052 5122 17108 5124
rect 17052 5070 17054 5122
rect 17054 5070 17106 5122
rect 17106 5070 17108 5122
rect 17052 5068 17108 5070
rect 17948 9324 18004 9380
rect 17612 5852 17668 5908
rect 17500 5122 17556 5124
rect 17500 5070 17502 5122
rect 17502 5070 17554 5122
rect 17554 5070 17556 5122
rect 17500 5068 17556 5070
rect 18172 9212 18228 9268
rect 18060 9042 18116 9044
rect 18060 8990 18062 9042
rect 18062 8990 18114 9042
rect 18114 8990 18116 9042
rect 18060 8988 18116 8990
rect 18284 9100 18340 9156
rect 18396 9436 18452 9492
rect 18620 8876 18676 8932
rect 18620 8204 18676 8260
rect 18508 7980 18564 8036
rect 18284 5906 18340 5908
rect 18284 5854 18286 5906
rect 18286 5854 18338 5906
rect 18338 5854 18340 5906
rect 18284 5852 18340 5854
rect 17724 5068 17780 5124
rect 17164 4956 17220 5012
rect 17500 3554 17556 3556
rect 17500 3502 17502 3554
rect 17502 3502 17554 3554
rect 17554 3502 17556 3554
rect 17500 3500 17556 3502
rect 14476 924 14532 980
rect 17500 1596 17556 1652
rect 18284 4396 18340 4452
rect 18508 6018 18564 6020
rect 18508 5966 18510 6018
rect 18510 5966 18562 6018
rect 18562 5966 18564 6018
rect 18508 5964 18564 5966
rect 18844 9938 18900 9940
rect 18844 9886 18846 9938
rect 18846 9886 18898 9938
rect 18898 9886 18900 9938
rect 18844 9884 18900 9886
rect 19628 10668 19684 10724
rect 19404 10332 19460 10388
rect 19516 10220 19572 10276
rect 19516 10050 19572 10052
rect 19516 9998 19518 10050
rect 19518 9998 19570 10050
rect 19570 9998 19572 10050
rect 19516 9996 19572 9998
rect 20188 12738 20244 12740
rect 20188 12686 20190 12738
rect 20190 12686 20242 12738
rect 20242 12686 20244 12738
rect 20188 12684 20244 12686
rect 20532 12570 20588 12572
rect 20532 12518 20534 12570
rect 20534 12518 20586 12570
rect 20586 12518 20588 12570
rect 20532 12516 20588 12518
rect 20636 12570 20692 12572
rect 20636 12518 20638 12570
rect 20638 12518 20690 12570
rect 20690 12518 20692 12570
rect 20636 12516 20692 12518
rect 20740 12570 20796 12572
rect 20740 12518 20742 12570
rect 20742 12518 20794 12570
rect 20794 12518 20796 12570
rect 20740 12516 20796 12518
rect 20860 12348 20916 12404
rect 21084 12402 21140 12404
rect 21084 12350 21086 12402
rect 21086 12350 21138 12402
rect 21138 12350 21140 12402
rect 21084 12348 21140 12350
rect 20076 11900 20132 11956
rect 20524 12124 20580 12180
rect 20524 11954 20580 11956
rect 20524 11902 20526 11954
rect 20526 11902 20578 11954
rect 20578 11902 20580 11954
rect 20524 11900 20580 11902
rect 20748 11900 20804 11956
rect 20860 12124 20916 12180
rect 21644 15538 21700 15540
rect 21644 15486 21646 15538
rect 21646 15486 21698 15538
rect 21698 15486 21700 15538
rect 21644 15484 21700 15486
rect 21868 15484 21924 15540
rect 22204 15148 22260 15204
rect 22316 16044 22372 16100
rect 21644 12850 21700 12852
rect 21644 12798 21646 12850
rect 21646 12798 21698 12850
rect 21698 12798 21700 12850
rect 21644 12796 21700 12798
rect 21084 11900 21140 11956
rect 21308 12012 21364 12068
rect 20532 11002 20588 11004
rect 20532 10950 20534 11002
rect 20534 10950 20586 11002
rect 20586 10950 20588 11002
rect 20532 10948 20588 10950
rect 20636 11002 20692 11004
rect 20636 10950 20638 11002
rect 20638 10950 20690 11002
rect 20690 10950 20692 11002
rect 20636 10948 20692 10950
rect 20740 11002 20796 11004
rect 20740 10950 20742 11002
rect 20742 10950 20794 11002
rect 20794 10950 20796 11002
rect 20740 10948 20796 10950
rect 20188 9996 20244 10052
rect 20300 10220 20356 10276
rect 19292 9154 19348 9156
rect 19292 9102 19294 9154
rect 19294 9102 19346 9154
rect 19346 9102 19348 9154
rect 19292 9100 19348 9102
rect 19516 9212 19572 9268
rect 21196 9996 21252 10052
rect 19068 8146 19124 8148
rect 19068 8094 19070 8146
rect 19070 8094 19122 8146
rect 19122 8094 19124 8146
rect 19068 8092 19124 8094
rect 20076 8370 20132 8372
rect 20076 8318 20078 8370
rect 20078 8318 20130 8370
rect 20130 8318 20132 8370
rect 20076 8316 20132 8318
rect 20188 8146 20244 8148
rect 20188 8094 20190 8146
rect 20190 8094 20242 8146
rect 20242 8094 20244 8146
rect 20188 8092 20244 8094
rect 19964 8034 20020 8036
rect 19964 7982 19966 8034
rect 19966 7982 20018 8034
rect 20018 7982 20020 8034
rect 19964 7980 20020 7982
rect 20532 9434 20588 9436
rect 20532 9382 20534 9434
rect 20534 9382 20586 9434
rect 20586 9382 20588 9434
rect 20532 9380 20588 9382
rect 20636 9434 20692 9436
rect 20636 9382 20638 9434
rect 20638 9382 20690 9434
rect 20690 9382 20692 9434
rect 20636 9380 20692 9382
rect 20740 9434 20796 9436
rect 20740 9382 20742 9434
rect 20742 9382 20794 9434
rect 20794 9382 20796 9434
rect 20740 9380 20796 9382
rect 20524 9212 20580 9268
rect 20524 8540 20580 8596
rect 20972 8930 21028 8932
rect 20972 8878 20974 8930
rect 20974 8878 21026 8930
rect 21026 8878 21028 8930
rect 20972 8876 21028 8878
rect 20532 7866 20588 7868
rect 20532 7814 20534 7866
rect 20534 7814 20586 7866
rect 20586 7814 20588 7866
rect 20532 7812 20588 7814
rect 20636 7866 20692 7868
rect 20636 7814 20638 7866
rect 20638 7814 20690 7866
rect 20690 7814 20692 7866
rect 20636 7812 20692 7814
rect 20740 7866 20796 7868
rect 20740 7814 20742 7866
rect 20742 7814 20794 7866
rect 20794 7814 20796 7866
rect 20740 7812 20796 7814
rect 19516 5964 19572 6020
rect 18844 5516 18900 5572
rect 18844 5292 18900 5348
rect 18732 5068 18788 5124
rect 18508 5010 18564 5012
rect 18508 4958 18510 5010
rect 18510 4958 18562 5010
rect 18562 4958 18564 5010
rect 18508 4956 18564 4958
rect 18956 4732 19012 4788
rect 19180 5122 19236 5124
rect 19180 5070 19182 5122
rect 19182 5070 19234 5122
rect 19234 5070 19236 5122
rect 19180 5068 19236 5070
rect 19068 4956 19124 5012
rect 18396 3612 18452 3668
rect 17948 3554 18004 3556
rect 17948 3502 17950 3554
rect 17950 3502 18002 3554
rect 18002 3502 18004 3554
rect 17948 3500 18004 3502
rect 18844 3554 18900 3556
rect 18844 3502 18846 3554
rect 18846 3502 18898 3554
rect 18898 3502 18900 3554
rect 18844 3500 18900 3502
rect 19964 5180 20020 5236
rect 19740 4956 19796 5012
rect 19740 4508 19796 4564
rect 19964 4898 20020 4900
rect 19964 4846 19966 4898
rect 19966 4846 20018 4898
rect 20018 4846 20020 4898
rect 19964 4844 20020 4846
rect 20076 4508 20132 4564
rect 19516 3836 19572 3892
rect 19068 2716 19124 2772
rect 19740 3500 19796 3556
rect 20412 7308 20468 7364
rect 21532 12066 21588 12068
rect 21532 12014 21534 12066
rect 21534 12014 21586 12066
rect 21586 12014 21588 12066
rect 21532 12012 21588 12014
rect 21644 11506 21700 11508
rect 21644 11454 21646 11506
rect 21646 11454 21698 11506
rect 21698 11454 21700 11506
rect 21644 11452 21700 11454
rect 22092 12850 22148 12852
rect 22092 12798 22094 12850
rect 22094 12798 22146 12850
rect 22146 12798 22148 12850
rect 22092 12796 22148 12798
rect 21980 12348 22036 12404
rect 22204 12348 22260 12404
rect 22652 16098 22708 16100
rect 22652 16046 22654 16098
rect 22654 16046 22706 16098
rect 22706 16046 22708 16098
rect 22652 16044 22708 16046
rect 23436 16156 23492 16212
rect 22876 15484 22932 15540
rect 23324 16044 23380 16100
rect 23772 16044 23828 16100
rect 24220 16098 24276 16100
rect 24220 16046 24222 16098
rect 24222 16046 24274 16098
rect 24274 16046 24276 16098
rect 24220 16044 24276 16046
rect 24780 16882 24836 16884
rect 24780 16830 24782 16882
rect 24782 16830 24834 16882
rect 24834 16830 24836 16882
rect 24780 16828 24836 16830
rect 24668 16044 24724 16100
rect 23436 15596 23492 15652
rect 23324 15372 23380 15428
rect 22876 15314 22932 15316
rect 22876 15262 22878 15314
rect 22878 15262 22930 15314
rect 22930 15262 22932 15314
rect 22876 15260 22932 15262
rect 22428 15202 22484 15204
rect 22428 15150 22430 15202
rect 22430 15150 22482 15202
rect 22482 15150 22484 15202
rect 22428 15148 22484 15150
rect 23100 13858 23156 13860
rect 23100 13806 23102 13858
rect 23102 13806 23154 13858
rect 23154 13806 23156 13858
rect 23100 13804 23156 13806
rect 24668 14812 24724 14868
rect 23996 13916 24052 13972
rect 23884 13804 23940 13860
rect 24556 13244 24612 13300
rect 22988 12908 23044 12964
rect 21980 11676 22036 11732
rect 21532 10722 21588 10724
rect 21532 10670 21534 10722
rect 21534 10670 21586 10722
rect 21586 10670 21588 10722
rect 21532 10668 21588 10670
rect 21644 9996 21700 10052
rect 21644 9266 21700 9268
rect 21644 9214 21646 9266
rect 21646 9214 21698 9266
rect 21698 9214 21700 9266
rect 21644 9212 21700 9214
rect 22876 11676 22932 11732
rect 22204 11394 22260 11396
rect 22204 11342 22206 11394
rect 22206 11342 22258 11394
rect 22258 11342 22260 11394
rect 22204 11340 22260 11342
rect 22316 10668 22372 10724
rect 22092 9884 22148 9940
rect 22316 9938 22372 9940
rect 22316 9886 22318 9938
rect 22318 9886 22370 9938
rect 22370 9886 22372 9938
rect 22316 9884 22372 9886
rect 23324 12402 23380 12404
rect 23324 12350 23326 12402
rect 23326 12350 23378 12402
rect 23378 12350 23380 12402
rect 23324 12348 23380 12350
rect 24332 11452 24388 11508
rect 22988 9884 23044 9940
rect 22652 9548 22708 9604
rect 22988 9602 23044 9604
rect 22988 9550 22990 9602
rect 22990 9550 23042 9602
rect 23042 9550 23044 9602
rect 22988 9548 23044 9550
rect 22652 9266 22708 9268
rect 22652 9214 22654 9266
rect 22654 9214 22706 9266
rect 22706 9214 22708 9266
rect 22652 9212 22708 9214
rect 22316 8988 22372 9044
rect 21420 8540 21476 8596
rect 21196 8428 21252 8484
rect 22652 8258 22708 8260
rect 22652 8206 22654 8258
rect 22654 8206 22706 8258
rect 22706 8206 22708 8258
rect 22652 8204 22708 8206
rect 21644 8034 21700 8036
rect 21644 7982 21646 8034
rect 21646 7982 21698 8034
rect 21698 7982 21700 8034
rect 21644 7980 21700 7982
rect 22428 8034 22484 8036
rect 22428 7982 22430 8034
rect 22430 7982 22482 8034
rect 22482 7982 22484 8034
rect 22428 7980 22484 7982
rect 22540 7868 22596 7924
rect 22204 7644 22260 7700
rect 21644 7532 21700 7588
rect 22092 7532 22148 7588
rect 20532 6298 20588 6300
rect 20532 6246 20534 6298
rect 20534 6246 20586 6298
rect 20586 6246 20588 6298
rect 20532 6244 20588 6246
rect 20636 6298 20692 6300
rect 20636 6246 20638 6298
rect 20638 6246 20690 6298
rect 20690 6246 20692 6298
rect 20636 6244 20692 6246
rect 20740 6298 20796 6300
rect 20740 6246 20742 6298
rect 20742 6246 20794 6298
rect 20794 6246 20796 6298
rect 20972 6300 21028 6356
rect 20740 6244 20796 6246
rect 20532 4730 20588 4732
rect 20532 4678 20534 4730
rect 20534 4678 20586 4730
rect 20586 4678 20588 4730
rect 20532 4676 20588 4678
rect 20636 4730 20692 4732
rect 20636 4678 20638 4730
rect 20638 4678 20690 4730
rect 20690 4678 20692 4730
rect 20636 4676 20692 4678
rect 20740 4730 20796 4732
rect 20740 4678 20742 4730
rect 20742 4678 20794 4730
rect 20794 4678 20796 4730
rect 20740 4676 20796 4678
rect 20300 4284 20356 4340
rect 20412 4172 20468 4228
rect 20188 3948 20244 4004
rect 21308 4172 21364 4228
rect 21420 4338 21476 4340
rect 21420 4286 21422 4338
rect 21422 4286 21474 4338
rect 21474 4286 21476 4338
rect 21420 4284 21476 4286
rect 20972 3500 21028 3556
rect 22316 7362 22372 7364
rect 22316 7310 22318 7362
rect 22318 7310 22370 7362
rect 22370 7310 22372 7362
rect 22316 7308 22372 7310
rect 22764 7532 22820 7588
rect 21980 5740 22036 5796
rect 22652 6690 22708 6692
rect 22652 6638 22654 6690
rect 22654 6638 22706 6690
rect 22706 6638 22708 6690
rect 22652 6636 22708 6638
rect 22876 5906 22932 5908
rect 22876 5854 22878 5906
rect 22878 5854 22930 5906
rect 22930 5854 22932 5906
rect 22876 5852 22932 5854
rect 22540 5740 22596 5796
rect 21980 5234 22036 5236
rect 21980 5182 21982 5234
rect 21982 5182 22034 5234
rect 22034 5182 22036 5234
rect 21980 5180 22036 5182
rect 23212 6188 23268 6244
rect 23548 9324 23604 9380
rect 23772 9324 23828 9380
rect 23996 9212 24052 9268
rect 24444 9602 24500 9604
rect 24444 9550 24446 9602
rect 24446 9550 24498 9602
rect 24498 9550 24500 9602
rect 24444 9548 24500 9550
rect 24332 9154 24388 9156
rect 24332 9102 24334 9154
rect 24334 9102 24386 9154
rect 24386 9102 24388 9154
rect 24332 9100 24388 9102
rect 23548 8428 23604 8484
rect 23436 8204 23492 8260
rect 23548 7980 23604 8036
rect 23660 7698 23716 7700
rect 23660 7646 23662 7698
rect 23662 7646 23714 7698
rect 23714 7646 23716 7698
rect 23660 7644 23716 7646
rect 24220 8370 24276 8372
rect 24220 8318 24222 8370
rect 24222 8318 24274 8370
rect 24274 8318 24276 8370
rect 24220 8316 24276 8318
rect 23884 7586 23940 7588
rect 23884 7534 23886 7586
rect 23886 7534 23938 7586
rect 23938 7534 23940 7586
rect 23884 7532 23940 7534
rect 23996 7308 24052 7364
rect 24220 7308 24276 7364
rect 23548 6636 23604 6692
rect 24108 6578 24164 6580
rect 24108 6526 24110 6578
rect 24110 6526 24162 6578
rect 24162 6526 24164 6578
rect 24108 6524 24164 6526
rect 23772 6300 23828 6356
rect 23660 6188 23716 6244
rect 23436 5794 23492 5796
rect 23436 5742 23438 5794
rect 23438 5742 23490 5794
rect 23490 5742 23492 5794
rect 23436 5740 23492 5742
rect 23436 4956 23492 5012
rect 23996 4732 24052 4788
rect 23100 4396 23156 4452
rect 21644 3948 21700 4004
rect 24108 4450 24164 4452
rect 24108 4398 24110 4450
rect 24110 4398 24162 4450
rect 24162 4398 24164 4450
rect 24108 4396 24164 4398
rect 24108 4060 24164 4116
rect 23996 3948 24052 4004
rect 22876 3836 22932 3892
rect 22652 3666 22708 3668
rect 22652 3614 22654 3666
rect 22654 3614 22706 3666
rect 22706 3614 22708 3666
rect 22652 3612 22708 3614
rect 20532 3162 20588 3164
rect 20532 3110 20534 3162
rect 20534 3110 20586 3162
rect 20586 3110 20588 3162
rect 20532 3108 20588 3110
rect 20636 3162 20692 3164
rect 20636 3110 20638 3162
rect 20638 3110 20690 3162
rect 20690 3110 20692 3162
rect 20636 3108 20692 3110
rect 20740 3162 20796 3164
rect 20740 3110 20742 3162
rect 20742 3110 20794 3162
rect 20794 3110 20796 3162
rect 21420 3164 21476 3220
rect 21868 3500 21924 3556
rect 20740 3108 20796 3110
rect 22092 3554 22148 3556
rect 22092 3502 22094 3554
rect 22094 3502 22146 3554
rect 22146 3502 22148 3554
rect 22092 3500 22148 3502
rect 23548 3442 23604 3444
rect 23548 3390 23550 3442
rect 23550 3390 23602 3442
rect 23602 3390 23604 3442
rect 23548 3388 23604 3390
rect 24332 6690 24388 6692
rect 24332 6638 24334 6690
rect 24334 6638 24386 6690
rect 24386 6638 24388 6690
rect 24332 6636 24388 6638
rect 24444 6300 24500 6356
rect 24444 5906 24500 5908
rect 24444 5854 24446 5906
rect 24446 5854 24498 5906
rect 24498 5854 24500 5906
rect 24444 5852 24500 5854
rect 25004 13746 25060 13748
rect 25004 13694 25006 13746
rect 25006 13694 25058 13746
rect 25058 13694 25060 13746
rect 25004 13692 25060 13694
rect 25004 12684 25060 12740
rect 24668 12124 24724 12180
rect 24892 11788 24948 11844
rect 25004 11506 25060 11508
rect 25004 11454 25006 11506
rect 25006 11454 25058 11506
rect 25058 11454 25060 11506
rect 25004 11452 25060 11454
rect 24892 11394 24948 11396
rect 24892 11342 24894 11394
rect 24894 11342 24946 11394
rect 24946 11342 24948 11394
rect 24892 11340 24948 11342
rect 26124 21586 26180 21588
rect 26124 21534 26126 21586
rect 26126 21534 26178 21586
rect 26178 21534 26180 21586
rect 26124 21532 26180 21534
rect 26684 22652 26740 22708
rect 26572 21532 26628 21588
rect 26796 22204 26852 22260
rect 28364 27298 28420 27300
rect 28364 27246 28366 27298
rect 28366 27246 28418 27298
rect 28418 27246 28420 27298
rect 28364 27244 28420 27246
rect 28252 26908 28308 26964
rect 27916 26796 27972 26852
rect 28028 25618 28084 25620
rect 28028 25566 28030 25618
rect 28030 25566 28082 25618
rect 28082 25566 28084 25618
rect 28028 25564 28084 25566
rect 27916 25506 27972 25508
rect 27916 25454 27918 25506
rect 27918 25454 27970 25506
rect 27970 25454 27972 25506
rect 27916 25452 27972 25454
rect 28700 28530 28756 28532
rect 28700 28478 28702 28530
rect 28702 28478 28754 28530
rect 28754 28478 28756 28530
rect 28700 28476 28756 28478
rect 28588 27970 28644 27972
rect 28588 27918 28590 27970
rect 28590 27918 28642 27970
rect 28642 27918 28644 27970
rect 28588 27916 28644 27918
rect 28700 27692 28756 27748
rect 27244 24050 27300 24052
rect 27244 23998 27246 24050
rect 27246 23998 27298 24050
rect 27298 23998 27300 24050
rect 27244 23996 27300 23998
rect 27356 23436 27412 23492
rect 28252 23996 28308 24052
rect 27916 23826 27972 23828
rect 27916 23774 27918 23826
rect 27918 23774 27970 23826
rect 27970 23774 27972 23826
rect 27916 23772 27972 23774
rect 28252 23772 28308 23828
rect 27132 22092 27188 22148
rect 26012 20860 26068 20916
rect 26460 20690 26516 20692
rect 26460 20638 26462 20690
rect 26462 20638 26514 20690
rect 26514 20638 26516 20690
rect 26460 20636 26516 20638
rect 25788 20188 25844 20244
rect 26124 20412 26180 20468
rect 25900 19516 25956 19572
rect 25676 18562 25732 18564
rect 25676 18510 25678 18562
rect 25678 18510 25730 18562
rect 25730 18510 25732 18562
rect 25676 18508 25732 18510
rect 25900 18396 25956 18452
rect 26012 18844 26068 18900
rect 25228 17612 25284 17668
rect 25900 17388 25956 17444
rect 25788 16828 25844 16884
rect 26572 20578 26628 20580
rect 26572 20526 26574 20578
rect 26574 20526 26626 20578
rect 26626 20526 26628 20578
rect 26572 20524 26628 20526
rect 26460 20300 26516 20356
rect 26348 19516 26404 19572
rect 26236 19458 26292 19460
rect 26236 19406 26238 19458
rect 26238 19406 26290 19458
rect 26290 19406 26292 19458
rect 26236 19404 26292 19406
rect 26348 19234 26404 19236
rect 26348 19182 26350 19234
rect 26350 19182 26402 19234
rect 26402 19182 26404 19234
rect 26348 19180 26404 19182
rect 26236 19122 26292 19124
rect 26236 19070 26238 19122
rect 26238 19070 26290 19122
rect 26290 19070 26292 19122
rect 26236 19068 26292 19070
rect 27692 22092 27748 22148
rect 27580 21980 27636 22036
rect 27580 21586 27636 21588
rect 27580 21534 27582 21586
rect 27582 21534 27634 21586
rect 27634 21534 27636 21586
rect 27580 21532 27636 21534
rect 27916 22652 27972 22708
rect 27468 20914 27524 20916
rect 27468 20862 27470 20914
rect 27470 20862 27522 20914
rect 27522 20862 27524 20914
rect 27468 20860 27524 20862
rect 28140 22146 28196 22148
rect 28140 22094 28142 22146
rect 28142 22094 28194 22146
rect 28194 22094 28196 22146
rect 28140 22092 28196 22094
rect 28588 21980 28644 22036
rect 28812 26962 28868 26964
rect 28812 26910 28814 26962
rect 28814 26910 28866 26962
rect 28866 26910 28868 26962
rect 28812 26908 28868 26910
rect 29036 27244 29092 27300
rect 28924 26796 28980 26852
rect 29148 22652 29204 22708
rect 27804 20578 27860 20580
rect 27804 20526 27806 20578
rect 27806 20526 27858 20578
rect 27858 20526 27860 20578
rect 27804 20524 27860 20526
rect 27468 20412 27524 20468
rect 27468 20242 27524 20244
rect 27468 20190 27470 20242
rect 27470 20190 27522 20242
rect 27522 20190 27524 20242
rect 27468 20188 27524 20190
rect 27804 20188 27860 20244
rect 26908 19906 26964 19908
rect 26908 19854 26910 19906
rect 26910 19854 26962 19906
rect 26962 19854 26964 19906
rect 26908 19852 26964 19854
rect 27692 19852 27748 19908
rect 26908 19122 26964 19124
rect 26908 19070 26910 19122
rect 26910 19070 26962 19122
rect 26962 19070 26964 19122
rect 26908 19068 26964 19070
rect 27468 19122 27524 19124
rect 27468 19070 27470 19122
rect 27470 19070 27522 19122
rect 27522 19070 27524 19122
rect 27468 19068 27524 19070
rect 26684 18450 26740 18452
rect 26684 18398 26686 18450
rect 26686 18398 26738 18450
rect 26738 18398 26740 18450
rect 26684 18396 26740 18398
rect 27132 18450 27188 18452
rect 27132 18398 27134 18450
rect 27134 18398 27186 18450
rect 27186 18398 27188 18450
rect 27132 18396 27188 18398
rect 26348 17554 26404 17556
rect 26348 17502 26350 17554
rect 26350 17502 26402 17554
rect 26402 17502 26404 17554
rect 26348 17500 26404 17502
rect 26124 16828 26180 16884
rect 26460 17442 26516 17444
rect 26460 17390 26462 17442
rect 26462 17390 26514 17442
rect 26514 17390 26516 17442
rect 26460 17388 26516 17390
rect 26572 17276 26628 17332
rect 26124 15932 26180 15988
rect 26460 16044 26516 16100
rect 27580 18396 27636 18452
rect 28364 20300 28420 20356
rect 27916 19740 27972 19796
rect 28252 19794 28308 19796
rect 28252 19742 28254 19794
rect 28254 19742 28306 19794
rect 28306 19742 28308 19794
rect 28252 19740 28308 19742
rect 28252 18844 28308 18900
rect 27468 17388 27524 17444
rect 27804 18396 27860 18452
rect 28028 18450 28084 18452
rect 28028 18398 28030 18450
rect 28030 18398 28082 18450
rect 28082 18398 28084 18450
rect 28028 18396 28084 18398
rect 28364 18284 28420 18340
rect 28812 20300 28868 20356
rect 29036 20636 29092 20692
rect 28700 19292 28756 19348
rect 29148 20188 29204 20244
rect 29036 19906 29092 19908
rect 29036 19854 29038 19906
rect 29038 19854 29090 19906
rect 29090 19854 29092 19906
rect 29036 19852 29092 19854
rect 28700 18844 28756 18900
rect 28028 16940 28084 16996
rect 28588 18338 28644 18340
rect 28588 18286 28590 18338
rect 28590 18286 28642 18338
rect 28642 18286 28644 18338
rect 28588 18284 28644 18286
rect 28028 16770 28084 16772
rect 28028 16718 28030 16770
rect 28030 16718 28082 16770
rect 28082 16718 28084 16770
rect 28028 16716 28084 16718
rect 27244 16098 27300 16100
rect 27244 16046 27246 16098
rect 27246 16046 27298 16098
rect 27298 16046 27300 16098
rect 27244 16044 27300 16046
rect 27132 15986 27188 15988
rect 27132 15934 27134 15986
rect 27134 15934 27186 15986
rect 27186 15934 27188 15986
rect 27132 15932 27188 15934
rect 25452 14812 25508 14868
rect 25452 13804 25508 13860
rect 25564 13746 25620 13748
rect 25564 13694 25566 13746
rect 25566 13694 25618 13746
rect 25618 13694 25620 13746
rect 25564 13692 25620 13694
rect 25452 13356 25508 13412
rect 25228 12124 25284 12180
rect 25116 10108 25172 10164
rect 25004 9772 25060 9828
rect 24668 8034 24724 8036
rect 24668 7982 24670 8034
rect 24670 7982 24722 8034
rect 24722 7982 24724 8034
rect 24668 7980 24724 7982
rect 24780 6524 24836 6580
rect 24668 4956 24724 5012
rect 24780 4732 24836 4788
rect 24892 4956 24948 5012
rect 24668 4508 24724 4564
rect 24556 4284 24612 4340
rect 24444 3612 24500 3668
rect 24780 3836 24836 3892
rect 24556 3554 24612 3556
rect 24556 3502 24558 3554
rect 24558 3502 24610 3554
rect 24610 3502 24612 3554
rect 24556 3500 24612 3502
rect 24108 2828 24164 2884
rect 26796 14364 26852 14420
rect 26012 13858 26068 13860
rect 26012 13806 26014 13858
rect 26014 13806 26066 13858
rect 26066 13806 26068 13858
rect 26012 13804 26068 13806
rect 26684 13858 26740 13860
rect 26684 13806 26686 13858
rect 26686 13806 26738 13858
rect 26738 13806 26740 13858
rect 26684 13804 26740 13806
rect 26124 13634 26180 13636
rect 26124 13582 26126 13634
rect 26126 13582 26178 13634
rect 26178 13582 26180 13634
rect 26124 13580 26180 13582
rect 27692 14418 27748 14420
rect 27692 14366 27694 14418
rect 27694 14366 27746 14418
rect 27746 14366 27748 14418
rect 27692 14364 27748 14366
rect 27468 14252 27524 14308
rect 27468 13746 27524 13748
rect 27468 13694 27470 13746
rect 27470 13694 27522 13746
rect 27522 13694 27524 13746
rect 27468 13692 27524 13694
rect 25452 9826 25508 9828
rect 25452 9774 25454 9826
rect 25454 9774 25506 9826
rect 25506 9774 25508 9826
rect 25452 9772 25508 9774
rect 27356 12738 27412 12740
rect 27356 12686 27358 12738
rect 27358 12686 27410 12738
rect 27410 12686 27412 12738
rect 27356 12684 27412 12686
rect 25676 11452 25732 11508
rect 26796 12124 26852 12180
rect 26012 11788 26068 11844
rect 26684 11788 26740 11844
rect 27580 11564 27636 11620
rect 25788 11394 25844 11396
rect 25788 11342 25790 11394
rect 25790 11342 25842 11394
rect 25842 11342 25844 11394
rect 25788 11340 25844 11342
rect 25788 11116 25844 11172
rect 26908 11394 26964 11396
rect 26908 11342 26910 11394
rect 26910 11342 26962 11394
rect 26962 11342 26964 11394
rect 26908 11340 26964 11342
rect 28812 17666 28868 17668
rect 28812 17614 28814 17666
rect 28814 17614 28866 17666
rect 28866 17614 28868 17666
rect 28812 17612 28868 17614
rect 29148 17612 29204 17668
rect 29148 17106 29204 17108
rect 29148 17054 29150 17106
rect 29150 17054 29202 17106
rect 29202 17054 29204 17106
rect 29148 17052 29204 17054
rect 30604 30716 30660 30772
rect 30192 30602 30248 30604
rect 30192 30550 30194 30602
rect 30194 30550 30246 30602
rect 30246 30550 30248 30602
rect 30192 30548 30248 30550
rect 30296 30602 30352 30604
rect 30296 30550 30298 30602
rect 30298 30550 30350 30602
rect 30350 30550 30352 30602
rect 30296 30548 30352 30550
rect 30400 30602 30456 30604
rect 30400 30550 30402 30602
rect 30402 30550 30454 30602
rect 30454 30550 30456 30602
rect 30400 30548 30456 30550
rect 30268 30268 30324 30324
rect 30044 30210 30100 30212
rect 30044 30158 30046 30210
rect 30046 30158 30098 30210
rect 30098 30158 30100 30210
rect 30044 30156 30100 30158
rect 31612 30940 31668 30996
rect 30604 30156 30660 30212
rect 30268 29932 30324 29988
rect 33404 32508 33460 32564
rect 32172 31948 32228 32004
rect 33404 31948 33460 32004
rect 33180 31500 33236 31556
rect 33964 34130 34020 34132
rect 33964 34078 33966 34130
rect 33966 34078 34018 34130
rect 34018 34078 34020 34130
rect 33964 34076 34020 34078
rect 35420 34860 35476 34916
rect 35644 34914 35700 34916
rect 35644 34862 35646 34914
rect 35646 34862 35698 34914
rect 35698 34862 35700 34914
rect 35644 34860 35700 34862
rect 36988 36204 37044 36260
rect 36988 35196 37044 35252
rect 36540 34914 36596 34916
rect 36540 34862 36542 34914
rect 36542 34862 36594 34914
rect 36594 34862 36596 34914
rect 36540 34860 36596 34862
rect 36652 34802 36708 34804
rect 36652 34750 36654 34802
rect 36654 34750 36706 34802
rect 36706 34750 36708 34802
rect 36652 34748 36708 34750
rect 36204 34636 36260 34692
rect 35756 34242 35812 34244
rect 35756 34190 35758 34242
rect 35758 34190 35810 34242
rect 35810 34190 35812 34242
rect 35756 34188 35812 34190
rect 36764 33852 36820 33908
rect 38668 36482 38724 36484
rect 38668 36430 38670 36482
rect 38670 36430 38722 36482
rect 38722 36430 38724 36482
rect 38668 36428 38724 36430
rect 37660 35532 37716 35588
rect 38108 35586 38164 35588
rect 38108 35534 38110 35586
rect 38110 35534 38162 35586
rect 38162 35534 38164 35586
rect 38108 35532 38164 35534
rect 37436 34860 37492 34916
rect 37548 34802 37604 34804
rect 37548 34750 37550 34802
rect 37550 34750 37602 34802
rect 37602 34750 37604 34802
rect 37548 34748 37604 34750
rect 37660 34690 37716 34692
rect 37660 34638 37662 34690
rect 37662 34638 37714 34690
rect 37714 34638 37716 34690
rect 37660 34636 37716 34638
rect 39852 36090 39908 36092
rect 39852 36038 39854 36090
rect 39854 36038 39906 36090
rect 39906 36038 39908 36090
rect 39852 36036 39908 36038
rect 39956 36090 40012 36092
rect 39956 36038 39958 36090
rect 39958 36038 40010 36090
rect 40010 36038 40012 36090
rect 39956 36036 40012 36038
rect 40060 36090 40116 36092
rect 40060 36038 40062 36090
rect 40062 36038 40114 36090
rect 40114 36038 40116 36090
rect 40060 36036 40116 36038
rect 40124 35868 40180 35924
rect 42588 36204 42644 36260
rect 43036 36258 43092 36260
rect 43036 36206 43038 36258
rect 43038 36206 43090 36258
rect 43090 36206 43092 36258
rect 43036 36204 43092 36206
rect 42700 36092 42756 36148
rect 40572 35922 40628 35924
rect 40572 35870 40574 35922
rect 40574 35870 40626 35922
rect 40626 35870 40628 35922
rect 40572 35868 40628 35870
rect 49512 36874 49568 36876
rect 49512 36822 49514 36874
rect 49514 36822 49566 36874
rect 49566 36822 49568 36874
rect 49512 36820 49568 36822
rect 49616 36874 49672 36876
rect 49616 36822 49618 36874
rect 49618 36822 49670 36874
rect 49670 36822 49672 36874
rect 49616 36820 49672 36822
rect 49720 36874 49776 36876
rect 49720 36822 49722 36874
rect 49722 36822 49774 36874
rect 49774 36822 49776 36874
rect 49720 36820 49776 36822
rect 48524 36540 48580 36596
rect 48972 36594 49028 36596
rect 48972 36542 48974 36594
rect 48974 36542 49026 36594
rect 49026 36542 49028 36594
rect 48972 36540 49028 36542
rect 52220 36764 52276 36820
rect 43820 36428 43876 36484
rect 40236 35196 40292 35252
rect 39852 34522 39908 34524
rect 39852 34470 39854 34522
rect 39854 34470 39906 34522
rect 39906 34470 39908 34522
rect 39852 34468 39908 34470
rect 39956 34522 40012 34524
rect 39956 34470 39958 34522
rect 39958 34470 40010 34522
rect 40010 34470 40012 34522
rect 39956 34468 40012 34470
rect 40060 34522 40116 34524
rect 40060 34470 40062 34522
rect 40062 34470 40114 34522
rect 40114 34470 40116 34522
rect 40060 34468 40116 34470
rect 39676 34300 39732 34356
rect 40460 34914 40516 34916
rect 40460 34862 40462 34914
rect 40462 34862 40514 34914
rect 40514 34862 40516 34914
rect 40460 34860 40516 34862
rect 41356 34914 41412 34916
rect 41356 34862 41358 34914
rect 41358 34862 41410 34914
rect 41410 34862 41412 34914
rect 41356 34860 41412 34862
rect 44156 35644 44212 35700
rect 44380 36204 44436 36260
rect 42028 34860 42084 34916
rect 40460 34354 40516 34356
rect 40460 34302 40462 34354
rect 40462 34302 40514 34354
rect 40514 34302 40516 34354
rect 40460 34300 40516 34302
rect 40684 34354 40740 34356
rect 40684 34302 40686 34354
rect 40686 34302 40738 34354
rect 40738 34302 40740 34354
rect 40684 34300 40740 34302
rect 37212 33906 37268 33908
rect 37212 33854 37214 33906
rect 37214 33854 37266 33906
rect 37266 33854 37268 33906
rect 37212 33852 37268 33854
rect 38668 33852 38724 33908
rect 37324 33292 37380 33348
rect 36876 33122 36932 33124
rect 36876 33070 36878 33122
rect 36878 33070 36930 33122
rect 36930 33070 36932 33122
rect 36876 33068 36932 33070
rect 33852 32562 33908 32564
rect 33852 32510 33854 32562
rect 33854 32510 33906 32562
rect 33906 32510 33908 32562
rect 33852 32508 33908 32510
rect 37996 33068 38052 33124
rect 38556 33068 38612 33124
rect 41468 34188 41524 34244
rect 41692 34188 41748 34244
rect 42812 34300 42868 34356
rect 42252 33906 42308 33908
rect 42252 33854 42254 33906
rect 42254 33854 42306 33906
rect 42306 33854 42308 33906
rect 42252 33852 42308 33854
rect 43484 34636 43540 34692
rect 43596 34300 43652 34356
rect 43932 34242 43988 34244
rect 43932 34190 43934 34242
rect 43934 34190 43986 34242
rect 43986 34190 43988 34242
rect 43932 34188 43988 34190
rect 42812 33740 42868 33796
rect 39340 33346 39396 33348
rect 39340 33294 39342 33346
rect 39342 33294 39394 33346
rect 39394 33294 39396 33346
rect 39340 33292 39396 33294
rect 39228 33068 39284 33124
rect 39852 32954 39908 32956
rect 39852 32902 39854 32954
rect 39854 32902 39906 32954
rect 39906 32902 39908 32954
rect 39852 32900 39908 32902
rect 39956 32954 40012 32956
rect 39956 32902 39958 32954
rect 39958 32902 40010 32954
rect 40010 32902 40012 32954
rect 39956 32900 40012 32902
rect 40060 32954 40116 32956
rect 40060 32902 40062 32954
rect 40062 32902 40114 32954
rect 40114 32902 40116 32954
rect 40060 32900 40116 32902
rect 43148 33346 43204 33348
rect 43148 33294 43150 33346
rect 43150 33294 43202 33346
rect 43202 33294 43204 33346
rect 43148 33292 43204 33294
rect 44044 33852 44100 33908
rect 43484 33292 43540 33348
rect 44268 33346 44324 33348
rect 44268 33294 44270 33346
rect 44270 33294 44322 33346
rect 44322 33294 44324 33346
rect 44268 33292 44324 33294
rect 43932 33180 43988 33236
rect 37100 32450 37156 32452
rect 37100 32398 37102 32450
rect 37102 32398 37154 32450
rect 37154 32398 37156 32450
rect 37100 32396 37156 32398
rect 37324 31948 37380 32004
rect 37548 32396 37604 32452
rect 33516 31500 33572 31556
rect 32060 30770 32116 30772
rect 32060 30718 32062 30770
rect 32062 30718 32114 30770
rect 32114 30718 32116 30770
rect 32060 30716 32116 30718
rect 32284 30268 32340 30324
rect 33740 30268 33796 30324
rect 31612 30098 31668 30100
rect 31612 30046 31614 30098
rect 31614 30046 31666 30098
rect 31666 30046 31668 30098
rect 31612 30044 31668 30046
rect 32172 30098 32228 30100
rect 32172 30046 32174 30098
rect 32174 30046 32226 30098
rect 32226 30046 32228 30098
rect 32172 30044 32228 30046
rect 29820 29708 29876 29764
rect 30192 29034 30248 29036
rect 30192 28982 30194 29034
rect 30194 28982 30246 29034
rect 30246 28982 30248 29034
rect 30192 28980 30248 28982
rect 30296 29034 30352 29036
rect 30296 28982 30298 29034
rect 30298 28982 30350 29034
rect 30350 28982 30352 29034
rect 30296 28980 30352 28982
rect 30400 29034 30456 29036
rect 30400 28982 30402 29034
rect 30402 28982 30454 29034
rect 30454 28982 30456 29034
rect 30400 28980 30456 28982
rect 34524 30604 34580 30660
rect 34524 30268 34580 30324
rect 33068 29484 33124 29540
rect 32396 29426 32452 29428
rect 32396 29374 32398 29426
rect 32398 29374 32450 29426
rect 32450 29374 32452 29426
rect 32396 29372 32452 29374
rect 32732 29314 32788 29316
rect 32732 29262 32734 29314
rect 32734 29262 32786 29314
rect 32786 29262 32788 29314
rect 32732 29260 32788 29262
rect 29708 28642 29764 28644
rect 29708 28590 29710 28642
rect 29710 28590 29762 28642
rect 29762 28590 29764 28642
rect 29708 28588 29764 28590
rect 29932 28476 29988 28532
rect 31052 28588 31108 28644
rect 30716 27970 30772 27972
rect 30716 27918 30718 27970
rect 30718 27918 30770 27970
rect 30770 27918 30772 27970
rect 30716 27916 30772 27918
rect 30044 27858 30100 27860
rect 30044 27806 30046 27858
rect 30046 27806 30098 27858
rect 30098 27806 30100 27858
rect 30044 27804 30100 27806
rect 30192 27466 30248 27468
rect 30192 27414 30194 27466
rect 30194 27414 30246 27466
rect 30246 27414 30248 27466
rect 30192 27412 30248 27414
rect 30296 27466 30352 27468
rect 30296 27414 30298 27466
rect 30298 27414 30350 27466
rect 30350 27414 30352 27466
rect 30296 27412 30352 27414
rect 30400 27466 30456 27468
rect 30400 27414 30402 27466
rect 30402 27414 30454 27466
rect 30454 27414 30456 27466
rect 30400 27412 30456 27414
rect 30828 27858 30884 27860
rect 30828 27806 30830 27858
rect 30830 27806 30882 27858
rect 30882 27806 30884 27858
rect 30828 27804 30884 27806
rect 30716 27634 30772 27636
rect 30716 27582 30718 27634
rect 30718 27582 30770 27634
rect 30770 27582 30772 27634
rect 30716 27580 30772 27582
rect 30940 26908 30996 26964
rect 29820 26290 29876 26292
rect 29820 26238 29822 26290
rect 29822 26238 29874 26290
rect 29874 26238 29876 26290
rect 29820 26236 29876 26238
rect 30940 26290 30996 26292
rect 30940 26238 30942 26290
rect 30942 26238 30994 26290
rect 30994 26238 30996 26290
rect 30940 26236 30996 26238
rect 29708 25564 29764 25620
rect 29820 26012 29876 26068
rect 29596 23324 29652 23380
rect 29708 23772 29764 23828
rect 30492 26012 30548 26068
rect 30192 25898 30248 25900
rect 30192 25846 30194 25898
rect 30194 25846 30246 25898
rect 30246 25846 30248 25898
rect 30192 25844 30248 25846
rect 30296 25898 30352 25900
rect 30296 25846 30298 25898
rect 30298 25846 30350 25898
rect 30350 25846 30352 25898
rect 30296 25844 30352 25846
rect 30400 25898 30456 25900
rect 30400 25846 30402 25898
rect 30402 25846 30454 25898
rect 30454 25846 30456 25898
rect 30400 25844 30456 25846
rect 30940 25340 30996 25396
rect 30604 24780 30660 24836
rect 30492 24722 30548 24724
rect 30492 24670 30494 24722
rect 30494 24670 30546 24722
rect 30546 24670 30548 24722
rect 30492 24668 30548 24670
rect 30192 24330 30248 24332
rect 30192 24278 30194 24330
rect 30194 24278 30246 24330
rect 30246 24278 30248 24330
rect 30192 24276 30248 24278
rect 30296 24330 30352 24332
rect 30296 24278 30298 24330
rect 30298 24278 30350 24330
rect 30350 24278 30352 24330
rect 30296 24276 30352 24278
rect 30400 24330 30456 24332
rect 30400 24278 30402 24330
rect 30402 24278 30454 24330
rect 30454 24278 30456 24330
rect 30400 24276 30456 24278
rect 30716 24668 30772 24724
rect 30044 23772 30100 23828
rect 30268 23826 30324 23828
rect 30268 23774 30270 23826
rect 30270 23774 30322 23826
rect 30322 23774 30324 23826
rect 30268 23772 30324 23774
rect 30380 23714 30436 23716
rect 30380 23662 30382 23714
rect 30382 23662 30434 23714
rect 30434 23662 30436 23714
rect 30380 23660 30436 23662
rect 31612 28642 31668 28644
rect 31612 28590 31614 28642
rect 31614 28590 31666 28642
rect 31666 28590 31668 28642
rect 31612 28588 31668 28590
rect 32508 28642 32564 28644
rect 32508 28590 32510 28642
rect 32510 28590 32562 28642
rect 32562 28590 32564 28642
rect 32508 28588 32564 28590
rect 32396 28476 32452 28532
rect 31164 27804 31220 27860
rect 31612 27580 31668 27636
rect 31724 27804 31780 27860
rect 31388 27020 31444 27076
rect 31500 26962 31556 26964
rect 31500 26910 31502 26962
rect 31502 26910 31554 26962
rect 31554 26910 31556 26962
rect 31500 26908 31556 26910
rect 31724 26962 31780 26964
rect 31724 26910 31726 26962
rect 31726 26910 31778 26962
rect 31778 26910 31780 26962
rect 31724 26908 31780 26910
rect 32060 27074 32116 27076
rect 32060 27022 32062 27074
rect 32062 27022 32114 27074
rect 32114 27022 32116 27074
rect 32060 27020 32116 27022
rect 32396 26962 32452 26964
rect 32396 26910 32398 26962
rect 32398 26910 32450 26962
rect 32450 26910 32452 26962
rect 32396 26908 32452 26910
rect 32284 26290 32340 26292
rect 32284 26238 32286 26290
rect 32286 26238 32338 26290
rect 32338 26238 32340 26290
rect 32284 26236 32340 26238
rect 32396 26178 32452 26180
rect 32396 26126 32398 26178
rect 32398 26126 32450 26178
rect 32450 26126 32452 26178
rect 32396 26124 32452 26126
rect 32508 26012 32564 26068
rect 33068 25452 33124 25508
rect 33180 25394 33236 25396
rect 33180 25342 33182 25394
rect 33182 25342 33234 25394
rect 33234 25342 33236 25394
rect 33180 25340 33236 25342
rect 32732 24834 32788 24836
rect 32732 24782 32734 24834
rect 32734 24782 32786 24834
rect 32786 24782 32788 24834
rect 32732 24780 32788 24782
rect 32508 24722 32564 24724
rect 32508 24670 32510 24722
rect 32510 24670 32562 24722
rect 32562 24670 32564 24722
rect 32508 24668 32564 24670
rect 31052 24444 31108 24500
rect 32844 24556 32900 24612
rect 30716 23660 30772 23716
rect 32620 23714 32676 23716
rect 32620 23662 32622 23714
rect 32622 23662 32674 23714
rect 32674 23662 32676 23714
rect 32620 23660 32676 23662
rect 30192 22762 30248 22764
rect 30192 22710 30194 22762
rect 30194 22710 30246 22762
rect 30246 22710 30248 22762
rect 30192 22708 30248 22710
rect 30296 22762 30352 22764
rect 30296 22710 30298 22762
rect 30298 22710 30350 22762
rect 30350 22710 30352 22762
rect 30296 22708 30352 22710
rect 30400 22762 30456 22764
rect 30400 22710 30402 22762
rect 30402 22710 30454 22762
rect 30454 22710 30456 22762
rect 30400 22708 30456 22710
rect 30716 22652 30772 22708
rect 30604 22092 30660 22148
rect 30192 21194 30248 21196
rect 30192 21142 30194 21194
rect 30194 21142 30246 21194
rect 30246 21142 30248 21194
rect 30192 21140 30248 21142
rect 30296 21194 30352 21196
rect 30296 21142 30298 21194
rect 30298 21142 30350 21194
rect 30350 21142 30352 21194
rect 30296 21140 30352 21142
rect 30400 21194 30456 21196
rect 30400 21142 30402 21194
rect 30402 21142 30454 21194
rect 30454 21142 30456 21194
rect 30400 21140 30456 21142
rect 30716 21644 30772 21700
rect 30604 20972 30660 21028
rect 29708 20636 29764 20692
rect 29596 20300 29652 20356
rect 29596 19852 29652 19908
rect 30828 20188 30884 20244
rect 30604 19740 30660 19796
rect 30192 19626 30248 19628
rect 30192 19574 30194 19626
rect 30194 19574 30246 19626
rect 30246 19574 30248 19626
rect 30192 19572 30248 19574
rect 30296 19626 30352 19628
rect 30296 19574 30298 19626
rect 30298 19574 30350 19626
rect 30350 19574 30352 19626
rect 30296 19572 30352 19574
rect 30400 19626 30456 19628
rect 30400 19574 30402 19626
rect 30402 19574 30454 19626
rect 30454 19574 30456 19626
rect 30400 19572 30456 19574
rect 30940 19180 30996 19236
rect 30492 19068 30548 19124
rect 29596 18844 29652 18900
rect 29596 17442 29652 17444
rect 29596 17390 29598 17442
rect 29598 17390 29650 17442
rect 29650 17390 29652 17442
rect 29596 17388 29652 17390
rect 29932 18562 29988 18564
rect 29932 18510 29934 18562
rect 29934 18510 29986 18562
rect 29986 18510 29988 18562
rect 29932 18508 29988 18510
rect 29260 16716 29316 16772
rect 29596 16770 29652 16772
rect 29596 16718 29598 16770
rect 29598 16718 29650 16770
rect 29650 16718 29652 16770
rect 29596 16716 29652 16718
rect 28588 16604 28644 16660
rect 28924 15820 28980 15876
rect 28028 14252 28084 14308
rect 28812 14418 28868 14420
rect 28812 14366 28814 14418
rect 28814 14366 28866 14418
rect 28866 14366 28868 14418
rect 28812 14364 28868 14366
rect 28700 14306 28756 14308
rect 28700 14254 28702 14306
rect 28702 14254 28754 14306
rect 28754 14254 28756 14306
rect 28700 14252 28756 14254
rect 28140 13746 28196 13748
rect 28140 13694 28142 13746
rect 28142 13694 28194 13746
rect 28194 13694 28196 13746
rect 28140 13692 28196 13694
rect 28812 13692 28868 13748
rect 28028 13634 28084 13636
rect 28028 13582 28030 13634
rect 28030 13582 28082 13634
rect 28082 13582 28084 13634
rect 28028 13580 28084 13582
rect 29708 16492 29764 16548
rect 29708 15874 29764 15876
rect 29708 15822 29710 15874
rect 29710 15822 29762 15874
rect 29762 15822 29764 15874
rect 29708 15820 29764 15822
rect 31052 18508 31108 18564
rect 31164 19852 31220 19908
rect 30156 18450 30212 18452
rect 30156 18398 30158 18450
rect 30158 18398 30210 18450
rect 30210 18398 30212 18450
rect 30156 18396 30212 18398
rect 30604 18284 30660 18340
rect 30192 18058 30248 18060
rect 30192 18006 30194 18058
rect 30194 18006 30246 18058
rect 30246 18006 30248 18058
rect 30192 18004 30248 18006
rect 30296 18058 30352 18060
rect 30296 18006 30298 18058
rect 30298 18006 30350 18058
rect 30350 18006 30352 18058
rect 30296 18004 30352 18006
rect 30400 18058 30456 18060
rect 30400 18006 30402 18058
rect 30402 18006 30454 18058
rect 30454 18006 30456 18058
rect 30400 18004 30456 18006
rect 32732 20524 32788 20580
rect 31724 19068 31780 19124
rect 31500 19010 31556 19012
rect 31500 18958 31502 19010
rect 31502 18958 31554 19010
rect 31554 18958 31556 19010
rect 31500 18956 31556 18958
rect 31388 18844 31444 18900
rect 31388 18674 31444 18676
rect 31388 18622 31390 18674
rect 31390 18622 31442 18674
rect 31442 18622 31444 18674
rect 31388 18620 31444 18622
rect 31276 18284 31332 18340
rect 30156 17388 30212 17444
rect 30268 17106 30324 17108
rect 30268 17054 30270 17106
rect 30270 17054 30322 17106
rect 30322 17054 30324 17106
rect 30268 17052 30324 17054
rect 30156 16716 30212 16772
rect 30828 16828 30884 16884
rect 30192 16490 30248 16492
rect 30192 16438 30194 16490
rect 30194 16438 30246 16490
rect 30246 16438 30248 16490
rect 30192 16436 30248 16438
rect 30296 16490 30352 16492
rect 30296 16438 30298 16490
rect 30298 16438 30350 16490
rect 30350 16438 30352 16490
rect 30296 16436 30352 16438
rect 30400 16490 30456 16492
rect 30400 16438 30402 16490
rect 30402 16438 30454 16490
rect 30454 16438 30456 16490
rect 30400 16436 30456 16438
rect 30268 16210 30324 16212
rect 30268 16158 30270 16210
rect 30270 16158 30322 16210
rect 30322 16158 30324 16210
rect 30268 16156 30324 16158
rect 30828 16156 30884 16212
rect 31164 15874 31220 15876
rect 31164 15822 31166 15874
rect 31166 15822 31218 15874
rect 31218 15822 31220 15874
rect 31164 15820 31220 15822
rect 29932 15372 29988 15428
rect 29596 15148 29652 15204
rect 30044 15202 30100 15204
rect 30044 15150 30046 15202
rect 30046 15150 30098 15202
rect 30098 15150 30100 15202
rect 30044 15148 30100 15150
rect 30716 15148 30772 15204
rect 30192 14922 30248 14924
rect 30192 14870 30194 14922
rect 30194 14870 30246 14922
rect 30246 14870 30248 14922
rect 30192 14868 30248 14870
rect 30296 14922 30352 14924
rect 30296 14870 30298 14922
rect 30298 14870 30350 14922
rect 30350 14870 30352 14922
rect 30296 14868 30352 14870
rect 30400 14922 30456 14924
rect 30400 14870 30402 14922
rect 30402 14870 30454 14922
rect 30454 14870 30456 14922
rect 30400 14868 30456 14870
rect 30156 13858 30212 13860
rect 30156 13806 30158 13858
rect 30158 13806 30210 13858
rect 30210 13806 30212 13858
rect 30156 13804 30212 13806
rect 29484 13746 29540 13748
rect 29484 13694 29486 13746
rect 29486 13694 29538 13746
rect 29538 13694 29540 13746
rect 29484 13692 29540 13694
rect 28924 13244 28980 13300
rect 30192 13354 30248 13356
rect 30192 13302 30194 13354
rect 30194 13302 30246 13354
rect 30246 13302 30248 13354
rect 30192 13300 30248 13302
rect 30296 13354 30352 13356
rect 30296 13302 30298 13354
rect 30298 13302 30350 13354
rect 30350 13302 30352 13354
rect 30296 13300 30352 13302
rect 30400 13354 30456 13356
rect 30400 13302 30402 13354
rect 30402 13302 30454 13354
rect 30454 13302 30456 13354
rect 30400 13300 30456 13302
rect 28476 13132 28532 13188
rect 28028 12738 28084 12740
rect 28028 12686 28030 12738
rect 28030 12686 28082 12738
rect 28082 12686 28084 12738
rect 28028 12684 28084 12686
rect 27916 12178 27972 12180
rect 27916 12126 27918 12178
rect 27918 12126 27970 12178
rect 27970 12126 27972 12178
rect 27916 12124 27972 12126
rect 28364 12012 28420 12068
rect 27916 11340 27972 11396
rect 28140 10780 28196 10836
rect 27020 10444 27076 10500
rect 26796 10332 26852 10388
rect 27020 9884 27076 9940
rect 25900 9266 25956 9268
rect 25900 9214 25902 9266
rect 25902 9214 25954 9266
rect 25954 9214 25956 9266
rect 25900 9212 25956 9214
rect 26124 9772 26180 9828
rect 26236 9266 26292 9268
rect 26236 9214 26238 9266
rect 26238 9214 26290 9266
rect 26290 9214 26292 9266
rect 26236 9212 26292 9214
rect 26012 9100 26068 9156
rect 26348 9154 26404 9156
rect 26348 9102 26350 9154
rect 26350 9102 26402 9154
rect 26402 9102 26404 9154
rect 26348 9100 26404 9102
rect 26908 8258 26964 8260
rect 26908 8206 26910 8258
rect 26910 8206 26962 8258
rect 26962 8206 26964 8258
rect 26908 8204 26964 8206
rect 26348 8146 26404 8148
rect 26348 8094 26350 8146
rect 26350 8094 26402 8146
rect 26402 8094 26404 8146
rect 26348 8092 26404 8094
rect 27804 9884 27860 9940
rect 28252 9772 28308 9828
rect 28140 9042 28196 9044
rect 28140 8990 28142 9042
rect 28142 8990 28194 9042
rect 28194 8990 28196 9042
rect 28140 8988 28196 8990
rect 26684 7756 26740 7812
rect 27244 8146 27300 8148
rect 27244 8094 27246 8146
rect 27246 8094 27298 8146
rect 27298 8094 27300 8146
rect 27244 8092 27300 8094
rect 25340 7308 25396 7364
rect 25116 6636 25172 6692
rect 25116 5964 25172 6020
rect 25228 6578 25284 6580
rect 25228 6526 25230 6578
rect 25230 6526 25282 6578
rect 25282 6526 25284 6578
rect 25228 6524 25284 6526
rect 25004 3500 25060 3556
rect 24780 2828 24836 2884
rect 25564 6524 25620 6580
rect 26348 7532 26404 7588
rect 26012 6636 26068 6692
rect 27692 7980 27748 8036
rect 28028 8092 28084 8148
rect 30716 13132 30772 13188
rect 29260 12796 29316 12852
rect 28588 12124 28644 12180
rect 28812 10780 28868 10836
rect 28476 10668 28532 10724
rect 28812 9884 28868 9940
rect 28476 9826 28532 9828
rect 28476 9774 28478 9826
rect 28478 9774 28530 9826
rect 28530 9774 28532 9826
rect 28476 9772 28532 9774
rect 29596 12684 29652 12740
rect 29708 12124 29764 12180
rect 29708 11900 29764 11956
rect 29596 11394 29652 11396
rect 29596 11342 29598 11394
rect 29598 11342 29650 11394
rect 29650 11342 29652 11394
rect 29596 11340 29652 11342
rect 30044 12684 30100 12740
rect 30268 12738 30324 12740
rect 30268 12686 30270 12738
rect 30270 12686 30322 12738
rect 30322 12686 30324 12738
rect 30268 12684 30324 12686
rect 30192 11786 30248 11788
rect 30192 11734 30194 11786
rect 30194 11734 30246 11786
rect 30246 11734 30248 11786
rect 30192 11732 30248 11734
rect 30296 11786 30352 11788
rect 30296 11734 30298 11786
rect 30298 11734 30350 11786
rect 30350 11734 30352 11786
rect 30296 11732 30352 11734
rect 30400 11786 30456 11788
rect 30400 11734 30402 11786
rect 30402 11734 30454 11786
rect 30454 11734 30456 11786
rect 30400 11732 30456 11734
rect 29820 10780 29876 10836
rect 29932 11004 29988 11060
rect 29820 10498 29876 10500
rect 29820 10446 29822 10498
rect 29822 10446 29874 10498
rect 29874 10446 29876 10498
rect 29820 10444 29876 10446
rect 28700 9042 28756 9044
rect 28700 8990 28702 9042
rect 28702 8990 28754 9042
rect 28754 8990 28756 9042
rect 28700 8988 28756 8990
rect 28812 8818 28868 8820
rect 28812 8766 28814 8818
rect 28814 8766 28866 8818
rect 28866 8766 28868 8818
rect 28812 8764 28868 8766
rect 28476 8204 28532 8260
rect 28812 8258 28868 8260
rect 28812 8206 28814 8258
rect 28814 8206 28866 8258
rect 28866 8206 28868 8258
rect 28812 8204 28868 8206
rect 25788 6466 25844 6468
rect 25788 6414 25790 6466
rect 25790 6414 25842 6466
rect 25842 6414 25844 6466
rect 25788 6412 25844 6414
rect 25676 5964 25732 6020
rect 25452 5180 25508 5236
rect 25452 4956 25508 5012
rect 25676 4620 25732 4676
rect 25676 4338 25732 4340
rect 25676 4286 25678 4338
rect 25678 4286 25730 4338
rect 25730 4286 25732 4338
rect 25676 4284 25732 4286
rect 26236 4732 26292 4788
rect 26124 4562 26180 4564
rect 26124 4510 26126 4562
rect 26126 4510 26178 4562
rect 26178 4510 26180 4562
rect 26124 4508 26180 4510
rect 26684 5404 26740 5460
rect 28140 6748 28196 6804
rect 28252 6972 28308 7028
rect 26012 4338 26068 4340
rect 26012 4286 26014 4338
rect 26014 4286 26066 4338
rect 26066 4286 26068 4338
rect 26012 4284 26068 4286
rect 26236 4226 26292 4228
rect 26236 4174 26238 4226
rect 26238 4174 26290 4226
rect 26290 4174 26292 4226
rect 26236 4172 26292 4174
rect 25900 3554 25956 3556
rect 25900 3502 25902 3554
rect 25902 3502 25954 3554
rect 25954 3502 25956 3554
rect 25900 3500 25956 3502
rect 25788 3276 25844 3332
rect 26124 3388 26180 3444
rect 25228 1148 25284 1204
rect 26348 3442 26404 3444
rect 26348 3390 26350 3442
rect 26350 3390 26402 3442
rect 26402 3390 26404 3442
rect 26348 3388 26404 3390
rect 27020 6188 27076 6244
rect 28140 6578 28196 6580
rect 28140 6526 28142 6578
rect 28142 6526 28194 6578
rect 28194 6526 28196 6578
rect 28140 6524 28196 6526
rect 28028 6466 28084 6468
rect 28028 6414 28030 6466
rect 28030 6414 28082 6466
rect 28082 6414 28084 6466
rect 28028 6412 28084 6414
rect 27468 5740 27524 5796
rect 27916 5404 27972 5460
rect 26460 2044 26516 2100
rect 28364 5122 28420 5124
rect 28364 5070 28366 5122
rect 28366 5070 28418 5122
rect 28418 5070 28420 5122
rect 28364 5068 28420 5070
rect 27916 4956 27972 5012
rect 28588 6972 28644 7028
rect 29484 9100 29540 9156
rect 30828 12290 30884 12292
rect 30828 12238 30830 12290
rect 30830 12238 30882 12290
rect 30882 12238 30884 12290
rect 30828 12236 30884 12238
rect 30192 10218 30248 10220
rect 30192 10166 30194 10218
rect 30194 10166 30246 10218
rect 30246 10166 30248 10218
rect 30192 10164 30248 10166
rect 30296 10218 30352 10220
rect 30296 10166 30298 10218
rect 30298 10166 30350 10218
rect 30350 10166 30352 10218
rect 30296 10164 30352 10166
rect 30400 10218 30456 10220
rect 30400 10166 30402 10218
rect 30402 10166 30454 10218
rect 30454 10166 30456 10218
rect 30400 10164 30456 10166
rect 30828 10834 30884 10836
rect 30828 10782 30830 10834
rect 30830 10782 30882 10834
rect 30882 10782 30884 10834
rect 30828 10780 30884 10782
rect 31052 10780 31108 10836
rect 32172 19010 32228 19012
rect 32172 18958 32174 19010
rect 32174 18958 32226 19010
rect 32226 18958 32228 19010
rect 32172 18956 32228 18958
rect 32172 18396 32228 18452
rect 31948 17052 32004 17108
rect 32284 18338 32340 18340
rect 32284 18286 32286 18338
rect 32286 18286 32338 18338
rect 32338 18286 32340 18338
rect 32284 18284 32340 18286
rect 32956 22370 33012 22372
rect 32956 22318 32958 22370
rect 32958 22318 33010 22370
rect 33010 22318 33012 22370
rect 32956 22316 33012 22318
rect 33964 30044 34020 30100
rect 35420 30322 35476 30324
rect 35420 30270 35422 30322
rect 35422 30270 35474 30322
rect 35474 30270 35476 30322
rect 35420 30268 35476 30270
rect 34748 30156 34804 30212
rect 35308 30210 35364 30212
rect 35308 30158 35310 30210
rect 35310 30158 35362 30210
rect 35362 30158 35364 30210
rect 35308 30156 35364 30158
rect 34076 29932 34132 29988
rect 33628 29538 33684 29540
rect 33628 29486 33630 29538
rect 33630 29486 33682 29538
rect 33682 29486 33684 29538
rect 33628 29484 33684 29486
rect 33740 28588 33796 28644
rect 33628 28530 33684 28532
rect 33628 28478 33630 28530
rect 33630 28478 33682 28530
rect 33682 28478 33684 28530
rect 33628 28476 33684 28478
rect 34636 29986 34692 29988
rect 34636 29934 34638 29986
rect 34638 29934 34690 29986
rect 34690 29934 34692 29986
rect 34636 29932 34692 29934
rect 38108 32172 38164 32228
rect 37772 32002 37828 32004
rect 37772 31950 37774 32002
rect 37774 31950 37826 32002
rect 37826 31950 37828 32002
rect 37772 31948 37828 31950
rect 38780 32172 38836 32228
rect 37884 30716 37940 30772
rect 36428 30604 36484 30660
rect 36652 30210 36708 30212
rect 36652 30158 36654 30210
rect 36654 30158 36706 30210
rect 36706 30158 36708 30210
rect 36652 30156 36708 30158
rect 37436 30210 37492 30212
rect 37436 30158 37438 30210
rect 37438 30158 37490 30210
rect 37490 30158 37492 30210
rect 37436 30156 37492 30158
rect 36092 29932 36148 29988
rect 36540 29986 36596 29988
rect 36540 29934 36542 29986
rect 36542 29934 36594 29986
rect 36594 29934 36596 29986
rect 36540 29932 36596 29934
rect 39852 31386 39908 31388
rect 39852 31334 39854 31386
rect 39854 31334 39906 31386
rect 39906 31334 39908 31386
rect 39852 31332 39908 31334
rect 39956 31386 40012 31388
rect 39956 31334 39958 31386
rect 39958 31334 40010 31386
rect 40010 31334 40012 31386
rect 39956 31332 40012 31334
rect 40060 31386 40116 31388
rect 40060 31334 40062 31386
rect 40062 31334 40114 31386
rect 40114 31334 40116 31386
rect 40060 31332 40116 31334
rect 39340 31052 39396 31108
rect 39116 30882 39172 30884
rect 39116 30830 39118 30882
rect 39118 30830 39170 30882
rect 39170 30830 39172 30882
rect 39116 30828 39172 30830
rect 39676 30940 39732 30996
rect 44716 35196 44772 35252
rect 44940 34860 44996 34916
rect 45276 36258 45332 36260
rect 45276 36206 45278 36258
rect 45278 36206 45330 36258
rect 45330 36206 45332 36258
rect 45276 36204 45332 36206
rect 45500 36092 45556 36148
rect 47180 36204 47236 36260
rect 45612 35698 45668 35700
rect 45612 35646 45614 35698
rect 45614 35646 45666 35698
rect 45666 35646 45668 35698
rect 45612 35644 45668 35646
rect 47180 35644 47236 35700
rect 46172 35420 46228 35476
rect 46508 35196 46564 35252
rect 45052 34188 45108 34244
rect 45388 34860 45444 34916
rect 46172 34860 46228 34916
rect 47180 34914 47236 34916
rect 47180 34862 47182 34914
rect 47182 34862 47234 34914
rect 47234 34862 47236 34914
rect 47180 34860 47236 34862
rect 46620 34802 46676 34804
rect 46620 34750 46622 34802
rect 46622 34750 46674 34802
rect 46674 34750 46676 34802
rect 46620 34748 46676 34750
rect 44716 33068 44772 33124
rect 44380 32956 44436 33012
rect 40460 31724 40516 31780
rect 41020 31778 41076 31780
rect 41020 31726 41022 31778
rect 41022 31726 41074 31778
rect 41074 31726 41076 31778
rect 41020 31724 41076 31726
rect 40460 31052 40516 31108
rect 42028 31106 42084 31108
rect 42028 31054 42030 31106
rect 42030 31054 42082 31106
rect 42082 31054 42084 31106
rect 42028 31052 42084 31054
rect 43596 31106 43652 31108
rect 43596 31054 43598 31106
rect 43598 31054 43650 31106
rect 43650 31054 43652 31106
rect 43596 31052 43652 31054
rect 40236 30882 40292 30884
rect 40236 30830 40238 30882
rect 40238 30830 40290 30882
rect 40290 30830 40292 30882
rect 40236 30828 40292 30830
rect 39340 30716 39396 30772
rect 39116 30268 39172 30324
rect 39004 30044 39060 30100
rect 44380 31388 44436 31444
rect 44492 32620 44548 32676
rect 47516 34802 47572 34804
rect 47516 34750 47518 34802
rect 47518 34750 47570 34802
rect 47570 34750 47572 34802
rect 47516 34748 47572 34750
rect 47180 33628 47236 33684
rect 45612 33292 45668 33348
rect 45500 33234 45556 33236
rect 45500 33182 45502 33234
rect 45502 33182 45554 33234
rect 45554 33182 45556 33234
rect 45500 33180 45556 33182
rect 45836 33234 45892 33236
rect 45836 33182 45838 33234
rect 45838 33182 45890 33234
rect 45890 33182 45892 33234
rect 45836 33180 45892 33182
rect 47852 35980 47908 36036
rect 48300 35980 48356 36036
rect 48076 35698 48132 35700
rect 48076 35646 48078 35698
rect 48078 35646 48130 35698
rect 48130 35646 48132 35698
rect 48076 35644 48132 35646
rect 48188 35196 48244 35252
rect 48524 35644 48580 35700
rect 48748 34860 48804 34916
rect 47740 34748 47796 34804
rect 48636 34802 48692 34804
rect 48636 34750 48638 34802
rect 48638 34750 48690 34802
rect 48690 34750 48692 34802
rect 48636 34748 48692 34750
rect 49756 35980 49812 36036
rect 53452 36540 53508 36596
rect 53676 37660 53732 37716
rect 54348 36594 54404 36596
rect 54348 36542 54350 36594
rect 54350 36542 54402 36594
rect 54402 36542 54404 36594
rect 54348 36540 54404 36542
rect 57708 37436 57764 37492
rect 52220 35868 52276 35924
rect 52108 35810 52164 35812
rect 52108 35758 52110 35810
rect 52110 35758 52162 35810
rect 52162 35758 52164 35810
rect 52108 35756 52164 35758
rect 51884 35532 51940 35588
rect 49308 35196 49364 35252
rect 49512 35306 49568 35308
rect 49512 35254 49514 35306
rect 49514 35254 49566 35306
rect 49566 35254 49568 35306
rect 49512 35252 49568 35254
rect 49616 35306 49672 35308
rect 49616 35254 49618 35306
rect 49618 35254 49670 35306
rect 49670 35254 49672 35306
rect 49616 35252 49672 35254
rect 49720 35306 49776 35308
rect 49720 35254 49722 35306
rect 49722 35254 49774 35306
rect 49774 35254 49776 35306
rect 49720 35252 49776 35254
rect 49756 34802 49812 34804
rect 49756 34750 49758 34802
rect 49758 34750 49810 34802
rect 49810 34750 49812 34802
rect 49756 34748 49812 34750
rect 48412 33628 48468 33684
rect 46060 33180 46116 33236
rect 44492 31276 44548 31332
rect 45388 31724 45444 31780
rect 44156 31218 44212 31220
rect 44156 31166 44158 31218
rect 44158 31166 44210 31218
rect 44210 31166 44212 31218
rect 44156 31164 44212 31166
rect 42140 30994 42196 30996
rect 42140 30942 42142 30994
rect 42142 30942 42194 30994
rect 42194 30942 42196 30994
rect 42140 30940 42196 30942
rect 41692 30098 41748 30100
rect 41692 30046 41694 30098
rect 41694 30046 41746 30098
rect 41746 30046 41748 30098
rect 41692 30044 41748 30046
rect 42140 30716 42196 30772
rect 40908 29932 40964 29988
rect 39852 29818 39908 29820
rect 39852 29766 39854 29818
rect 39854 29766 39906 29818
rect 39906 29766 39908 29818
rect 39852 29764 39908 29766
rect 39956 29818 40012 29820
rect 39956 29766 39958 29818
rect 39958 29766 40010 29818
rect 40010 29766 40012 29818
rect 39956 29764 40012 29766
rect 40060 29818 40116 29820
rect 40060 29766 40062 29818
rect 40062 29766 40114 29818
rect 40114 29766 40116 29818
rect 40060 29764 40116 29766
rect 40460 29650 40516 29652
rect 40460 29598 40462 29650
rect 40462 29598 40514 29650
rect 40514 29598 40516 29650
rect 40460 29596 40516 29598
rect 35532 29260 35588 29316
rect 35756 29148 35812 29204
rect 34300 28642 34356 28644
rect 34300 28590 34302 28642
rect 34302 28590 34354 28642
rect 34354 28590 34356 28642
rect 34300 28588 34356 28590
rect 35196 28364 35252 28420
rect 35644 28418 35700 28420
rect 35644 28366 35646 28418
rect 35646 28366 35698 28418
rect 35698 28366 35700 28418
rect 35644 28364 35700 28366
rect 36876 28642 36932 28644
rect 36876 28590 36878 28642
rect 36878 28590 36930 28642
rect 36930 28590 36932 28642
rect 36876 28588 36932 28590
rect 35756 28028 35812 28084
rect 36092 28418 36148 28420
rect 36092 28366 36094 28418
rect 36094 28366 36146 28418
rect 36146 28366 36148 28418
rect 36092 28364 36148 28366
rect 34636 27186 34692 27188
rect 34636 27134 34638 27186
rect 34638 27134 34690 27186
rect 34690 27134 34692 27186
rect 34636 27132 34692 27134
rect 33628 24556 33684 24612
rect 34300 26460 34356 26516
rect 32844 17500 32900 17556
rect 33180 20076 33236 20132
rect 32844 17276 32900 17332
rect 32732 17164 32788 17220
rect 31836 16940 31892 16996
rect 31724 16268 31780 16324
rect 31724 15820 31780 15876
rect 31948 16098 32004 16100
rect 31948 16046 31950 16098
rect 31950 16046 32002 16098
rect 32002 16046 32004 16098
rect 31948 16044 32004 16046
rect 32172 16044 32228 16100
rect 32060 15932 32116 15988
rect 32508 16994 32564 16996
rect 32508 16942 32510 16994
rect 32510 16942 32562 16994
rect 32562 16942 32564 16994
rect 32508 16940 32564 16942
rect 32844 16828 32900 16884
rect 32732 16604 32788 16660
rect 32396 15932 32452 15988
rect 32620 15986 32676 15988
rect 32620 15934 32622 15986
rect 32622 15934 32674 15986
rect 32674 15934 32676 15986
rect 32620 15932 32676 15934
rect 32508 15820 32564 15876
rect 32396 15708 32452 15764
rect 31948 15372 32004 15428
rect 31836 15314 31892 15316
rect 31836 15262 31838 15314
rect 31838 15262 31890 15314
rect 31890 15262 31892 15314
rect 31836 15260 31892 15262
rect 32172 15202 32228 15204
rect 32172 15150 32174 15202
rect 32174 15150 32226 15202
rect 32226 15150 32228 15202
rect 32172 15148 32228 15150
rect 32396 14700 32452 14756
rect 32620 13692 32676 13748
rect 31500 12738 31556 12740
rect 31500 12686 31502 12738
rect 31502 12686 31554 12738
rect 31554 12686 31556 12738
rect 31500 12684 31556 12686
rect 32732 13468 32788 13524
rect 32172 12684 32228 12740
rect 31500 12124 31556 12180
rect 31836 10780 31892 10836
rect 30268 9938 30324 9940
rect 30268 9886 30270 9938
rect 30270 9886 30322 9938
rect 30322 9886 30324 9938
rect 30268 9884 30324 9886
rect 31276 10556 31332 10612
rect 30940 9938 30996 9940
rect 30940 9886 30942 9938
rect 30942 9886 30994 9938
rect 30994 9886 30996 9938
rect 30940 9884 30996 9886
rect 29708 9212 29764 9268
rect 32284 10668 32340 10724
rect 32396 10610 32452 10612
rect 32396 10558 32398 10610
rect 32398 10558 32450 10610
rect 32450 10558 32452 10610
rect 32396 10556 32452 10558
rect 32844 12572 32900 12628
rect 33628 23660 33684 23716
rect 33292 17164 33348 17220
rect 33516 19516 33572 19572
rect 33516 18956 33572 19012
rect 34300 26012 34356 26068
rect 33852 25340 33908 25396
rect 34300 25506 34356 25508
rect 34300 25454 34302 25506
rect 34302 25454 34354 25506
rect 34354 25454 34356 25506
rect 34300 25452 34356 25454
rect 33852 24722 33908 24724
rect 33852 24670 33854 24722
rect 33854 24670 33906 24722
rect 33906 24670 33908 24722
rect 33852 24668 33908 24670
rect 34076 24668 34132 24724
rect 34524 24722 34580 24724
rect 34524 24670 34526 24722
rect 34526 24670 34578 24722
rect 34578 24670 34580 24722
rect 34524 24668 34580 24670
rect 34636 24610 34692 24612
rect 34636 24558 34638 24610
rect 34638 24558 34690 24610
rect 34690 24558 34692 24610
rect 34636 24556 34692 24558
rect 33964 23938 34020 23940
rect 33964 23886 33966 23938
rect 33966 23886 34018 23938
rect 34018 23886 34020 23938
rect 33964 23884 34020 23886
rect 34636 23938 34692 23940
rect 34636 23886 34638 23938
rect 34638 23886 34690 23938
rect 34690 23886 34692 23938
rect 34636 23884 34692 23886
rect 34748 23714 34804 23716
rect 34748 23662 34750 23714
rect 34750 23662 34802 23714
rect 34802 23662 34804 23714
rect 34748 23660 34804 23662
rect 34972 23714 35028 23716
rect 34972 23662 34974 23714
rect 34974 23662 35026 23714
rect 35026 23662 35028 23714
rect 34972 23660 35028 23662
rect 33740 22540 33796 22596
rect 34076 23154 34132 23156
rect 34076 23102 34078 23154
rect 34078 23102 34130 23154
rect 34130 23102 34132 23154
rect 34076 23100 34132 23102
rect 34076 22370 34132 22372
rect 34076 22318 34078 22370
rect 34078 22318 34130 22370
rect 34130 22318 34132 22370
rect 34076 22316 34132 22318
rect 33964 21644 34020 21700
rect 34972 21026 35028 21028
rect 34972 20974 34974 21026
rect 34974 20974 35026 21026
rect 35026 20974 35028 21026
rect 34972 20972 35028 20974
rect 33740 19628 33796 19684
rect 35532 27746 35588 27748
rect 35532 27694 35534 27746
rect 35534 27694 35586 27746
rect 35586 27694 35588 27746
rect 35532 27692 35588 27694
rect 36652 28418 36708 28420
rect 36652 28366 36654 28418
rect 36654 28366 36706 28418
rect 36706 28366 36708 28418
rect 36652 28364 36708 28366
rect 37100 28364 37156 28420
rect 36428 28252 36484 28308
rect 36092 27692 36148 27748
rect 36316 27692 36372 27748
rect 36316 27298 36372 27300
rect 36316 27246 36318 27298
rect 36318 27246 36370 27298
rect 36370 27246 36372 27298
rect 36316 27244 36372 27246
rect 37996 29260 38052 29316
rect 37436 28642 37492 28644
rect 37436 28590 37438 28642
rect 37438 28590 37490 28642
rect 37490 28590 37492 28642
rect 37436 28588 37492 28590
rect 39116 29314 39172 29316
rect 39116 29262 39118 29314
rect 39118 29262 39170 29314
rect 39170 29262 39172 29314
rect 39116 29260 39172 29262
rect 40572 29426 40628 29428
rect 40572 29374 40574 29426
rect 40574 29374 40626 29426
rect 40626 29374 40628 29426
rect 40572 29372 40628 29374
rect 38556 29148 38612 29204
rect 38108 28418 38164 28420
rect 38108 28366 38110 28418
rect 38110 28366 38162 28418
rect 38162 28366 38164 28418
rect 38108 28364 38164 28366
rect 39340 29202 39396 29204
rect 39340 29150 39342 29202
rect 39342 29150 39394 29202
rect 39394 29150 39396 29202
rect 39340 29148 39396 29150
rect 40796 29372 40852 29428
rect 39340 28700 39396 28756
rect 40012 28754 40068 28756
rect 40012 28702 40014 28754
rect 40014 28702 40066 28754
rect 40066 28702 40068 28754
rect 40012 28700 40068 28702
rect 40236 28476 40292 28532
rect 39852 28250 39908 28252
rect 39852 28198 39854 28250
rect 39854 28198 39906 28250
rect 39906 28198 39908 28250
rect 39852 28196 39908 28198
rect 39956 28250 40012 28252
rect 39956 28198 39958 28250
rect 39958 28198 40010 28250
rect 40010 28198 40012 28250
rect 39956 28196 40012 28198
rect 40060 28250 40116 28252
rect 40060 28198 40062 28250
rect 40062 28198 40114 28250
rect 40114 28198 40116 28250
rect 40060 28196 40116 28198
rect 37100 27244 37156 27300
rect 35644 26236 35700 26292
rect 36652 26796 36708 26852
rect 36540 26514 36596 26516
rect 36540 26462 36542 26514
rect 36542 26462 36594 26514
rect 36594 26462 36596 26514
rect 36540 26460 36596 26462
rect 36204 26290 36260 26292
rect 36204 26238 36206 26290
rect 36206 26238 36258 26290
rect 36258 26238 36260 26290
rect 36204 26236 36260 26238
rect 35980 26178 36036 26180
rect 35980 26126 35982 26178
rect 35982 26126 36034 26178
rect 36034 26126 36036 26178
rect 35980 26124 36036 26126
rect 35420 24834 35476 24836
rect 35420 24782 35422 24834
rect 35422 24782 35474 24834
rect 35474 24782 35476 24834
rect 35420 24780 35476 24782
rect 35308 24722 35364 24724
rect 35308 24670 35310 24722
rect 35310 24670 35362 24722
rect 35362 24670 35364 24722
rect 35308 24668 35364 24670
rect 35756 24220 35812 24276
rect 35532 23714 35588 23716
rect 35532 23662 35534 23714
rect 35534 23662 35586 23714
rect 35586 23662 35588 23714
rect 35532 23660 35588 23662
rect 36204 23042 36260 23044
rect 36204 22990 36206 23042
rect 36206 22990 36258 23042
rect 36258 22990 36260 23042
rect 36204 22988 36260 22990
rect 39228 27244 39284 27300
rect 38556 27074 38612 27076
rect 38556 27022 38558 27074
rect 38558 27022 38610 27074
rect 38610 27022 38612 27074
rect 38556 27020 38612 27022
rect 39004 27020 39060 27076
rect 38668 26684 38724 26740
rect 38332 26290 38388 26292
rect 38332 26238 38334 26290
rect 38334 26238 38386 26290
rect 38386 26238 38388 26290
rect 38332 26236 38388 26238
rect 38332 26066 38388 26068
rect 38332 26014 38334 26066
rect 38334 26014 38386 26066
rect 38386 26014 38388 26066
rect 38332 26012 38388 26014
rect 38668 25788 38724 25844
rect 39900 27580 39956 27636
rect 39676 27298 39732 27300
rect 39676 27246 39678 27298
rect 39678 27246 39730 27298
rect 39730 27246 39732 27298
rect 39676 27244 39732 27246
rect 40124 27692 40180 27748
rect 40124 27244 40180 27300
rect 39900 27132 39956 27188
rect 39788 27074 39844 27076
rect 39788 27022 39790 27074
rect 39790 27022 39842 27074
rect 39842 27022 39844 27074
rect 39788 27020 39844 27022
rect 39116 26684 39172 26740
rect 39676 26796 39732 26852
rect 39564 26572 39620 26628
rect 39452 26178 39508 26180
rect 39452 26126 39454 26178
rect 39454 26126 39506 26178
rect 39506 26126 39508 26178
rect 39452 26124 39508 26126
rect 39116 25452 39172 25508
rect 39340 25452 39396 25508
rect 37100 24556 37156 24612
rect 37996 24556 38052 24612
rect 36876 23714 36932 23716
rect 36876 23662 36878 23714
rect 36878 23662 36930 23714
rect 36930 23662 36932 23714
rect 36876 23660 36932 23662
rect 36764 22988 36820 23044
rect 36204 21980 36260 22036
rect 35756 21698 35812 21700
rect 35756 21646 35758 21698
rect 35758 21646 35810 21698
rect 35810 21646 35812 21698
rect 35756 21644 35812 21646
rect 35196 20076 35252 20132
rect 35868 20524 35924 20580
rect 34636 19852 34692 19908
rect 35196 19906 35252 19908
rect 35196 19854 35198 19906
rect 35198 19854 35250 19906
rect 35250 19854 35252 19906
rect 35196 19852 35252 19854
rect 34076 19234 34132 19236
rect 34076 19182 34078 19234
rect 34078 19182 34130 19234
rect 34130 19182 34132 19234
rect 34076 19180 34132 19182
rect 33852 18620 33908 18676
rect 35308 19628 35364 19684
rect 35532 19628 35588 19684
rect 34636 19180 34692 19236
rect 34748 19122 34804 19124
rect 34748 19070 34750 19122
rect 34750 19070 34802 19122
rect 34802 19070 34804 19122
rect 34748 19068 34804 19070
rect 34748 18508 34804 18564
rect 33628 18172 33684 18228
rect 33628 17778 33684 17780
rect 33628 17726 33630 17778
rect 33630 17726 33682 17778
rect 33682 17726 33684 17778
rect 33628 17724 33684 17726
rect 33516 17276 33572 17332
rect 34188 18060 34244 18116
rect 34524 17778 34580 17780
rect 34524 17726 34526 17778
rect 34526 17726 34578 17778
rect 34578 17726 34580 17778
rect 34524 17724 34580 17726
rect 33516 15986 33572 15988
rect 33516 15934 33518 15986
rect 33518 15934 33570 15986
rect 33570 15934 33572 15986
rect 33516 15932 33572 15934
rect 33740 15874 33796 15876
rect 33740 15822 33742 15874
rect 33742 15822 33794 15874
rect 33794 15822 33796 15874
rect 33740 15820 33796 15822
rect 34412 15986 34468 15988
rect 34412 15934 34414 15986
rect 34414 15934 34466 15986
rect 34466 15934 34468 15986
rect 34412 15932 34468 15934
rect 34524 15874 34580 15876
rect 34524 15822 34526 15874
rect 34526 15822 34578 15874
rect 34578 15822 34580 15874
rect 34524 15820 34580 15822
rect 34300 15708 34356 15764
rect 33628 14476 33684 14532
rect 33852 15036 33908 15092
rect 33404 13804 33460 13860
rect 33180 12236 33236 12292
rect 33404 12012 33460 12068
rect 32844 10444 32900 10500
rect 33180 10444 33236 10500
rect 32956 10220 33012 10276
rect 32284 9212 32340 9268
rect 32844 9884 32900 9940
rect 30044 9100 30100 9156
rect 29932 8988 29988 9044
rect 29596 8316 29652 8372
rect 29708 8764 29764 8820
rect 29484 7532 29540 7588
rect 30604 9154 30660 9156
rect 30604 9102 30606 9154
rect 30606 9102 30658 9154
rect 30658 9102 30660 9154
rect 30604 9100 30660 9102
rect 30492 9042 30548 9044
rect 30492 8990 30494 9042
rect 30494 8990 30546 9042
rect 30546 8990 30548 9042
rect 30492 8988 30548 8990
rect 31500 9042 31556 9044
rect 31500 8990 31502 9042
rect 31502 8990 31554 9042
rect 31554 8990 31556 9042
rect 31500 8988 31556 8990
rect 30192 8650 30248 8652
rect 30192 8598 30194 8650
rect 30194 8598 30246 8650
rect 30246 8598 30248 8650
rect 30192 8596 30248 8598
rect 30296 8650 30352 8652
rect 30296 8598 30298 8650
rect 30298 8598 30350 8650
rect 30350 8598 30352 8650
rect 30296 8596 30352 8598
rect 30400 8650 30456 8652
rect 30400 8598 30402 8650
rect 30402 8598 30454 8650
rect 30454 8598 30456 8650
rect 30400 8596 30456 8598
rect 31388 8258 31444 8260
rect 31388 8206 31390 8258
rect 31390 8206 31442 8258
rect 31442 8206 31444 8258
rect 31388 8204 31444 8206
rect 31724 8204 31780 8260
rect 31612 8092 31668 8148
rect 29820 7532 29876 7588
rect 31164 7420 31220 7476
rect 30940 7362 30996 7364
rect 30940 7310 30942 7362
rect 30942 7310 30994 7362
rect 30994 7310 30996 7362
rect 30940 7308 30996 7310
rect 30192 7082 30248 7084
rect 30192 7030 30194 7082
rect 30194 7030 30246 7082
rect 30246 7030 30248 7082
rect 30192 7028 30248 7030
rect 30296 7082 30352 7084
rect 30296 7030 30298 7082
rect 30298 7030 30350 7082
rect 30350 7030 30352 7082
rect 30296 7028 30352 7030
rect 30400 7082 30456 7084
rect 30400 7030 30402 7082
rect 30402 7030 30454 7082
rect 30454 7030 30456 7082
rect 30400 7028 30456 7030
rect 28924 6748 28980 6804
rect 29484 6802 29540 6804
rect 29484 6750 29486 6802
rect 29486 6750 29538 6802
rect 29538 6750 29540 6802
rect 29484 6748 29540 6750
rect 28812 6636 28868 6692
rect 27692 4732 27748 4788
rect 27244 4620 27300 4676
rect 28140 4732 28196 4788
rect 27804 4620 27860 4676
rect 27356 4338 27412 4340
rect 27356 4286 27358 4338
rect 27358 4286 27410 4338
rect 27410 4286 27412 4338
rect 27356 4284 27412 4286
rect 27020 4060 27076 4116
rect 27804 3948 27860 4004
rect 27132 2940 27188 2996
rect 27244 1484 27300 1540
rect 28252 3500 28308 3556
rect 26908 1260 26964 1316
rect 28364 3276 28420 3332
rect 28588 3442 28644 3444
rect 28588 3390 28590 3442
rect 28590 3390 28642 3442
rect 28642 3390 28644 3442
rect 28588 3388 28644 3390
rect 28476 3164 28532 3220
rect 29708 5852 29764 5908
rect 29708 5404 29764 5460
rect 28924 4956 28980 5012
rect 29148 5068 29204 5124
rect 29260 3554 29316 3556
rect 29260 3502 29262 3554
rect 29262 3502 29314 3554
rect 29314 3502 29316 3554
rect 29260 3500 29316 3502
rect 29596 3330 29652 3332
rect 29596 3278 29598 3330
rect 29598 3278 29650 3330
rect 29650 3278 29652 3330
rect 29596 3276 29652 3278
rect 29820 5180 29876 5236
rect 30604 6300 30660 6356
rect 30044 5906 30100 5908
rect 30044 5854 30046 5906
rect 30046 5854 30098 5906
rect 30098 5854 30100 5906
rect 30044 5852 30100 5854
rect 30380 5794 30436 5796
rect 30380 5742 30382 5794
rect 30382 5742 30434 5794
rect 30434 5742 30436 5794
rect 30380 5740 30436 5742
rect 30192 5514 30248 5516
rect 30192 5462 30194 5514
rect 30194 5462 30246 5514
rect 30246 5462 30248 5514
rect 30192 5460 30248 5462
rect 30296 5514 30352 5516
rect 30296 5462 30298 5514
rect 30298 5462 30350 5514
rect 30350 5462 30352 5514
rect 30296 5460 30352 5462
rect 30400 5514 30456 5516
rect 30400 5462 30402 5514
rect 30402 5462 30454 5514
rect 30454 5462 30456 5514
rect 30400 5460 30456 5462
rect 29932 4396 29988 4452
rect 30044 5180 30100 5236
rect 30492 5122 30548 5124
rect 30492 5070 30494 5122
rect 30494 5070 30546 5122
rect 30546 5070 30548 5122
rect 30492 5068 30548 5070
rect 30156 4396 30212 4452
rect 31500 6748 31556 6804
rect 32732 9266 32788 9268
rect 32732 9214 32734 9266
rect 32734 9214 32786 9266
rect 32786 9214 32788 9266
rect 32732 9212 32788 9214
rect 32844 8540 32900 8596
rect 32620 7474 32676 7476
rect 32620 7422 32622 7474
rect 32622 7422 32674 7474
rect 32674 7422 32676 7474
rect 32620 7420 32676 7422
rect 32060 6802 32116 6804
rect 32060 6750 32062 6802
rect 32062 6750 32114 6802
rect 32114 6750 32116 6802
rect 32060 6748 32116 6750
rect 31612 6636 31668 6692
rect 32396 6690 32452 6692
rect 32396 6638 32398 6690
rect 32398 6638 32450 6690
rect 32450 6638 32452 6690
rect 32396 6636 32452 6638
rect 31052 6578 31108 6580
rect 31052 6526 31054 6578
rect 31054 6526 31106 6578
rect 31106 6526 31108 6578
rect 31052 6524 31108 6526
rect 32060 6524 32116 6580
rect 30940 5906 30996 5908
rect 30940 5854 30942 5906
rect 30942 5854 30994 5906
rect 30994 5854 30996 5906
rect 30940 5852 30996 5854
rect 32732 5906 32788 5908
rect 32732 5854 32734 5906
rect 32734 5854 32786 5906
rect 32786 5854 32788 5906
rect 32732 5852 32788 5854
rect 30828 5010 30884 5012
rect 30828 4958 30830 5010
rect 30830 4958 30882 5010
rect 30882 4958 30884 5010
rect 30828 4956 30884 4958
rect 30716 4732 30772 4788
rect 30192 3946 30248 3948
rect 30192 3894 30194 3946
rect 30194 3894 30246 3946
rect 30246 3894 30248 3946
rect 30192 3892 30248 3894
rect 30296 3946 30352 3948
rect 30296 3894 30298 3946
rect 30298 3894 30350 3946
rect 30350 3894 30352 3946
rect 30296 3892 30352 3894
rect 30400 3946 30456 3948
rect 30400 3894 30402 3946
rect 30402 3894 30454 3946
rect 30454 3894 30456 3946
rect 30400 3892 30456 3894
rect 30044 3724 30100 3780
rect 29820 2492 29876 2548
rect 30156 3666 30212 3668
rect 30156 3614 30158 3666
rect 30158 3614 30210 3666
rect 30210 3614 30212 3666
rect 30156 3612 30212 3614
rect 30156 2380 30212 2436
rect 30604 3442 30660 3444
rect 30604 3390 30606 3442
rect 30606 3390 30658 3442
rect 30658 3390 30660 3442
rect 30604 3388 30660 3390
rect 29708 2268 29764 2324
rect 32284 5234 32340 5236
rect 32284 5182 32286 5234
rect 32286 5182 32338 5234
rect 32338 5182 32340 5234
rect 32284 5180 32340 5182
rect 33068 8540 33124 8596
rect 33404 10332 33460 10388
rect 35308 18060 35364 18116
rect 35196 17724 35252 17780
rect 34972 17052 35028 17108
rect 35196 17164 35252 17220
rect 34972 16268 35028 16324
rect 35420 16156 35476 16212
rect 36204 20860 36260 20916
rect 36764 22146 36820 22148
rect 36764 22094 36766 22146
rect 36766 22094 36818 22146
rect 36818 22094 36820 22146
rect 36764 22092 36820 22094
rect 36316 21420 36372 21476
rect 36092 20636 36148 20692
rect 36092 19628 36148 19684
rect 36652 21980 36708 22036
rect 35980 19068 36036 19124
rect 34412 14700 34468 14756
rect 34860 14812 34916 14868
rect 33964 14476 34020 14532
rect 34076 13634 34132 13636
rect 34076 13582 34078 13634
rect 34078 13582 34130 13634
rect 34130 13582 34132 13634
rect 34076 13580 34132 13582
rect 34748 14252 34804 14308
rect 34972 14530 35028 14532
rect 34972 14478 34974 14530
rect 34974 14478 35026 14530
rect 35026 14478 35028 14530
rect 34972 14476 35028 14478
rect 35644 18172 35700 18228
rect 35308 14306 35364 14308
rect 35308 14254 35310 14306
rect 35310 14254 35362 14306
rect 35362 14254 35364 14306
rect 35308 14252 35364 14254
rect 34860 13746 34916 13748
rect 34860 13694 34862 13746
rect 34862 13694 34914 13746
rect 34914 13694 34916 13746
rect 34860 13692 34916 13694
rect 35308 13746 35364 13748
rect 35308 13694 35310 13746
rect 35310 13694 35362 13746
rect 35362 13694 35364 13746
rect 35308 13692 35364 13694
rect 34636 13580 34692 13636
rect 34076 12684 34132 12740
rect 34748 12290 34804 12292
rect 34748 12238 34750 12290
rect 34750 12238 34802 12290
rect 34802 12238 34804 12290
rect 34748 12236 34804 12238
rect 34300 11506 34356 11508
rect 34300 11454 34302 11506
rect 34302 11454 34354 11506
rect 34354 11454 34356 11506
rect 34300 11452 34356 11454
rect 36540 21532 36596 21588
rect 36652 20972 36708 21028
rect 36428 18844 36484 18900
rect 36652 18674 36708 18676
rect 36652 18622 36654 18674
rect 36654 18622 36706 18674
rect 36706 18622 36708 18674
rect 36652 18620 36708 18622
rect 36540 17724 36596 17780
rect 36764 17666 36820 17668
rect 36764 17614 36766 17666
rect 36766 17614 36818 17666
rect 36818 17614 36820 17666
rect 36764 17612 36820 17614
rect 35868 16882 35924 16884
rect 35868 16830 35870 16882
rect 35870 16830 35922 16882
rect 35922 16830 35924 16882
rect 35868 16828 35924 16830
rect 35868 16210 35924 16212
rect 35868 16158 35870 16210
rect 35870 16158 35922 16210
rect 35922 16158 35924 16210
rect 35868 16156 35924 16158
rect 35756 14812 35812 14868
rect 35644 14700 35700 14756
rect 35980 14476 36036 14532
rect 35756 13634 35812 13636
rect 35756 13582 35758 13634
rect 35758 13582 35810 13634
rect 35810 13582 35812 13634
rect 35756 13580 35812 13582
rect 35644 13244 35700 13300
rect 35532 12738 35588 12740
rect 35532 12686 35534 12738
rect 35534 12686 35586 12738
rect 35586 12686 35588 12738
rect 35532 12684 35588 12686
rect 35532 11900 35588 11956
rect 35420 11676 35476 11732
rect 33964 10498 34020 10500
rect 33964 10446 33966 10498
rect 33966 10446 34018 10498
rect 34018 10446 34020 10498
rect 33964 10444 34020 10446
rect 31164 4844 31220 4900
rect 31948 4898 32004 4900
rect 31948 4846 31950 4898
rect 31950 4846 32002 4898
rect 32002 4846 32004 4898
rect 31948 4844 32004 4846
rect 32172 4844 32228 4900
rect 31388 4732 31444 4788
rect 31276 4562 31332 4564
rect 31276 4510 31278 4562
rect 31278 4510 31330 4562
rect 31330 4510 31332 4562
rect 31276 4508 31332 4510
rect 31388 4172 31444 4228
rect 31948 4508 32004 4564
rect 33068 4898 33124 4900
rect 33068 4846 33070 4898
rect 33070 4846 33122 4898
rect 33122 4846 33124 4898
rect 33068 4844 33124 4846
rect 34076 9212 34132 9268
rect 34188 10444 34244 10500
rect 35532 11564 35588 11620
rect 34972 11170 35028 11172
rect 34972 11118 34974 11170
rect 34974 11118 35026 11170
rect 35026 11118 35028 11170
rect 34972 11116 35028 11118
rect 35980 12796 36036 12852
rect 35980 12066 36036 12068
rect 35980 12014 35982 12066
rect 35982 12014 36034 12066
rect 36034 12014 36036 12066
rect 35980 12012 36036 12014
rect 35644 11170 35700 11172
rect 35644 11118 35646 11170
rect 35646 11118 35698 11170
rect 35698 11118 35700 11170
rect 35644 11116 35700 11118
rect 34972 10668 35028 10724
rect 35420 10610 35476 10612
rect 35420 10558 35422 10610
rect 35422 10558 35474 10610
rect 35474 10558 35476 10610
rect 35420 10556 35476 10558
rect 37772 23714 37828 23716
rect 37772 23662 37774 23714
rect 37774 23662 37826 23714
rect 37826 23662 37828 23714
rect 37772 23660 37828 23662
rect 38108 24050 38164 24052
rect 38108 23998 38110 24050
rect 38110 23998 38162 24050
rect 38162 23998 38164 24050
rect 38108 23996 38164 23998
rect 39228 25228 39284 25284
rect 37212 23212 37268 23268
rect 36988 22092 37044 22148
rect 37660 22092 37716 22148
rect 37996 22092 38052 22148
rect 37884 21698 37940 21700
rect 37884 21646 37886 21698
rect 37886 21646 37938 21698
rect 37938 21646 37940 21698
rect 37884 21644 37940 21646
rect 37772 21586 37828 21588
rect 37772 21534 37774 21586
rect 37774 21534 37826 21586
rect 37826 21534 37828 21586
rect 37772 21532 37828 21534
rect 37324 21420 37380 21476
rect 38108 20914 38164 20916
rect 38108 20862 38110 20914
rect 38110 20862 38162 20914
rect 38162 20862 38164 20914
rect 38108 20860 38164 20862
rect 37772 20412 37828 20468
rect 38892 23996 38948 24052
rect 38668 23154 38724 23156
rect 38668 23102 38670 23154
rect 38670 23102 38722 23154
rect 38722 23102 38724 23154
rect 38668 23100 38724 23102
rect 38444 22092 38500 22148
rect 39564 25788 39620 25844
rect 39900 26796 39956 26852
rect 39852 26682 39908 26684
rect 39852 26630 39854 26682
rect 39854 26630 39906 26682
rect 39906 26630 39908 26682
rect 39852 26628 39908 26630
rect 39956 26682 40012 26684
rect 39956 26630 39958 26682
rect 39958 26630 40010 26682
rect 40010 26630 40012 26682
rect 39956 26628 40012 26630
rect 40060 26682 40116 26684
rect 40060 26630 40062 26682
rect 40062 26630 40114 26682
rect 40114 26630 40116 26682
rect 40060 26628 40116 26630
rect 39900 26348 39956 26404
rect 39788 26236 39844 26292
rect 41356 29986 41412 29988
rect 41356 29934 41358 29986
rect 41358 29934 41410 29986
rect 41410 29934 41412 29986
rect 41356 29932 41412 29934
rect 41804 29426 41860 29428
rect 41804 29374 41806 29426
rect 41806 29374 41858 29426
rect 41858 29374 41860 29426
rect 41804 29372 41860 29374
rect 40908 28700 40964 28756
rect 41132 29260 41188 29316
rect 41692 29314 41748 29316
rect 41692 29262 41694 29314
rect 41694 29262 41746 29314
rect 41746 29262 41748 29314
rect 41692 29260 41748 29262
rect 43148 29932 43204 29988
rect 45388 30716 45444 30772
rect 44716 30156 44772 30212
rect 44380 28476 44436 28532
rect 44492 29820 44548 29876
rect 41580 27746 41636 27748
rect 41580 27694 41582 27746
rect 41582 27694 41634 27746
rect 41634 27694 41636 27746
rect 41580 27692 41636 27694
rect 41804 27634 41860 27636
rect 41804 27582 41806 27634
rect 41806 27582 41858 27634
rect 41858 27582 41860 27634
rect 41804 27580 41860 27582
rect 41692 27468 41748 27524
rect 40796 27132 40852 27188
rect 40348 25788 40404 25844
rect 39900 25506 39956 25508
rect 39900 25454 39902 25506
rect 39902 25454 39954 25506
rect 39954 25454 39956 25506
rect 39900 25452 39956 25454
rect 40124 25506 40180 25508
rect 40124 25454 40126 25506
rect 40126 25454 40178 25506
rect 40178 25454 40180 25506
rect 40124 25452 40180 25454
rect 39676 25340 39732 25396
rect 41244 27132 41300 27188
rect 42252 27356 42308 27412
rect 42140 27186 42196 27188
rect 42140 27134 42142 27186
rect 42142 27134 42194 27186
rect 42194 27134 42196 27186
rect 42140 27132 42196 27134
rect 41692 26850 41748 26852
rect 41692 26798 41694 26850
rect 41694 26798 41746 26850
rect 41746 26798 41748 26850
rect 41692 26796 41748 26798
rect 41916 26402 41972 26404
rect 41916 26350 41918 26402
rect 41918 26350 41970 26402
rect 41970 26350 41972 26402
rect 41916 26348 41972 26350
rect 40796 25452 40852 25508
rect 39852 25114 39908 25116
rect 39852 25062 39854 25114
rect 39854 25062 39906 25114
rect 39906 25062 39908 25114
rect 39852 25060 39908 25062
rect 39956 25114 40012 25116
rect 39956 25062 39958 25114
rect 39958 25062 40010 25114
rect 40010 25062 40012 25114
rect 39956 25060 40012 25062
rect 40060 25114 40116 25116
rect 40060 25062 40062 25114
rect 40062 25062 40114 25114
rect 40114 25062 40116 25114
rect 40060 25060 40116 25062
rect 41244 25394 41300 25396
rect 41244 25342 41246 25394
rect 41246 25342 41298 25394
rect 41298 25342 41300 25394
rect 41244 25340 41300 25342
rect 42028 26290 42084 26292
rect 42028 26238 42030 26290
rect 42030 26238 42082 26290
rect 42082 26238 42084 26290
rect 42028 26236 42084 26238
rect 42140 26124 42196 26180
rect 41468 25228 41524 25284
rect 42028 25228 42084 25284
rect 39852 23546 39908 23548
rect 39852 23494 39854 23546
rect 39854 23494 39906 23546
rect 39906 23494 39908 23546
rect 39852 23492 39908 23494
rect 39956 23546 40012 23548
rect 39956 23494 39958 23546
rect 39958 23494 40010 23546
rect 40010 23494 40012 23546
rect 39956 23492 40012 23494
rect 40060 23546 40116 23548
rect 40060 23494 40062 23546
rect 40062 23494 40114 23546
rect 40114 23494 40116 23546
rect 40060 23492 40116 23494
rect 39564 23154 39620 23156
rect 39564 23102 39566 23154
rect 39566 23102 39618 23154
rect 39618 23102 39620 23154
rect 39564 23100 39620 23102
rect 41132 23826 41188 23828
rect 41132 23774 41134 23826
rect 41134 23774 41186 23826
rect 41186 23774 41188 23826
rect 41132 23772 41188 23774
rect 41692 23660 41748 23716
rect 42140 23714 42196 23716
rect 42140 23662 42142 23714
rect 42142 23662 42194 23714
rect 42194 23662 42196 23714
rect 42140 23660 42196 23662
rect 44604 29596 44660 29652
rect 45276 29596 45332 29652
rect 46508 32508 46564 32564
rect 46620 31724 46676 31780
rect 46956 31724 47012 31780
rect 46844 31666 46900 31668
rect 46844 31614 46846 31666
rect 46846 31614 46898 31666
rect 46898 31614 46900 31666
rect 46844 31612 46900 31614
rect 46396 31164 46452 31220
rect 45948 30716 46004 30772
rect 46172 30882 46228 30884
rect 46172 30830 46174 30882
rect 46174 30830 46226 30882
rect 46226 30830 46228 30882
rect 46172 30828 46228 30830
rect 45500 29484 45556 29540
rect 47292 31666 47348 31668
rect 47292 31614 47294 31666
rect 47294 31614 47346 31666
rect 47346 31614 47348 31666
rect 47292 31612 47348 31614
rect 46956 30828 47012 30884
rect 46060 30210 46116 30212
rect 46060 30158 46062 30210
rect 46062 30158 46114 30210
rect 46114 30158 46116 30210
rect 46060 30156 46116 30158
rect 47180 30098 47236 30100
rect 47180 30046 47182 30098
rect 47182 30046 47234 30098
rect 47234 30046 47236 30098
rect 47180 30044 47236 30046
rect 45052 28476 45108 28532
rect 45388 28700 45444 28756
rect 46508 29538 46564 29540
rect 46508 29486 46510 29538
rect 46510 29486 46562 29538
rect 46562 29486 46564 29538
rect 46508 29484 46564 29486
rect 46844 29426 46900 29428
rect 46844 29374 46846 29426
rect 46846 29374 46898 29426
rect 46898 29374 46900 29426
rect 46844 29372 46900 29374
rect 45052 27916 45108 27972
rect 45276 27858 45332 27860
rect 45276 27806 45278 27858
rect 45278 27806 45330 27858
rect 45330 27806 45332 27858
rect 45276 27804 45332 27806
rect 46396 28588 46452 28644
rect 46620 28700 46676 28756
rect 47292 28140 47348 28196
rect 45724 27916 45780 27972
rect 45500 27804 45556 27860
rect 44492 27132 44548 27188
rect 44716 27186 44772 27188
rect 44716 27134 44718 27186
rect 44718 27134 44770 27186
rect 44770 27134 44772 27186
rect 44716 27132 44772 27134
rect 45500 27132 45556 27188
rect 43260 26684 43316 26740
rect 43148 26514 43204 26516
rect 43148 26462 43150 26514
rect 43150 26462 43202 26514
rect 43202 26462 43204 26514
rect 43148 26460 43204 26462
rect 42364 24220 42420 24276
rect 42700 23772 42756 23828
rect 42252 23324 42308 23380
rect 40236 23154 40292 23156
rect 40236 23102 40238 23154
rect 40238 23102 40290 23154
rect 40290 23102 40292 23154
rect 40236 23100 40292 23102
rect 40908 23100 40964 23156
rect 40572 22652 40628 22708
rect 40348 22316 40404 22372
rect 39852 21978 39908 21980
rect 39852 21926 39854 21978
rect 39854 21926 39906 21978
rect 39906 21926 39908 21978
rect 39852 21924 39908 21926
rect 39956 21978 40012 21980
rect 39956 21926 39958 21978
rect 39958 21926 40010 21978
rect 40010 21926 40012 21978
rect 39956 21924 40012 21926
rect 40060 21978 40116 21980
rect 40060 21926 40062 21978
rect 40062 21926 40114 21978
rect 40114 21926 40116 21978
rect 40060 21924 40116 21926
rect 38668 20860 38724 20916
rect 39228 20914 39284 20916
rect 39228 20862 39230 20914
rect 39230 20862 39282 20914
rect 39282 20862 39284 20914
rect 39228 20860 39284 20862
rect 37100 19628 37156 19684
rect 38108 20076 38164 20132
rect 37100 18620 37156 18676
rect 37212 19068 37268 19124
rect 36204 14700 36260 14756
rect 36316 13692 36372 13748
rect 36988 16940 37044 16996
rect 36540 12850 36596 12852
rect 36540 12798 36542 12850
rect 36542 12798 36594 12850
rect 36594 12798 36596 12850
rect 36540 12796 36596 12798
rect 36652 12738 36708 12740
rect 36652 12686 36654 12738
rect 36654 12686 36706 12738
rect 36706 12686 36708 12738
rect 36652 12684 36708 12686
rect 37660 19964 37716 20020
rect 37660 18620 37716 18676
rect 37996 18338 38052 18340
rect 37996 18286 37998 18338
rect 37998 18286 38050 18338
rect 38050 18286 38052 18338
rect 37996 18284 38052 18286
rect 37548 17612 37604 17668
rect 37884 17666 37940 17668
rect 37884 17614 37886 17666
rect 37886 17614 37938 17666
rect 37938 17614 37940 17666
rect 37884 17612 37940 17614
rect 37772 16882 37828 16884
rect 37772 16830 37774 16882
rect 37774 16830 37826 16882
rect 37826 16830 37828 16882
rect 37772 16828 37828 16830
rect 37884 16716 37940 16772
rect 37212 16156 37268 16212
rect 37660 16044 37716 16100
rect 37548 15260 37604 15316
rect 37324 13804 37380 13860
rect 37772 14252 37828 14308
rect 37548 13804 37604 13860
rect 37884 13858 37940 13860
rect 37884 13806 37886 13858
rect 37886 13806 37938 13858
rect 37938 13806 37940 13858
rect 37884 13804 37940 13806
rect 37100 12572 37156 12628
rect 37212 12684 37268 12740
rect 36204 11564 36260 11620
rect 36092 11004 36148 11060
rect 35756 10332 35812 10388
rect 35644 9996 35700 10052
rect 34748 9660 34804 9716
rect 34300 9324 34356 9380
rect 34188 8988 34244 9044
rect 34972 9714 35028 9716
rect 34972 9662 34974 9714
rect 34974 9662 35026 9714
rect 35026 9662 35028 9714
rect 34972 9660 35028 9662
rect 34860 9324 34916 9380
rect 34972 9266 35028 9268
rect 34972 9214 34974 9266
rect 34974 9214 35026 9266
rect 35026 9214 35028 9266
rect 34972 9212 35028 9214
rect 35308 9212 35364 9268
rect 34860 9154 34916 9156
rect 34860 9102 34862 9154
rect 34862 9102 34914 9154
rect 34914 9102 34916 9154
rect 34860 9100 34916 9102
rect 33404 7868 33460 7924
rect 36316 10498 36372 10500
rect 36316 10446 36318 10498
rect 36318 10446 36370 10498
rect 36370 10446 36372 10498
rect 36316 10444 36372 10446
rect 35756 9660 35812 9716
rect 36540 9714 36596 9716
rect 36540 9662 36542 9714
rect 36542 9662 36594 9714
rect 36594 9662 36596 9714
rect 36540 9660 36596 9662
rect 36428 9436 36484 9492
rect 36540 9266 36596 9268
rect 36540 9214 36542 9266
rect 36542 9214 36594 9266
rect 36594 9214 36596 9266
rect 36540 9212 36596 9214
rect 35756 8428 35812 8484
rect 36540 8818 36596 8820
rect 36540 8766 36542 8818
rect 36542 8766 36594 8818
rect 36594 8766 36596 8818
rect 36540 8764 36596 8766
rect 36764 8258 36820 8260
rect 36764 8206 36766 8258
rect 36766 8206 36818 8258
rect 36818 8206 36820 8258
rect 36764 8204 36820 8206
rect 37212 9548 37268 9604
rect 38668 20018 38724 20020
rect 38668 19966 38670 20018
rect 38670 19966 38722 20018
rect 38722 19966 38724 20018
rect 38668 19964 38724 19966
rect 39116 20412 39172 20468
rect 38668 19180 38724 19236
rect 39004 19234 39060 19236
rect 39004 19182 39006 19234
rect 39006 19182 39058 19234
rect 39058 19182 39060 19234
rect 39004 19180 39060 19182
rect 39116 18844 39172 18900
rect 38892 18674 38948 18676
rect 38892 18622 38894 18674
rect 38894 18622 38946 18674
rect 38946 18622 38948 18674
rect 38892 18620 38948 18622
rect 39228 18620 39284 18676
rect 38668 18450 38724 18452
rect 38668 18398 38670 18450
rect 38670 18398 38722 18450
rect 38722 18398 38724 18450
rect 38668 18396 38724 18398
rect 39004 18284 39060 18340
rect 38892 17612 38948 17668
rect 39452 21474 39508 21476
rect 39452 21422 39454 21474
rect 39454 21422 39506 21474
rect 39506 21422 39508 21474
rect 39452 21420 39508 21422
rect 39452 20300 39508 20356
rect 40124 21420 40180 21476
rect 39900 20524 39956 20580
rect 39852 20410 39908 20412
rect 39852 20358 39854 20410
rect 39854 20358 39906 20410
rect 39906 20358 39908 20410
rect 39852 20356 39908 20358
rect 39956 20410 40012 20412
rect 39956 20358 39958 20410
rect 39958 20358 40010 20410
rect 40010 20358 40012 20410
rect 39956 20356 40012 20358
rect 40060 20410 40116 20412
rect 40060 20358 40062 20410
rect 40062 20358 40114 20410
rect 40114 20358 40116 20410
rect 40060 20356 40116 20358
rect 39564 20130 39620 20132
rect 39564 20078 39566 20130
rect 39566 20078 39618 20130
rect 39618 20078 39620 20130
rect 39564 20076 39620 20078
rect 39676 19964 39732 20020
rect 39340 18060 39396 18116
rect 39900 19292 39956 19348
rect 39900 19010 39956 19012
rect 39900 18958 39902 19010
rect 39902 18958 39954 19010
rect 39954 18958 39956 19010
rect 39900 18956 39956 18958
rect 40348 20076 40404 20132
rect 41916 23154 41972 23156
rect 41916 23102 41918 23154
rect 41918 23102 41970 23154
rect 41970 23102 41972 23154
rect 41916 23100 41972 23102
rect 40908 22370 40964 22372
rect 40908 22318 40910 22370
rect 40910 22318 40962 22370
rect 40962 22318 40964 22370
rect 40908 22316 40964 22318
rect 41580 22652 41636 22708
rect 42476 22316 42532 22372
rect 40908 20188 40964 20244
rect 40684 20018 40740 20020
rect 40684 19966 40686 20018
rect 40686 19966 40738 20018
rect 40738 19966 40740 20018
rect 40684 19964 40740 19966
rect 40460 19180 40516 19236
rect 40348 19122 40404 19124
rect 40348 19070 40350 19122
rect 40350 19070 40402 19122
rect 40402 19070 40404 19122
rect 40348 19068 40404 19070
rect 39852 18842 39908 18844
rect 39852 18790 39854 18842
rect 39854 18790 39906 18842
rect 39906 18790 39908 18842
rect 39852 18788 39908 18790
rect 39956 18842 40012 18844
rect 39956 18790 39958 18842
rect 39958 18790 40010 18842
rect 40010 18790 40012 18842
rect 39956 18788 40012 18790
rect 40060 18842 40116 18844
rect 40060 18790 40062 18842
rect 40062 18790 40114 18842
rect 40114 18790 40116 18842
rect 40060 18788 40116 18790
rect 40236 18844 40292 18900
rect 40124 18620 40180 18676
rect 40572 18956 40628 19012
rect 39452 18396 39508 18452
rect 39340 17666 39396 17668
rect 39340 17614 39342 17666
rect 39342 17614 39394 17666
rect 39394 17614 39396 17666
rect 39340 17612 39396 17614
rect 39228 17388 39284 17444
rect 40460 18396 40516 18452
rect 39788 18226 39844 18228
rect 39788 18174 39790 18226
rect 39790 18174 39842 18226
rect 39842 18174 39844 18226
rect 39788 18172 39844 18174
rect 39676 17778 39732 17780
rect 39676 17726 39678 17778
rect 39678 17726 39730 17778
rect 39730 17726 39732 17778
rect 39676 17724 39732 17726
rect 39452 17052 39508 17108
rect 40348 17442 40404 17444
rect 40348 17390 40350 17442
rect 40350 17390 40402 17442
rect 40402 17390 40404 17442
rect 40348 17388 40404 17390
rect 40572 17442 40628 17444
rect 40572 17390 40574 17442
rect 40574 17390 40626 17442
rect 40626 17390 40628 17442
rect 40572 17388 40628 17390
rect 39852 17274 39908 17276
rect 39852 17222 39854 17274
rect 39854 17222 39906 17274
rect 39906 17222 39908 17274
rect 39852 17220 39908 17222
rect 39956 17274 40012 17276
rect 39956 17222 39958 17274
rect 39958 17222 40010 17274
rect 40010 17222 40012 17274
rect 39956 17220 40012 17222
rect 40060 17274 40116 17276
rect 40060 17222 40062 17274
rect 40062 17222 40114 17274
rect 40114 17222 40116 17274
rect 40236 17276 40292 17332
rect 40060 17220 40116 17222
rect 40796 18396 40852 18452
rect 41020 19292 41076 19348
rect 41580 19122 41636 19124
rect 41580 19070 41582 19122
rect 41582 19070 41634 19122
rect 41634 19070 41636 19122
rect 41580 19068 41636 19070
rect 41020 18732 41076 18788
rect 43036 22258 43092 22260
rect 43036 22206 43038 22258
rect 43038 22206 43090 22258
rect 43090 22206 43092 22258
rect 43036 22204 43092 22206
rect 41916 20914 41972 20916
rect 41916 20862 41918 20914
rect 41918 20862 41970 20914
rect 41970 20862 41972 20914
rect 41916 20860 41972 20862
rect 41804 20130 41860 20132
rect 41804 20078 41806 20130
rect 41806 20078 41858 20130
rect 41858 20078 41860 20130
rect 41804 20076 41860 20078
rect 42140 19964 42196 20020
rect 42700 19346 42756 19348
rect 42700 19294 42702 19346
rect 42702 19294 42754 19346
rect 42754 19294 42756 19346
rect 42700 19292 42756 19294
rect 41692 18732 41748 18788
rect 41916 18732 41972 18788
rect 41580 18396 41636 18452
rect 40908 17276 40964 17332
rect 40908 17106 40964 17108
rect 40908 17054 40910 17106
rect 40910 17054 40962 17106
rect 40962 17054 40964 17106
rect 40908 17052 40964 17054
rect 38444 16098 38500 16100
rect 38444 16046 38446 16098
rect 38446 16046 38498 16098
rect 38498 16046 38500 16098
rect 38444 16044 38500 16046
rect 38668 15820 38724 15876
rect 39004 15820 39060 15876
rect 39116 16044 39172 16100
rect 38892 15708 38948 15764
rect 39564 15932 39620 15988
rect 40572 16604 40628 16660
rect 40460 16380 40516 16436
rect 40124 16156 40180 16212
rect 39900 16098 39956 16100
rect 39900 16046 39902 16098
rect 39902 16046 39954 16098
rect 39954 16046 39956 16098
rect 39900 16044 39956 16046
rect 40236 15874 40292 15876
rect 40236 15822 40238 15874
rect 40238 15822 40290 15874
rect 40290 15822 40292 15874
rect 40236 15820 40292 15822
rect 39852 15706 39908 15708
rect 39852 15654 39854 15706
rect 39854 15654 39906 15706
rect 39906 15654 39908 15706
rect 39852 15652 39908 15654
rect 39956 15706 40012 15708
rect 39956 15654 39958 15706
rect 39958 15654 40010 15706
rect 40010 15654 40012 15706
rect 39956 15652 40012 15654
rect 40060 15706 40116 15708
rect 40060 15654 40062 15706
rect 40062 15654 40114 15706
rect 40114 15654 40116 15706
rect 40060 15652 40116 15654
rect 38892 15148 38948 15204
rect 38444 13804 38500 13860
rect 39788 14924 39844 14980
rect 40236 14588 40292 14644
rect 39116 14476 39172 14532
rect 39900 14418 39956 14420
rect 39900 14366 39902 14418
rect 39902 14366 39954 14418
rect 39954 14366 39956 14418
rect 39900 14364 39956 14366
rect 40348 14418 40404 14420
rect 40348 14366 40350 14418
rect 40350 14366 40402 14418
rect 40402 14366 40404 14418
rect 40348 14364 40404 14366
rect 39788 14306 39844 14308
rect 39788 14254 39790 14306
rect 39790 14254 39842 14306
rect 39842 14254 39844 14306
rect 39788 14252 39844 14254
rect 39852 14138 39908 14140
rect 39852 14086 39854 14138
rect 39854 14086 39906 14138
rect 39906 14086 39908 14138
rect 39852 14084 39908 14086
rect 39956 14138 40012 14140
rect 39956 14086 39958 14138
rect 39958 14086 40010 14138
rect 40010 14086 40012 14138
rect 39956 14084 40012 14086
rect 40060 14138 40116 14140
rect 40060 14086 40062 14138
rect 40062 14086 40114 14138
rect 40114 14086 40116 14138
rect 40060 14084 40116 14086
rect 39676 13746 39732 13748
rect 39676 13694 39678 13746
rect 39678 13694 39730 13746
rect 39730 13694 39732 13746
rect 39676 13692 39732 13694
rect 39900 13580 39956 13636
rect 37884 12796 37940 12852
rect 37772 12684 37828 12740
rect 38556 11116 38612 11172
rect 39116 11170 39172 11172
rect 39116 11118 39118 11170
rect 39118 11118 39170 11170
rect 39170 11118 39172 11170
rect 39116 11116 39172 11118
rect 37436 9602 37492 9604
rect 37436 9550 37438 9602
rect 37438 9550 37490 9602
rect 37490 9550 37492 9602
rect 37436 9548 37492 9550
rect 38668 10498 38724 10500
rect 38668 10446 38670 10498
rect 38670 10446 38722 10498
rect 38722 10446 38724 10498
rect 38668 10444 38724 10446
rect 39852 12570 39908 12572
rect 39852 12518 39854 12570
rect 39854 12518 39906 12570
rect 39906 12518 39908 12570
rect 39852 12516 39908 12518
rect 39956 12570 40012 12572
rect 39956 12518 39958 12570
rect 39958 12518 40010 12570
rect 40010 12518 40012 12570
rect 39956 12516 40012 12518
rect 40060 12570 40116 12572
rect 40060 12518 40062 12570
rect 40062 12518 40114 12570
rect 40114 12518 40116 12570
rect 40060 12516 40116 12518
rect 40348 13692 40404 13748
rect 40348 12460 40404 12516
rect 40124 12012 40180 12068
rect 39228 10444 39284 10500
rect 39116 10220 39172 10276
rect 38220 9548 38276 9604
rect 37884 9436 37940 9492
rect 37212 9212 37268 9268
rect 36876 8092 36932 8148
rect 36428 7756 36484 7812
rect 35196 7308 35252 7364
rect 36316 7362 36372 7364
rect 36316 7310 36318 7362
rect 36318 7310 36370 7362
rect 36370 7310 36372 7362
rect 36316 7308 36372 7310
rect 34972 6690 35028 6692
rect 34972 6638 34974 6690
rect 34974 6638 35026 6690
rect 35026 6638 35028 6690
rect 34972 6636 35028 6638
rect 34860 6578 34916 6580
rect 34860 6526 34862 6578
rect 34862 6526 34914 6578
rect 34914 6526 34916 6578
rect 34860 6524 34916 6526
rect 34188 6466 34244 6468
rect 34188 6414 34190 6466
rect 34190 6414 34242 6466
rect 34242 6414 34244 6466
rect 34188 6412 34244 6414
rect 32732 4338 32788 4340
rect 32732 4286 32734 4338
rect 32734 4286 32786 4338
rect 32786 4286 32788 4338
rect 32732 4284 32788 4286
rect 35084 6466 35140 6468
rect 35084 6414 35086 6466
rect 35086 6414 35138 6466
rect 35138 6414 35140 6466
rect 35084 6412 35140 6414
rect 35084 5964 35140 6020
rect 34188 5292 34244 5348
rect 34076 5234 34132 5236
rect 34076 5182 34078 5234
rect 34078 5182 34130 5234
rect 34130 5182 34132 5234
rect 34076 5180 34132 5182
rect 34412 5068 34468 5124
rect 34860 5068 34916 5124
rect 37212 7196 37268 7252
rect 37324 8428 37380 8484
rect 36428 6578 36484 6580
rect 36428 6526 36430 6578
rect 36430 6526 36482 6578
rect 36482 6526 36484 6578
rect 36428 6524 36484 6526
rect 35980 6412 36036 6468
rect 35196 5292 35252 5348
rect 35532 5740 35588 5796
rect 35980 5628 36036 5684
rect 36988 6076 37044 6132
rect 35532 5180 35588 5236
rect 33852 4396 33908 4452
rect 33628 4338 33684 4340
rect 33628 4286 33630 4338
rect 33630 4286 33682 4338
rect 33682 4286 33684 4338
rect 33628 4284 33684 4286
rect 33516 3724 33572 3780
rect 32172 3612 32228 3668
rect 32508 3554 32564 3556
rect 32508 3502 32510 3554
rect 32510 3502 32562 3554
rect 32562 3502 32564 3554
rect 32508 3500 32564 3502
rect 31612 3442 31668 3444
rect 31612 3390 31614 3442
rect 31614 3390 31666 3442
rect 31666 3390 31668 3442
rect 31612 3388 31668 3390
rect 32396 3388 32452 3444
rect 33180 3442 33236 3444
rect 33180 3390 33182 3442
rect 33182 3390 33234 3442
rect 33234 3390 33236 3442
rect 33180 3388 33236 3390
rect 34076 4508 34132 4564
rect 35644 4450 35700 4452
rect 35644 4398 35646 4450
rect 35646 4398 35698 4450
rect 35698 4398 35700 4450
rect 35644 4396 35700 4398
rect 34412 4226 34468 4228
rect 34412 4174 34414 4226
rect 34414 4174 34466 4226
rect 34466 4174 34468 4226
rect 34412 4172 34468 4174
rect 34188 3778 34244 3780
rect 34188 3726 34190 3778
rect 34190 3726 34242 3778
rect 34242 3726 34244 3778
rect 34188 3724 34244 3726
rect 34860 3554 34916 3556
rect 34860 3502 34862 3554
rect 34862 3502 34914 3554
rect 34914 3502 34916 3554
rect 34860 3500 34916 3502
rect 28812 1260 28868 1316
rect 35980 3554 36036 3556
rect 35980 3502 35982 3554
rect 35982 3502 36034 3554
rect 36034 3502 36036 3554
rect 35980 3500 36036 3502
rect 35084 1596 35140 1652
rect 35308 2716 35364 2772
rect 36316 5740 36372 5796
rect 36540 6018 36596 6020
rect 36540 5966 36542 6018
rect 36542 5966 36594 6018
rect 36594 5966 36596 6018
rect 36540 5964 36596 5966
rect 36204 5628 36260 5684
rect 36876 5794 36932 5796
rect 36876 5742 36878 5794
rect 36878 5742 36930 5794
rect 36930 5742 36932 5794
rect 36876 5740 36932 5742
rect 36764 5010 36820 5012
rect 36764 4958 36766 5010
rect 36766 4958 36818 5010
rect 36818 4958 36820 5010
rect 36764 4956 36820 4958
rect 37548 8876 37604 8932
rect 37884 8428 37940 8484
rect 39788 11170 39844 11172
rect 39788 11118 39790 11170
rect 39790 11118 39842 11170
rect 39842 11118 39844 11170
rect 39788 11116 39844 11118
rect 39852 11002 39908 11004
rect 39852 10950 39854 11002
rect 39854 10950 39906 11002
rect 39906 10950 39908 11002
rect 39852 10948 39908 10950
rect 39956 11002 40012 11004
rect 39956 10950 39958 11002
rect 39958 10950 40010 11002
rect 40010 10950 40012 11002
rect 39956 10948 40012 10950
rect 40060 11002 40116 11004
rect 40060 10950 40062 11002
rect 40062 10950 40114 11002
rect 40114 10950 40116 11002
rect 40060 10948 40116 10950
rect 40124 10610 40180 10612
rect 40124 10558 40126 10610
rect 40126 10558 40178 10610
rect 40178 10558 40180 10610
rect 40124 10556 40180 10558
rect 40012 10498 40068 10500
rect 40012 10446 40014 10498
rect 40014 10446 40066 10498
rect 40066 10446 40068 10498
rect 40012 10444 40068 10446
rect 39900 10108 39956 10164
rect 38668 9602 38724 9604
rect 38668 9550 38670 9602
rect 38670 9550 38722 9602
rect 38722 9550 38724 9602
rect 38668 9548 38724 9550
rect 40012 9602 40068 9604
rect 40012 9550 40014 9602
rect 40014 9550 40066 9602
rect 40066 9550 40068 9602
rect 40012 9548 40068 9550
rect 37772 8258 37828 8260
rect 37772 8206 37774 8258
rect 37774 8206 37826 8258
rect 37826 8206 37828 8258
rect 37772 8204 37828 8206
rect 38220 8146 38276 8148
rect 38220 8094 38222 8146
rect 38222 8094 38274 8146
rect 38274 8094 38276 8146
rect 38220 8092 38276 8094
rect 37772 7756 37828 7812
rect 37548 7308 37604 7364
rect 37660 7196 37716 7252
rect 37436 6466 37492 6468
rect 37436 6414 37438 6466
rect 37438 6414 37490 6466
rect 37490 6414 37492 6466
rect 37436 6412 37492 6414
rect 37324 5628 37380 5684
rect 36988 4396 37044 4452
rect 36204 4226 36260 4228
rect 36204 4174 36206 4226
rect 36206 4174 36258 4226
rect 36258 4174 36260 4226
rect 36204 4172 36260 4174
rect 37100 4226 37156 4228
rect 37100 4174 37102 4226
rect 37102 4174 37154 4226
rect 37154 4174 37156 4226
rect 37100 4172 37156 4174
rect 36764 3500 36820 3556
rect 36428 3442 36484 3444
rect 36428 3390 36430 3442
rect 36430 3390 36482 3442
rect 36482 3390 36484 3442
rect 36428 3388 36484 3390
rect 36092 2156 36148 2212
rect 35308 1372 35364 1428
rect 37100 3554 37156 3556
rect 37100 3502 37102 3554
rect 37102 3502 37154 3554
rect 37154 3502 37156 3554
rect 37100 3500 37156 3502
rect 37436 2716 37492 2772
rect 37436 2268 37492 2324
rect 37660 6412 37716 6468
rect 39852 9434 39908 9436
rect 39852 9382 39854 9434
rect 39854 9382 39906 9434
rect 39906 9382 39908 9434
rect 39852 9380 39908 9382
rect 39956 9434 40012 9436
rect 39956 9382 39958 9434
rect 39958 9382 40010 9434
rect 40010 9382 40012 9434
rect 39956 9380 40012 9382
rect 40060 9434 40116 9436
rect 40060 9382 40062 9434
rect 40062 9382 40114 9434
rect 40114 9382 40116 9434
rect 40060 9380 40116 9382
rect 39564 9266 39620 9268
rect 39564 9214 39566 9266
rect 39566 9214 39618 9266
rect 39618 9214 39620 9266
rect 39564 9212 39620 9214
rect 38444 7362 38500 7364
rect 38444 7310 38446 7362
rect 38446 7310 38498 7362
rect 38498 7310 38500 7362
rect 38444 7308 38500 7310
rect 38332 7196 38388 7252
rect 37996 5964 38052 6020
rect 38892 6972 38948 7028
rect 38668 5906 38724 5908
rect 38668 5854 38670 5906
rect 38670 5854 38722 5906
rect 38722 5854 38724 5906
rect 38668 5852 38724 5854
rect 37660 5292 37716 5348
rect 38108 5122 38164 5124
rect 38108 5070 38110 5122
rect 38110 5070 38162 5122
rect 38162 5070 38164 5122
rect 38108 5068 38164 5070
rect 37772 4508 37828 4564
rect 37884 4844 37940 4900
rect 40012 9154 40068 9156
rect 40012 9102 40014 9154
rect 40014 9102 40066 9154
rect 40066 9102 40068 9154
rect 40012 9100 40068 9102
rect 39852 7866 39908 7868
rect 39852 7814 39854 7866
rect 39854 7814 39906 7866
rect 39906 7814 39908 7866
rect 39852 7812 39908 7814
rect 39956 7866 40012 7868
rect 39956 7814 39958 7866
rect 39958 7814 40010 7866
rect 40010 7814 40012 7866
rect 39956 7812 40012 7814
rect 40060 7866 40116 7868
rect 40060 7814 40062 7866
rect 40062 7814 40114 7866
rect 40114 7814 40116 7866
rect 40060 7812 40116 7814
rect 41804 18284 41860 18340
rect 41692 17778 41748 17780
rect 41692 17726 41694 17778
rect 41694 17726 41746 17778
rect 41746 17726 41748 17778
rect 41692 17724 41748 17726
rect 41804 17052 41860 17108
rect 41804 16828 41860 16884
rect 41692 15820 41748 15876
rect 40572 15148 40628 15204
rect 42588 19010 42644 19012
rect 42588 18958 42590 19010
rect 42590 18958 42642 19010
rect 42642 18958 42644 19010
rect 42588 18956 42644 18958
rect 42364 18508 42420 18564
rect 42252 18450 42308 18452
rect 42252 18398 42254 18450
rect 42254 18398 42306 18450
rect 42306 18398 42308 18450
rect 42252 18396 42308 18398
rect 42588 18338 42644 18340
rect 42588 18286 42590 18338
rect 42590 18286 42642 18338
rect 42642 18286 42644 18338
rect 42588 18284 42644 18286
rect 42588 18060 42644 18116
rect 42028 17388 42084 17444
rect 42028 16940 42084 16996
rect 42476 16994 42532 16996
rect 42476 16942 42478 16994
rect 42478 16942 42530 16994
rect 42530 16942 42532 16994
rect 42476 16940 42532 16942
rect 41916 16268 41972 16324
rect 42028 16770 42084 16772
rect 42028 16718 42030 16770
rect 42030 16718 42082 16770
rect 42082 16718 42084 16770
rect 42028 16716 42084 16718
rect 42028 16492 42084 16548
rect 42476 15314 42532 15316
rect 42476 15262 42478 15314
rect 42478 15262 42530 15314
rect 42530 15262 42532 15314
rect 42476 15260 42532 15262
rect 41916 14700 41972 14756
rect 42028 15036 42084 15092
rect 40684 14530 40740 14532
rect 40684 14478 40686 14530
rect 40686 14478 40738 14530
rect 40738 14478 40740 14530
rect 40684 14476 40740 14478
rect 41580 14306 41636 14308
rect 41580 14254 41582 14306
rect 41582 14254 41634 14306
rect 41634 14254 41636 14306
rect 41580 14252 41636 14254
rect 40684 14140 40740 14196
rect 40572 13746 40628 13748
rect 40572 13694 40574 13746
rect 40574 13694 40626 13746
rect 40626 13694 40628 13746
rect 40572 13692 40628 13694
rect 40796 13580 40852 13636
rect 41580 13468 41636 13524
rect 42476 14588 42532 14644
rect 42252 14252 42308 14308
rect 42700 15874 42756 15876
rect 42700 15822 42702 15874
rect 42702 15822 42754 15874
rect 42754 15822 42756 15874
rect 42700 15820 42756 15822
rect 43036 15314 43092 15316
rect 43036 15262 43038 15314
rect 43038 15262 43090 15314
rect 43090 15262 43092 15314
rect 43036 15260 43092 15262
rect 43932 26460 43988 26516
rect 43372 26348 43428 26404
rect 43820 26402 43876 26404
rect 43820 26350 43822 26402
rect 43822 26350 43874 26402
rect 43874 26350 43876 26402
rect 43820 26348 43876 26350
rect 45052 27020 45108 27076
rect 44044 26236 44100 26292
rect 44380 26348 44436 26404
rect 44492 26290 44548 26292
rect 44492 26238 44494 26290
rect 44494 26238 44546 26290
rect 44546 26238 44548 26290
rect 44492 26236 44548 26238
rect 44380 25452 44436 25508
rect 46284 27970 46340 27972
rect 46284 27918 46286 27970
rect 46286 27918 46338 27970
rect 46338 27918 46340 27970
rect 46284 27916 46340 27918
rect 45948 27580 46004 27636
rect 46620 27858 46676 27860
rect 46620 27806 46622 27858
rect 46622 27806 46674 27858
rect 46674 27806 46676 27858
rect 46620 27804 46676 27806
rect 46508 27746 46564 27748
rect 46508 27694 46510 27746
rect 46510 27694 46562 27746
rect 46562 27694 46564 27746
rect 46508 27692 46564 27694
rect 46844 27580 46900 27636
rect 46060 27074 46116 27076
rect 46060 27022 46062 27074
rect 46062 27022 46114 27074
rect 46114 27022 46116 27074
rect 46060 27020 46116 27022
rect 46284 27020 46340 27076
rect 45500 26514 45556 26516
rect 45500 26462 45502 26514
rect 45502 26462 45554 26514
rect 45554 26462 45556 26514
rect 45500 26460 45556 26462
rect 44604 25340 44660 25396
rect 43484 24834 43540 24836
rect 43484 24782 43486 24834
rect 43486 24782 43538 24834
rect 43538 24782 43540 24834
rect 43484 24780 43540 24782
rect 44044 24834 44100 24836
rect 44044 24782 44046 24834
rect 44046 24782 44098 24834
rect 44098 24782 44100 24834
rect 44044 24780 44100 24782
rect 44268 24556 44324 24612
rect 44940 25452 44996 25508
rect 45500 25394 45556 25396
rect 45500 25342 45502 25394
rect 45502 25342 45554 25394
rect 45554 25342 45556 25394
rect 45500 25340 45556 25342
rect 45612 25282 45668 25284
rect 45612 25230 45614 25282
rect 45614 25230 45666 25282
rect 45666 25230 45668 25282
rect 45612 25228 45668 25230
rect 48412 32956 48468 33012
rect 48076 32786 48132 32788
rect 48076 32734 48078 32786
rect 48078 32734 48130 32786
rect 48130 32734 48132 32786
rect 48076 32732 48132 32734
rect 47628 31778 47684 31780
rect 47628 31726 47630 31778
rect 47630 31726 47682 31778
rect 47682 31726 47684 31778
rect 47628 31724 47684 31726
rect 47516 31554 47572 31556
rect 47516 31502 47518 31554
rect 47518 31502 47570 31554
rect 47570 31502 47572 31554
rect 47516 31500 47572 31502
rect 47852 31500 47908 31556
rect 48076 31554 48132 31556
rect 48076 31502 48078 31554
rect 48078 31502 48130 31554
rect 48130 31502 48132 31554
rect 48076 31500 48132 31502
rect 48748 30268 48804 30324
rect 47740 30098 47796 30100
rect 47740 30046 47742 30098
rect 47742 30046 47794 30098
rect 47794 30046 47796 30098
rect 47740 30044 47796 30046
rect 48188 28700 48244 28756
rect 48076 28588 48132 28644
rect 48748 29202 48804 29204
rect 48748 29150 48750 29202
rect 48750 29150 48802 29202
rect 48802 29150 48804 29202
rect 48748 29148 48804 29150
rect 48300 28642 48356 28644
rect 48300 28590 48302 28642
rect 48302 28590 48354 28642
rect 48354 28590 48356 28642
rect 48300 28588 48356 28590
rect 48412 28700 48468 28756
rect 48636 28642 48692 28644
rect 48636 28590 48638 28642
rect 48638 28590 48690 28642
rect 48690 28590 48692 28642
rect 48636 28588 48692 28590
rect 48748 27692 48804 27748
rect 48524 27074 48580 27076
rect 48524 27022 48526 27074
rect 48526 27022 48578 27074
rect 48578 27022 48580 27074
rect 48524 27020 48580 27022
rect 47404 26796 47460 26852
rect 49512 33738 49568 33740
rect 49512 33686 49514 33738
rect 49514 33686 49566 33738
rect 49566 33686 49568 33738
rect 49512 33684 49568 33686
rect 49616 33738 49672 33740
rect 49616 33686 49618 33738
rect 49618 33686 49670 33738
rect 49670 33686 49672 33738
rect 49616 33684 49672 33686
rect 49720 33738 49776 33740
rect 49720 33686 49722 33738
rect 49722 33686 49774 33738
rect 49774 33686 49776 33738
rect 49720 33684 49776 33686
rect 49644 33346 49700 33348
rect 49644 33294 49646 33346
rect 49646 33294 49698 33346
rect 49698 33294 49700 33346
rect 49644 33292 49700 33294
rect 49980 34636 50036 34692
rect 50316 34690 50372 34692
rect 50316 34638 50318 34690
rect 50318 34638 50370 34690
rect 50370 34638 50372 34690
rect 50316 34636 50372 34638
rect 50876 34914 50932 34916
rect 50876 34862 50878 34914
rect 50878 34862 50930 34914
rect 50930 34862 50932 34914
rect 50876 34860 50932 34862
rect 51212 34412 51268 34468
rect 52780 35756 52836 35812
rect 53116 35868 53172 35924
rect 53116 35644 53172 35700
rect 58380 36540 58436 36596
rect 58828 36594 58884 36596
rect 58828 36542 58830 36594
rect 58830 36542 58882 36594
rect 58882 36542 58884 36594
rect 58828 36540 58884 36542
rect 63196 37548 63252 37604
rect 52556 35586 52612 35588
rect 52556 35534 52558 35586
rect 52558 35534 52610 35586
rect 52610 35534 52612 35586
rect 52556 35532 52612 35534
rect 51996 34636 52052 34692
rect 50092 33292 50148 33348
rect 49532 32562 49588 32564
rect 49532 32510 49534 32562
rect 49534 32510 49586 32562
rect 49586 32510 49588 32562
rect 49532 32508 49588 32510
rect 49512 32170 49568 32172
rect 49512 32118 49514 32170
rect 49514 32118 49566 32170
rect 49566 32118 49568 32170
rect 49512 32116 49568 32118
rect 49616 32170 49672 32172
rect 49616 32118 49618 32170
rect 49618 32118 49670 32170
rect 49670 32118 49672 32170
rect 49616 32116 49672 32118
rect 49720 32170 49776 32172
rect 49720 32118 49722 32170
rect 49722 32118 49774 32170
rect 49774 32118 49776 32170
rect 49720 32116 49776 32118
rect 49308 31724 49364 31780
rect 50428 33346 50484 33348
rect 50428 33294 50430 33346
rect 50430 33294 50482 33346
rect 50482 33294 50484 33346
rect 50428 33292 50484 33294
rect 51884 34130 51940 34132
rect 51884 34078 51886 34130
rect 51886 34078 51938 34130
rect 51938 34078 51940 34130
rect 51884 34076 51940 34078
rect 50988 33346 51044 33348
rect 50988 33294 50990 33346
rect 50990 33294 51042 33346
rect 51042 33294 51044 33346
rect 50988 33292 51044 33294
rect 50652 33068 50708 33124
rect 51548 33180 51604 33236
rect 51772 33234 51828 33236
rect 51772 33182 51774 33234
rect 51774 33182 51826 33234
rect 51826 33182 51828 33234
rect 51772 33180 51828 33182
rect 50988 33068 51044 33124
rect 50764 32732 50820 32788
rect 51660 33122 51716 33124
rect 51660 33070 51662 33122
rect 51662 33070 51714 33122
rect 51714 33070 51716 33122
rect 51660 33068 51716 33070
rect 52780 34130 52836 34132
rect 52780 34078 52782 34130
rect 52782 34078 52834 34130
rect 52834 34078 52836 34130
rect 52780 34076 52836 34078
rect 52556 33292 52612 33348
rect 53116 33292 53172 33348
rect 52332 33180 52388 33236
rect 52220 32674 52276 32676
rect 52220 32622 52222 32674
rect 52222 32622 52274 32674
rect 52274 32622 52276 32674
rect 52220 32620 52276 32622
rect 52332 32284 52388 32340
rect 52780 33122 52836 33124
rect 52780 33070 52782 33122
rect 52782 33070 52834 33122
rect 52834 33070 52836 33122
rect 52780 33068 52836 33070
rect 49980 31778 50036 31780
rect 49980 31726 49982 31778
rect 49982 31726 50034 31778
rect 50034 31726 50036 31778
rect 49980 31724 50036 31726
rect 49756 31052 49812 31108
rect 51100 31666 51156 31668
rect 51100 31614 51102 31666
rect 51102 31614 51154 31666
rect 51154 31614 51156 31666
rect 51100 31612 51156 31614
rect 50428 31106 50484 31108
rect 50428 31054 50430 31106
rect 50430 31054 50482 31106
rect 50482 31054 50484 31106
rect 50428 31052 50484 31054
rect 49512 30602 49568 30604
rect 49512 30550 49514 30602
rect 49514 30550 49566 30602
rect 49566 30550 49568 30602
rect 49512 30548 49568 30550
rect 49616 30602 49672 30604
rect 49616 30550 49618 30602
rect 49618 30550 49670 30602
rect 49670 30550 49672 30602
rect 49616 30548 49672 30550
rect 49720 30602 49776 30604
rect 49720 30550 49722 30602
rect 49722 30550 49774 30602
rect 49774 30550 49776 30602
rect 49720 30548 49776 30550
rect 49756 30322 49812 30324
rect 49756 30270 49758 30322
rect 49758 30270 49810 30322
rect 49810 30270 49812 30322
rect 49756 30268 49812 30270
rect 51212 31554 51268 31556
rect 51212 31502 51214 31554
rect 51214 31502 51266 31554
rect 51266 31502 51268 31554
rect 51212 31500 51268 31502
rect 50988 30604 51044 30660
rect 50428 29596 50484 29652
rect 49644 29426 49700 29428
rect 49644 29374 49646 29426
rect 49646 29374 49698 29426
rect 49698 29374 49700 29426
rect 49644 29372 49700 29374
rect 49868 29148 49924 29204
rect 49512 29034 49568 29036
rect 49512 28982 49514 29034
rect 49514 28982 49566 29034
rect 49566 28982 49568 29034
rect 49512 28980 49568 28982
rect 49616 29034 49672 29036
rect 49616 28982 49618 29034
rect 49618 28982 49670 29034
rect 49670 28982 49672 29034
rect 49616 28980 49672 28982
rect 49720 29034 49776 29036
rect 49720 28982 49722 29034
rect 49722 28982 49774 29034
rect 49774 28982 49776 29034
rect 49720 28980 49776 28982
rect 49868 27692 49924 27748
rect 51100 29650 51156 29652
rect 51100 29598 51102 29650
rect 51102 29598 51154 29650
rect 51154 29598 51156 29650
rect 51100 29596 51156 29598
rect 50540 28700 50596 28756
rect 50204 27692 50260 27748
rect 49756 27580 49812 27636
rect 49512 27466 49568 27468
rect 49512 27414 49514 27466
rect 49514 27414 49566 27466
rect 49566 27414 49568 27466
rect 49512 27412 49568 27414
rect 49616 27466 49672 27468
rect 49616 27414 49618 27466
rect 49618 27414 49670 27466
rect 49670 27414 49672 27466
rect 49616 27412 49672 27414
rect 49720 27466 49776 27468
rect 49720 27414 49722 27466
rect 49722 27414 49774 27466
rect 49774 27414 49776 27466
rect 49720 27412 49776 27414
rect 49308 26908 49364 26964
rect 49196 26684 49252 26740
rect 48188 26348 48244 26404
rect 49756 26402 49812 26404
rect 49756 26350 49758 26402
rect 49758 26350 49810 26402
rect 49810 26350 49812 26402
rect 49756 26348 49812 26350
rect 49196 26236 49252 26292
rect 50428 26236 50484 26292
rect 50764 26290 50820 26292
rect 50764 26238 50766 26290
rect 50766 26238 50818 26290
rect 50818 26238 50820 26290
rect 50764 26236 50820 26238
rect 47404 25676 47460 25732
rect 45388 24610 45444 24612
rect 45388 24558 45390 24610
rect 45390 24558 45442 24610
rect 45442 24558 45444 24610
rect 45388 24556 45444 24558
rect 44268 23100 44324 23156
rect 46956 23772 47012 23828
rect 46172 23266 46228 23268
rect 46172 23214 46174 23266
rect 46174 23214 46226 23266
rect 46226 23214 46228 23266
rect 46172 23212 46228 23214
rect 44492 22988 44548 23044
rect 43820 22204 43876 22260
rect 45500 23154 45556 23156
rect 45500 23102 45502 23154
rect 45502 23102 45554 23154
rect 45554 23102 45556 23154
rect 45500 23100 45556 23102
rect 45612 23042 45668 23044
rect 45612 22990 45614 23042
rect 45614 22990 45666 23042
rect 45666 22990 45668 23042
rect 45612 22988 45668 22990
rect 47516 23772 47572 23828
rect 47180 23266 47236 23268
rect 47180 23214 47182 23266
rect 47182 23214 47234 23266
rect 47234 23214 47236 23266
rect 47180 23212 47236 23214
rect 48412 26066 48468 26068
rect 48412 26014 48414 26066
rect 48414 26014 48466 26066
rect 48466 26014 48468 26066
rect 48412 26012 48468 26014
rect 49532 26066 49588 26068
rect 49532 26014 49534 26066
rect 49534 26014 49586 26066
rect 49586 26014 49588 26066
rect 49532 26012 49588 26014
rect 49512 25898 49568 25900
rect 49512 25846 49514 25898
rect 49514 25846 49566 25898
rect 49566 25846 49568 25898
rect 49512 25844 49568 25846
rect 49616 25898 49672 25900
rect 49616 25846 49618 25898
rect 49618 25846 49670 25898
rect 49670 25846 49672 25898
rect 49616 25844 49672 25846
rect 49720 25898 49776 25900
rect 49720 25846 49722 25898
rect 49722 25846 49774 25898
rect 49774 25846 49776 25898
rect 49720 25844 49776 25846
rect 49308 24892 49364 24948
rect 48748 24108 48804 24164
rect 47740 23212 47796 23268
rect 45724 22370 45780 22372
rect 45724 22318 45726 22370
rect 45726 22318 45778 22370
rect 45778 22318 45780 22370
rect 45724 22316 45780 22318
rect 44828 22204 44884 22260
rect 45388 22092 45444 22148
rect 45948 22092 46004 22148
rect 44268 21698 44324 21700
rect 44268 21646 44270 21698
rect 44270 21646 44322 21698
rect 44322 21646 44324 21698
rect 44268 21644 44324 21646
rect 43372 19906 43428 19908
rect 43372 19854 43374 19906
rect 43374 19854 43426 19906
rect 43426 19854 43428 19906
rect 43372 19852 43428 19854
rect 43596 19346 43652 19348
rect 43596 19294 43598 19346
rect 43598 19294 43650 19346
rect 43650 19294 43652 19346
rect 43596 19292 43652 19294
rect 46508 21532 46564 21588
rect 44604 20690 44660 20692
rect 44604 20638 44606 20690
rect 44606 20638 44658 20690
rect 44658 20638 44660 20690
rect 44604 20636 44660 20638
rect 44380 20578 44436 20580
rect 44380 20526 44382 20578
rect 44382 20526 44434 20578
rect 44434 20526 44436 20578
rect 44380 20524 44436 20526
rect 45388 20524 45444 20580
rect 44716 20076 44772 20132
rect 44156 20018 44212 20020
rect 44156 19966 44158 20018
rect 44158 19966 44210 20018
rect 44210 19966 44212 20018
rect 44156 19964 44212 19966
rect 43932 19906 43988 19908
rect 43932 19854 43934 19906
rect 43934 19854 43986 19906
rect 43986 19854 43988 19906
rect 43932 19852 43988 19854
rect 43372 18620 43428 18676
rect 43596 18508 43652 18564
rect 43484 18338 43540 18340
rect 43484 18286 43486 18338
rect 43486 18286 43538 18338
rect 43538 18286 43540 18338
rect 43484 18284 43540 18286
rect 43708 18396 43764 18452
rect 43596 17836 43652 17892
rect 43820 16828 43876 16884
rect 47292 22930 47348 22932
rect 47292 22878 47294 22930
rect 47294 22878 47346 22930
rect 47346 22878 47348 22930
rect 47292 22876 47348 22878
rect 47404 22540 47460 22596
rect 47292 22146 47348 22148
rect 47292 22094 47294 22146
rect 47294 22094 47346 22146
rect 47346 22094 47348 22146
rect 47292 22092 47348 22094
rect 46956 21532 47012 21588
rect 46172 20018 46228 20020
rect 46172 19966 46174 20018
rect 46174 19966 46226 20018
rect 46226 19966 46228 20018
rect 46172 19964 46228 19966
rect 45500 19906 45556 19908
rect 45500 19854 45502 19906
rect 45502 19854 45554 19906
rect 45554 19854 45556 19906
rect 45500 19852 45556 19854
rect 45276 19516 45332 19572
rect 44492 18060 44548 18116
rect 44940 18396 44996 18452
rect 43932 16380 43988 16436
rect 43372 15426 43428 15428
rect 43372 15374 43374 15426
rect 43374 15374 43426 15426
rect 43426 15374 43428 15426
rect 43372 15372 43428 15374
rect 43596 14812 43652 14868
rect 43372 14588 43428 14644
rect 43260 14028 43316 14084
rect 44044 15260 44100 15316
rect 44156 15426 44212 15428
rect 44156 15374 44158 15426
rect 44158 15374 44210 15426
rect 44210 15374 44212 15426
rect 44156 15372 44212 15374
rect 44268 16716 44324 16772
rect 44604 15314 44660 15316
rect 44604 15262 44606 15314
rect 44606 15262 44658 15314
rect 44658 15262 44660 15314
rect 44604 15260 44660 15262
rect 45276 17052 45332 17108
rect 46508 20130 46564 20132
rect 46508 20078 46510 20130
rect 46510 20078 46562 20130
rect 46562 20078 46564 20130
rect 46508 20076 46564 20078
rect 46284 19740 46340 19796
rect 46844 19740 46900 19796
rect 47068 19628 47124 19684
rect 45836 18674 45892 18676
rect 45836 18622 45838 18674
rect 45838 18622 45890 18674
rect 45890 18622 45892 18674
rect 45836 18620 45892 18622
rect 45500 18450 45556 18452
rect 45500 18398 45502 18450
rect 45502 18398 45554 18450
rect 45554 18398 45556 18450
rect 45500 18396 45556 18398
rect 45836 18396 45892 18452
rect 45724 17724 45780 17780
rect 47068 18396 47124 18452
rect 46956 17612 47012 17668
rect 47180 17388 47236 17444
rect 45388 16716 45444 16772
rect 45612 16492 45668 16548
rect 46284 16492 46340 16548
rect 46396 16940 46452 16996
rect 44716 14924 44772 14980
rect 46508 15708 46564 15764
rect 46060 14476 46116 14532
rect 45948 14140 46004 14196
rect 45388 13858 45444 13860
rect 45388 13806 45390 13858
rect 45390 13806 45442 13858
rect 45442 13806 45444 13858
rect 45388 13804 45444 13806
rect 46284 14140 46340 14196
rect 47068 16770 47124 16772
rect 47068 16718 47070 16770
rect 47070 16718 47122 16770
rect 47122 16718 47124 16770
rect 47068 16716 47124 16718
rect 46844 15314 46900 15316
rect 46844 15262 46846 15314
rect 46846 15262 46898 15314
rect 46898 15262 46900 15314
rect 46844 15260 46900 15262
rect 47852 22988 47908 23044
rect 48636 23042 48692 23044
rect 48636 22990 48638 23042
rect 48638 22990 48690 23042
rect 48690 22990 48692 23042
rect 48636 22988 48692 22990
rect 48076 22876 48132 22932
rect 47852 22092 47908 22148
rect 48076 22316 48132 22372
rect 48188 22204 48244 22260
rect 47740 21586 47796 21588
rect 47740 21534 47742 21586
rect 47742 21534 47794 21586
rect 47794 21534 47796 21586
rect 47740 21532 47796 21534
rect 48300 21532 48356 21588
rect 48300 20636 48356 20692
rect 48412 20748 48468 20804
rect 47628 20188 47684 20244
rect 48412 20188 48468 20244
rect 48524 20300 48580 20356
rect 48076 19964 48132 20020
rect 48636 19852 48692 19908
rect 48188 18620 48244 18676
rect 47852 18396 47908 18452
rect 47516 17666 47572 17668
rect 47516 17614 47518 17666
rect 47518 17614 47570 17666
rect 47570 17614 47572 17666
rect 47516 17612 47572 17614
rect 47740 17442 47796 17444
rect 47740 17390 47742 17442
rect 47742 17390 47794 17442
rect 47794 17390 47796 17442
rect 47740 17388 47796 17390
rect 47628 17106 47684 17108
rect 47628 17054 47630 17106
rect 47630 17054 47682 17106
rect 47682 17054 47684 17106
rect 47628 17052 47684 17054
rect 47404 16940 47460 16996
rect 47628 16268 47684 16324
rect 47292 15708 47348 15764
rect 48636 17106 48692 17108
rect 48636 17054 48638 17106
rect 48638 17054 48690 17106
rect 48690 17054 48692 17106
rect 48636 17052 48692 17054
rect 48188 16940 48244 16996
rect 49512 24330 49568 24332
rect 49512 24278 49514 24330
rect 49514 24278 49566 24330
rect 49566 24278 49568 24330
rect 49512 24276 49568 24278
rect 49616 24330 49672 24332
rect 49616 24278 49618 24330
rect 49618 24278 49670 24330
rect 49670 24278 49672 24330
rect 49616 24276 49672 24278
rect 49720 24330 49776 24332
rect 49720 24278 49722 24330
rect 49722 24278 49774 24330
rect 49774 24278 49776 24330
rect 49720 24276 49776 24278
rect 49308 24050 49364 24052
rect 49308 23998 49310 24050
rect 49310 23998 49362 24050
rect 49362 23998 49364 24050
rect 49308 23996 49364 23998
rect 49756 24108 49812 24164
rect 50316 24108 50372 24164
rect 49868 23996 49924 24052
rect 49980 23660 50036 23716
rect 49512 22762 49568 22764
rect 49512 22710 49514 22762
rect 49514 22710 49566 22762
rect 49566 22710 49568 22762
rect 49512 22708 49568 22710
rect 49616 22762 49672 22764
rect 49616 22710 49618 22762
rect 49618 22710 49670 22762
rect 49670 22710 49672 22762
rect 49616 22708 49672 22710
rect 49720 22762 49776 22764
rect 49720 22710 49722 22762
rect 49722 22710 49774 22762
rect 49774 22710 49776 22762
rect 49720 22708 49776 22710
rect 49532 22594 49588 22596
rect 49532 22542 49534 22594
rect 49534 22542 49586 22594
rect 49586 22542 49588 22594
rect 49532 22540 49588 22542
rect 50092 23436 50148 23492
rect 50988 23436 51044 23492
rect 49420 22370 49476 22372
rect 49420 22318 49422 22370
rect 49422 22318 49474 22370
rect 49474 22318 49476 22370
rect 49420 22316 49476 22318
rect 49980 22092 50036 22148
rect 50988 22652 51044 22708
rect 50204 21868 50260 21924
rect 50316 21644 50372 21700
rect 49868 21586 49924 21588
rect 49868 21534 49870 21586
rect 49870 21534 49922 21586
rect 49922 21534 49924 21586
rect 49868 21532 49924 21534
rect 49512 21194 49568 21196
rect 49512 21142 49514 21194
rect 49514 21142 49566 21194
rect 49566 21142 49568 21194
rect 49512 21140 49568 21142
rect 49616 21194 49672 21196
rect 49616 21142 49618 21194
rect 49618 21142 49670 21194
rect 49670 21142 49672 21194
rect 49616 21140 49672 21142
rect 49720 21194 49776 21196
rect 49720 21142 49722 21194
rect 49722 21142 49774 21194
rect 49774 21142 49776 21194
rect 49720 21140 49776 21142
rect 49644 20802 49700 20804
rect 49644 20750 49646 20802
rect 49646 20750 49698 20802
rect 49698 20750 49700 20802
rect 49644 20748 49700 20750
rect 50092 20300 50148 20356
rect 49532 20018 49588 20020
rect 49532 19966 49534 20018
rect 49534 19966 49586 20018
rect 49586 19966 49588 20018
rect 49532 19964 49588 19966
rect 49512 19626 49568 19628
rect 49512 19574 49514 19626
rect 49514 19574 49566 19626
rect 49566 19574 49568 19626
rect 49512 19572 49568 19574
rect 49616 19626 49672 19628
rect 49616 19574 49618 19626
rect 49618 19574 49670 19626
rect 49670 19574 49672 19626
rect 49616 19572 49672 19574
rect 49720 19626 49776 19628
rect 49720 19574 49722 19626
rect 49722 19574 49774 19626
rect 49774 19574 49776 19626
rect 49720 19572 49776 19574
rect 49644 19404 49700 19460
rect 49308 18732 49364 18788
rect 48972 16716 49028 16772
rect 48524 16098 48580 16100
rect 48524 16046 48526 16098
rect 48526 16046 48578 16098
rect 48578 16046 48580 16098
rect 48524 16044 48580 16046
rect 48076 14588 48132 14644
rect 46172 13858 46228 13860
rect 46172 13806 46174 13858
rect 46174 13806 46226 13858
rect 46226 13806 46228 13858
rect 46172 13804 46228 13806
rect 42028 13020 42084 13076
rect 40796 12962 40852 12964
rect 40796 12910 40798 12962
rect 40798 12910 40850 12962
rect 40850 12910 40852 12962
rect 40796 12908 40852 12910
rect 42476 12962 42532 12964
rect 42476 12910 42478 12962
rect 42478 12910 42530 12962
rect 42530 12910 42532 12962
rect 42476 12908 42532 12910
rect 40460 12236 40516 12292
rect 43596 12908 43652 12964
rect 45948 13580 46004 13636
rect 46844 13356 46900 13412
rect 44940 12908 44996 12964
rect 45836 12962 45892 12964
rect 45836 12910 45838 12962
rect 45838 12910 45890 12962
rect 45890 12910 45892 12962
rect 45836 12908 45892 12910
rect 44492 12796 44548 12852
rect 44268 12684 44324 12740
rect 42588 12066 42644 12068
rect 42588 12014 42590 12066
rect 42590 12014 42642 12066
rect 42642 12014 42644 12066
rect 42588 12012 42644 12014
rect 43932 12124 43988 12180
rect 43596 12012 43652 12068
rect 41916 11452 41972 11508
rect 43932 11564 43988 11620
rect 43596 11116 43652 11172
rect 46060 12850 46116 12852
rect 46060 12798 46062 12850
rect 46062 12798 46114 12850
rect 46114 12798 46116 12850
rect 46060 12796 46116 12798
rect 45612 12738 45668 12740
rect 45612 12686 45614 12738
rect 45614 12686 45666 12738
rect 45666 12686 45668 12738
rect 45612 12684 45668 12686
rect 45388 12236 45444 12292
rect 42252 10668 42308 10724
rect 44268 11170 44324 11172
rect 44268 11118 44270 11170
rect 44270 11118 44322 11170
rect 44322 11118 44324 11170
rect 44268 11116 44324 11118
rect 40572 10556 40628 10612
rect 40796 10610 40852 10612
rect 40796 10558 40798 10610
rect 40798 10558 40850 10610
rect 40850 10558 40852 10610
rect 40796 10556 40852 10558
rect 41468 10498 41524 10500
rect 41468 10446 41470 10498
rect 41470 10446 41522 10498
rect 41522 10446 41524 10498
rect 41468 10444 41524 10446
rect 40460 10108 40516 10164
rect 40572 9772 40628 9828
rect 40348 9548 40404 9604
rect 40684 9266 40740 9268
rect 40684 9214 40686 9266
rect 40686 9214 40738 9266
rect 40738 9214 40740 9266
rect 40684 9212 40740 9214
rect 40460 8764 40516 8820
rect 40572 9154 40628 9156
rect 40572 9102 40574 9154
rect 40574 9102 40626 9154
rect 40626 9102 40628 9154
rect 40572 9100 40628 9102
rect 40908 9042 40964 9044
rect 40908 8990 40910 9042
rect 40910 8990 40962 9042
rect 40962 8990 40964 9042
rect 40908 8988 40964 8990
rect 40572 8540 40628 8596
rect 41356 9826 41412 9828
rect 41356 9774 41358 9826
rect 41358 9774 41410 9826
rect 41410 9774 41412 9826
rect 41356 9772 41412 9774
rect 41580 9042 41636 9044
rect 41580 8990 41582 9042
rect 41582 8990 41634 9042
rect 41634 8990 41636 9042
rect 41580 8988 41636 8990
rect 42140 9602 42196 9604
rect 42140 9550 42142 9602
rect 42142 9550 42194 9602
rect 42194 9550 42196 9602
rect 42140 9548 42196 9550
rect 42476 10386 42532 10388
rect 42476 10334 42478 10386
rect 42478 10334 42530 10386
rect 42530 10334 42532 10386
rect 42476 10332 42532 10334
rect 42812 10386 42868 10388
rect 42812 10334 42814 10386
rect 42814 10334 42866 10386
rect 42866 10334 42868 10386
rect 42812 10332 42868 10334
rect 43820 10610 43876 10612
rect 43820 10558 43822 10610
rect 43822 10558 43874 10610
rect 43874 10558 43876 10610
rect 43820 10556 43876 10558
rect 44044 10498 44100 10500
rect 44044 10446 44046 10498
rect 44046 10446 44098 10498
rect 44098 10446 44100 10498
rect 44044 10444 44100 10446
rect 45276 10610 45332 10612
rect 45276 10558 45278 10610
rect 45278 10558 45330 10610
rect 45330 10558 45332 10610
rect 45276 10556 45332 10558
rect 45500 10444 45556 10500
rect 44716 9826 44772 9828
rect 44716 9774 44718 9826
rect 44718 9774 44770 9826
rect 44770 9774 44772 9826
rect 44716 9772 44772 9774
rect 45724 9826 45780 9828
rect 45724 9774 45726 9826
rect 45726 9774 45778 9826
rect 45778 9774 45780 9826
rect 45724 9772 45780 9774
rect 42364 9548 42420 9604
rect 42364 9100 42420 9156
rect 40796 8316 40852 8372
rect 41692 8764 41748 8820
rect 41692 8540 41748 8596
rect 41580 8316 41636 8372
rect 40684 7868 40740 7924
rect 39564 7084 39620 7140
rect 39340 6524 39396 6580
rect 39340 5852 39396 5908
rect 39676 6690 39732 6692
rect 39676 6638 39678 6690
rect 39678 6638 39730 6690
rect 39730 6638 39732 6690
rect 39676 6636 39732 6638
rect 40124 6524 40180 6580
rect 41356 6690 41412 6692
rect 41356 6638 41358 6690
rect 41358 6638 41410 6690
rect 41410 6638 41412 6690
rect 41356 6636 41412 6638
rect 40348 6412 40404 6468
rect 39676 6300 39732 6356
rect 39564 5906 39620 5908
rect 39564 5854 39566 5906
rect 39566 5854 39618 5906
rect 39618 5854 39620 5906
rect 39564 5852 39620 5854
rect 39852 6298 39908 6300
rect 39852 6246 39854 6298
rect 39854 6246 39906 6298
rect 39906 6246 39908 6298
rect 39852 6244 39908 6246
rect 39956 6298 40012 6300
rect 39956 6246 39958 6298
rect 39958 6246 40010 6298
rect 40010 6246 40012 6298
rect 39956 6244 40012 6246
rect 40060 6298 40116 6300
rect 40060 6246 40062 6298
rect 40062 6246 40114 6298
rect 40114 6246 40116 6298
rect 40060 6244 40116 6246
rect 39116 5234 39172 5236
rect 39116 5182 39118 5234
rect 39118 5182 39170 5234
rect 39170 5182 39172 5234
rect 39116 5180 39172 5182
rect 38892 5068 38948 5124
rect 39004 5010 39060 5012
rect 39004 4958 39006 5010
rect 39006 4958 39058 5010
rect 39058 4958 39060 5010
rect 39004 4956 39060 4958
rect 38668 4226 38724 4228
rect 38668 4174 38670 4226
rect 38670 4174 38722 4226
rect 38722 4174 38724 4226
rect 38668 4172 38724 4174
rect 39116 4508 39172 4564
rect 39452 4844 39508 4900
rect 39228 4172 39284 4228
rect 38220 3554 38276 3556
rect 38220 3502 38222 3554
rect 38222 3502 38274 3554
rect 38274 3502 38276 3554
rect 38220 3500 38276 3502
rect 41244 6466 41300 6468
rect 41244 6414 41246 6466
rect 41246 6414 41298 6466
rect 41298 6414 41300 6466
rect 41244 6412 41300 6414
rect 40796 5906 40852 5908
rect 40796 5854 40798 5906
rect 40798 5854 40850 5906
rect 40850 5854 40852 5906
rect 40796 5852 40852 5854
rect 42700 9602 42756 9604
rect 42700 9550 42702 9602
rect 42702 9550 42754 9602
rect 42754 9550 42756 9602
rect 42700 9548 42756 9550
rect 42252 8876 42308 8932
rect 43260 9602 43316 9604
rect 43260 9550 43262 9602
rect 43262 9550 43314 9602
rect 43314 9550 43316 9602
rect 43260 9548 43316 9550
rect 44604 9714 44660 9716
rect 44604 9662 44606 9714
rect 44606 9662 44658 9714
rect 44658 9662 44660 9714
rect 44604 9660 44660 9662
rect 43484 9436 43540 9492
rect 43932 9436 43988 9492
rect 42700 8652 42756 8708
rect 42924 9324 42980 9380
rect 43036 9266 43092 9268
rect 43036 9214 43038 9266
rect 43038 9214 43090 9266
rect 43090 9214 43092 9266
rect 43036 9212 43092 9214
rect 44044 9266 44100 9268
rect 44044 9214 44046 9266
rect 44046 9214 44098 9266
rect 44098 9214 44100 9266
rect 44044 9212 44100 9214
rect 43260 8652 43316 8708
rect 42924 8428 42980 8484
rect 45388 9548 45444 9604
rect 45276 9212 45332 9268
rect 45276 8764 45332 8820
rect 43484 8258 43540 8260
rect 43484 8206 43486 8258
rect 43486 8206 43538 8258
rect 43538 8206 43540 8258
rect 43484 8204 43540 8206
rect 43260 7868 43316 7924
rect 42028 7644 42084 7700
rect 45948 9660 46004 9716
rect 46284 8258 46340 8260
rect 46284 8206 46286 8258
rect 46286 8206 46338 8258
rect 46338 8206 46340 8258
rect 46284 8204 46340 8206
rect 46732 8258 46788 8260
rect 46732 8206 46734 8258
rect 46734 8206 46786 8258
rect 46786 8206 46788 8258
rect 46732 8204 46788 8206
rect 45388 8092 45444 8148
rect 42924 7420 42980 7476
rect 42812 7196 42868 7252
rect 42588 6690 42644 6692
rect 42588 6638 42590 6690
rect 42590 6638 42642 6690
rect 42642 6638 42644 6690
rect 42588 6636 42644 6638
rect 40348 5180 40404 5236
rect 40460 5292 40516 5348
rect 39788 5068 39844 5124
rect 40124 4956 40180 5012
rect 41020 5122 41076 5124
rect 41020 5070 41022 5122
rect 41022 5070 41074 5122
rect 41074 5070 41076 5122
rect 41020 5068 41076 5070
rect 40348 4898 40404 4900
rect 40348 4846 40350 4898
rect 40350 4846 40402 4898
rect 40402 4846 40404 4898
rect 40348 4844 40404 4846
rect 39852 4730 39908 4732
rect 39852 4678 39854 4730
rect 39854 4678 39906 4730
rect 39906 4678 39908 4730
rect 39852 4676 39908 4678
rect 39956 4730 40012 4732
rect 39956 4678 39958 4730
rect 39958 4678 40010 4730
rect 40010 4678 40012 4730
rect 39956 4676 40012 4678
rect 40060 4730 40116 4732
rect 40060 4678 40062 4730
rect 40062 4678 40114 4730
rect 40114 4678 40116 4730
rect 40060 4676 40116 4678
rect 40236 4732 40292 4788
rect 41468 4732 41524 4788
rect 41804 4956 41860 5012
rect 41356 4620 41412 4676
rect 40460 4508 40516 4564
rect 40348 4450 40404 4452
rect 40348 4398 40350 4450
rect 40350 4398 40402 4450
rect 40402 4398 40404 4450
rect 40348 4396 40404 4398
rect 41356 4284 41412 4340
rect 41580 4620 41636 4676
rect 40236 3948 40292 4004
rect 37660 1596 37716 1652
rect 37548 812 37604 868
rect 40124 3500 40180 3556
rect 39452 3442 39508 3444
rect 39452 3390 39454 3442
rect 39454 3390 39506 3442
rect 39506 3390 39508 3442
rect 39452 3388 39508 3390
rect 40236 3388 40292 3444
rect 41692 4562 41748 4564
rect 41692 4510 41694 4562
rect 41694 4510 41746 4562
rect 41746 4510 41748 4562
rect 41692 4508 41748 4510
rect 41916 4898 41972 4900
rect 41916 4846 41918 4898
rect 41918 4846 41970 4898
rect 41970 4846 41972 4898
rect 41916 4844 41972 4846
rect 42140 5906 42196 5908
rect 42140 5854 42142 5906
rect 42142 5854 42194 5906
rect 42194 5854 42196 5906
rect 42140 5852 42196 5854
rect 42028 4620 42084 4676
rect 42140 5404 42196 5460
rect 42476 5628 42532 5684
rect 42252 4844 42308 4900
rect 42252 4450 42308 4452
rect 42252 4398 42254 4450
rect 42254 4398 42306 4450
rect 42306 4398 42308 4450
rect 42252 4396 42308 4398
rect 42364 4732 42420 4788
rect 41804 4338 41860 4340
rect 41804 4286 41806 4338
rect 41806 4286 41858 4338
rect 41858 4286 41860 4338
rect 41804 4284 41860 4286
rect 43932 7420 43988 7476
rect 43036 7308 43092 7364
rect 43484 6802 43540 6804
rect 43484 6750 43486 6802
rect 43486 6750 43538 6802
rect 43538 6750 43540 6802
rect 43484 6748 43540 6750
rect 42924 6188 42980 6244
rect 42924 5404 42980 5460
rect 42700 4562 42756 4564
rect 42700 4510 42702 4562
rect 42702 4510 42754 4562
rect 42754 4510 42756 4562
rect 42700 4508 42756 4510
rect 42364 4284 42420 4340
rect 42924 3778 42980 3780
rect 42924 3726 42926 3778
rect 42926 3726 42978 3778
rect 42978 3726 42980 3778
rect 42924 3724 42980 3726
rect 41580 3612 41636 3668
rect 39852 3162 39908 3164
rect 39852 3110 39854 3162
rect 39854 3110 39906 3162
rect 39906 3110 39908 3162
rect 39852 3108 39908 3110
rect 39956 3162 40012 3164
rect 39956 3110 39958 3162
rect 39958 3110 40010 3162
rect 40010 3110 40012 3162
rect 39956 3108 40012 3110
rect 40060 3162 40116 3164
rect 40060 3110 40062 3162
rect 40062 3110 40114 3162
rect 40114 3110 40116 3162
rect 40060 3108 40116 3110
rect 41244 3442 41300 3444
rect 41244 3390 41246 3442
rect 41246 3390 41298 3442
rect 41298 3390 41300 3442
rect 41244 3388 41300 3390
rect 40236 2044 40292 2100
rect 42812 3612 42868 3668
rect 42028 3442 42084 3444
rect 42028 3390 42030 3442
rect 42030 3390 42082 3442
rect 42082 3390 42084 3442
rect 42028 3388 42084 3390
rect 42924 3164 42980 3220
rect 43036 924 43092 980
rect 43372 4732 43428 4788
rect 43596 4844 43652 4900
rect 43596 2828 43652 2884
rect 43708 4732 43764 4788
rect 43708 1484 43764 1540
rect 44492 7308 44548 7364
rect 44156 6748 44212 6804
rect 44604 6300 44660 6356
rect 44828 5180 44884 5236
rect 44268 4898 44324 4900
rect 44268 4846 44270 4898
rect 44270 4846 44322 4898
rect 44322 4846 44324 4898
rect 44268 4844 44324 4846
rect 44156 4732 44212 4788
rect 44156 4508 44212 4564
rect 44044 4284 44100 4340
rect 48412 15314 48468 15316
rect 48412 15262 48414 15314
rect 48414 15262 48466 15314
rect 48466 15262 48468 15314
rect 48412 15260 48468 15262
rect 49868 19292 49924 19348
rect 50988 19964 51044 20020
rect 51100 19292 51156 19348
rect 49868 18732 49924 18788
rect 50204 18956 50260 19012
rect 49756 18674 49812 18676
rect 49756 18622 49758 18674
rect 49758 18622 49810 18674
rect 49810 18622 49812 18674
rect 49756 18620 49812 18622
rect 50764 19010 50820 19012
rect 50764 18958 50766 19010
rect 50766 18958 50818 19010
rect 50818 18958 50820 19010
rect 50764 18956 50820 18958
rect 50316 18844 50372 18900
rect 49512 18058 49568 18060
rect 49512 18006 49514 18058
rect 49514 18006 49566 18058
rect 49566 18006 49568 18058
rect 49512 18004 49568 18006
rect 49616 18058 49672 18060
rect 49616 18006 49618 18058
rect 49618 18006 49670 18058
rect 49670 18006 49672 18058
rect 49616 18004 49672 18006
rect 49720 18058 49776 18060
rect 49720 18006 49722 18058
rect 49722 18006 49774 18058
rect 49774 18006 49776 18058
rect 49720 18004 49776 18006
rect 49980 17836 50036 17892
rect 49420 16940 49476 16996
rect 50876 18732 50932 18788
rect 50652 18450 50708 18452
rect 50652 18398 50654 18450
rect 50654 18398 50706 18450
rect 50706 18398 50708 18450
rect 50652 18396 50708 18398
rect 50316 17612 50372 17668
rect 50764 17554 50820 17556
rect 50764 17502 50766 17554
rect 50766 17502 50818 17554
rect 50818 17502 50820 17554
rect 50764 17500 50820 17502
rect 49756 16716 49812 16772
rect 50540 17388 50596 17444
rect 50092 16716 50148 16772
rect 49512 16490 49568 16492
rect 49512 16438 49514 16490
rect 49514 16438 49566 16490
rect 49566 16438 49568 16490
rect 49512 16436 49568 16438
rect 49616 16490 49672 16492
rect 49616 16438 49618 16490
rect 49618 16438 49670 16490
rect 49670 16438 49672 16490
rect 49616 16436 49672 16438
rect 49720 16490 49776 16492
rect 49720 16438 49722 16490
rect 49722 16438 49774 16490
rect 49774 16438 49776 16490
rect 49720 16436 49776 16438
rect 49868 16268 49924 16324
rect 49420 16098 49476 16100
rect 49420 16046 49422 16098
rect 49422 16046 49474 16098
rect 49474 16046 49476 16098
rect 49420 16044 49476 16046
rect 49980 15260 50036 15316
rect 50428 15820 50484 15876
rect 49512 14922 49568 14924
rect 49512 14870 49514 14922
rect 49514 14870 49566 14922
rect 49566 14870 49568 14922
rect 49512 14868 49568 14870
rect 49616 14922 49672 14924
rect 49616 14870 49618 14922
rect 49618 14870 49670 14922
rect 49670 14870 49672 14922
rect 49616 14868 49672 14870
rect 49720 14922 49776 14924
rect 49720 14870 49722 14922
rect 49722 14870 49774 14922
rect 49774 14870 49776 14922
rect 49720 14868 49776 14870
rect 48412 14252 48468 14308
rect 48748 14028 48804 14084
rect 50316 14418 50372 14420
rect 50316 14366 50318 14418
rect 50318 14366 50370 14418
rect 50370 14366 50372 14418
rect 50316 14364 50372 14366
rect 50092 14028 50148 14084
rect 50652 16716 50708 16772
rect 51100 18396 51156 18452
rect 50988 16882 51044 16884
rect 50988 16830 50990 16882
rect 50990 16830 51042 16882
rect 51042 16830 51044 16882
rect 50988 16828 51044 16830
rect 50876 16716 50932 16772
rect 50652 15426 50708 15428
rect 50652 15374 50654 15426
rect 50654 15374 50706 15426
rect 50706 15374 50708 15426
rect 50652 15372 50708 15374
rect 50540 15260 50596 15316
rect 50876 15820 50932 15876
rect 50764 15148 50820 15204
rect 51436 30940 51492 30996
rect 51548 30828 51604 30884
rect 51324 29148 51380 29204
rect 51436 28588 51492 28644
rect 52220 31666 52276 31668
rect 52220 31614 52222 31666
rect 52222 31614 52274 31666
rect 52274 31614 52276 31666
rect 52220 31612 52276 31614
rect 51772 31554 51828 31556
rect 51772 31502 51774 31554
rect 51774 31502 51826 31554
rect 51826 31502 51828 31554
rect 51772 31500 51828 31502
rect 55356 35698 55412 35700
rect 55356 35646 55358 35698
rect 55358 35646 55410 35698
rect 55410 35646 55412 35698
rect 55356 35644 55412 35646
rect 55916 35698 55972 35700
rect 55916 35646 55918 35698
rect 55918 35646 55970 35698
rect 55970 35646 55972 35698
rect 55916 35644 55972 35646
rect 55132 34242 55188 34244
rect 55132 34190 55134 34242
rect 55134 34190 55186 34242
rect 55186 34190 55188 34242
rect 55132 34188 55188 34190
rect 56028 35196 56084 35252
rect 58044 35644 58100 35700
rect 56588 35586 56644 35588
rect 56588 35534 56590 35586
rect 56590 35534 56642 35586
rect 56642 35534 56644 35586
rect 56588 35532 56644 35534
rect 57484 35586 57540 35588
rect 57484 35534 57486 35586
rect 57486 35534 57538 35586
rect 57538 35534 57540 35586
rect 57484 35532 57540 35534
rect 57036 35420 57092 35476
rect 57708 35474 57764 35476
rect 57708 35422 57710 35474
rect 57710 35422 57762 35474
rect 57762 35422 57764 35474
rect 57708 35420 57764 35422
rect 57260 35196 57316 35252
rect 55916 34748 55972 34804
rect 56812 34802 56868 34804
rect 56812 34750 56814 34802
rect 56814 34750 56866 34802
rect 56866 34750 56868 34802
rect 56812 34748 56868 34750
rect 55692 33964 55748 34020
rect 54908 33906 54964 33908
rect 54908 33854 54910 33906
rect 54910 33854 54962 33906
rect 54962 33854 54964 33906
rect 54908 33852 54964 33854
rect 53900 33180 53956 33236
rect 53788 32620 53844 32676
rect 52780 31500 52836 31556
rect 53788 32450 53844 32452
rect 53788 32398 53790 32450
rect 53790 32398 53842 32450
rect 53842 32398 53844 32450
rect 53788 32396 53844 32398
rect 52444 30882 52500 30884
rect 52444 30830 52446 30882
rect 52446 30830 52498 30882
rect 52498 30830 52500 30882
rect 52444 30828 52500 30830
rect 52444 29596 52500 29652
rect 54124 31948 54180 32004
rect 54012 31612 54068 31668
rect 53788 31388 53844 31444
rect 53900 31554 53956 31556
rect 53900 31502 53902 31554
rect 53902 31502 53954 31554
rect 53954 31502 53956 31554
rect 53900 31500 53956 31502
rect 56588 33346 56644 33348
rect 56588 33294 56590 33346
rect 56590 33294 56642 33346
rect 56642 33294 56644 33346
rect 56588 33292 56644 33294
rect 57148 33180 57204 33236
rect 54572 31948 54628 32004
rect 55692 32562 55748 32564
rect 55692 32510 55694 32562
rect 55694 32510 55746 32562
rect 55746 32510 55748 32562
rect 55692 32508 55748 32510
rect 55356 31948 55412 32004
rect 54012 31052 54068 31108
rect 53564 30268 53620 30324
rect 54236 30994 54292 30996
rect 54236 30942 54238 30994
rect 54238 30942 54290 30994
rect 54290 30942 54292 30994
rect 54236 30940 54292 30942
rect 54236 30716 54292 30772
rect 54684 30882 54740 30884
rect 54684 30830 54686 30882
rect 54686 30830 54738 30882
rect 54738 30830 54740 30882
rect 54684 30828 54740 30830
rect 55580 31724 55636 31780
rect 55356 31106 55412 31108
rect 55356 31054 55358 31106
rect 55358 31054 55410 31106
rect 55410 31054 55412 31106
rect 55356 31052 55412 31054
rect 54796 30716 54852 30772
rect 55356 30492 55412 30548
rect 56364 32562 56420 32564
rect 56364 32510 56366 32562
rect 56366 32510 56418 32562
rect 56418 32510 56420 32562
rect 56364 32508 56420 32510
rect 56140 31778 56196 31780
rect 56140 31726 56142 31778
rect 56142 31726 56194 31778
rect 56194 31726 56196 31778
rect 56140 31724 56196 31726
rect 55916 31500 55972 31556
rect 55580 30828 55636 30884
rect 55916 30716 55972 30772
rect 55692 30268 55748 30324
rect 56812 31666 56868 31668
rect 56812 31614 56814 31666
rect 56814 31614 56866 31666
rect 56866 31614 56868 31666
rect 56812 31612 56868 31614
rect 57260 31554 57316 31556
rect 57260 31502 57262 31554
rect 57262 31502 57314 31554
rect 57314 31502 57316 31554
rect 57260 31500 57316 31502
rect 54796 30156 54852 30212
rect 54684 30098 54740 30100
rect 54684 30046 54686 30098
rect 54686 30046 54738 30098
rect 54738 30046 54740 30098
rect 54684 30044 54740 30046
rect 55692 30098 55748 30100
rect 55692 30046 55694 30098
rect 55694 30046 55746 30098
rect 55746 30046 55748 30098
rect 55692 30044 55748 30046
rect 53452 29820 53508 29876
rect 54012 29820 54068 29876
rect 55580 29986 55636 29988
rect 55580 29934 55582 29986
rect 55582 29934 55634 29986
rect 55634 29934 55636 29986
rect 55580 29932 55636 29934
rect 54796 29820 54852 29876
rect 51884 29148 51940 29204
rect 52668 29148 52724 29204
rect 52332 28754 52388 28756
rect 52332 28702 52334 28754
rect 52334 28702 52386 28754
rect 52386 28702 52388 28754
rect 52332 28700 52388 28702
rect 52444 27916 52500 27972
rect 54908 29538 54964 29540
rect 54908 29486 54910 29538
rect 54910 29486 54962 29538
rect 54962 29486 54964 29538
rect 54908 29484 54964 29486
rect 54572 29426 54628 29428
rect 54572 29374 54574 29426
rect 54574 29374 54626 29426
rect 54626 29374 54628 29426
rect 54572 29372 54628 29374
rect 53004 28700 53060 28756
rect 53116 28476 53172 28532
rect 52892 27692 52948 27748
rect 53564 28140 53620 28196
rect 54012 28364 54068 28420
rect 54572 28530 54628 28532
rect 54572 28478 54574 28530
rect 54574 28478 54626 28530
rect 54626 28478 54628 28530
rect 54572 28476 54628 28478
rect 54460 28364 54516 28420
rect 51436 22428 51492 22484
rect 51772 22258 51828 22260
rect 51772 22206 51774 22258
rect 51774 22206 51826 22258
rect 51826 22206 51828 22258
rect 51772 22204 51828 22206
rect 52332 26850 52388 26852
rect 52332 26798 52334 26850
rect 52334 26798 52386 26850
rect 52386 26798 52388 26850
rect 52332 26796 52388 26798
rect 54348 28140 54404 28196
rect 55468 28418 55524 28420
rect 55468 28366 55470 28418
rect 55470 28366 55522 28418
rect 55522 28366 55524 28418
rect 55468 28364 55524 28366
rect 54572 27970 54628 27972
rect 54572 27918 54574 27970
rect 54574 27918 54626 27970
rect 54626 27918 54628 27970
rect 54572 27916 54628 27918
rect 54684 27692 54740 27748
rect 53788 27244 53844 27300
rect 53564 27020 53620 27076
rect 52668 26460 52724 26516
rect 52780 26572 52836 26628
rect 52668 26290 52724 26292
rect 52668 26238 52670 26290
rect 52670 26238 52722 26290
rect 52722 26238 52724 26290
rect 52668 26236 52724 26238
rect 53564 26572 53620 26628
rect 53452 26460 53508 26516
rect 52556 23714 52612 23716
rect 52556 23662 52558 23714
rect 52558 23662 52610 23714
rect 52610 23662 52612 23714
rect 52556 23660 52612 23662
rect 52220 22540 52276 22596
rect 52556 23324 52612 23380
rect 51884 21868 51940 21924
rect 51324 18732 51380 18788
rect 51660 18674 51716 18676
rect 51660 18622 51662 18674
rect 51662 18622 51714 18674
rect 51714 18622 51716 18674
rect 51660 18620 51716 18622
rect 51436 18284 51492 18340
rect 51212 18172 51268 18228
rect 51212 17724 51268 17780
rect 51436 17554 51492 17556
rect 51436 17502 51438 17554
rect 51438 17502 51490 17554
rect 51490 17502 51492 17554
rect 51436 17500 51492 17502
rect 51324 17276 51380 17332
rect 51660 17052 51716 17108
rect 51884 16940 51940 16996
rect 51884 16770 51940 16772
rect 51884 16718 51886 16770
rect 51886 16718 51938 16770
rect 51938 16718 51940 16770
rect 51884 16716 51940 16718
rect 51212 15426 51268 15428
rect 51212 15374 51214 15426
rect 51214 15374 51266 15426
rect 51266 15374 51268 15426
rect 51212 15372 51268 15374
rect 51660 15314 51716 15316
rect 51660 15262 51662 15314
rect 51662 15262 51714 15314
rect 51714 15262 51716 15314
rect 51660 15260 51716 15262
rect 52108 21756 52164 21812
rect 50764 14418 50820 14420
rect 50764 14366 50766 14418
rect 50766 14366 50818 14418
rect 50818 14366 50820 14418
rect 50764 14364 50820 14366
rect 50876 14306 50932 14308
rect 50876 14254 50878 14306
rect 50878 14254 50930 14306
rect 50930 14254 50932 14306
rect 50876 14252 50932 14254
rect 50428 13804 50484 13860
rect 48636 13580 48692 13636
rect 48300 13356 48356 13412
rect 49980 13580 50036 13636
rect 49512 13354 49568 13356
rect 49512 13302 49514 13354
rect 49514 13302 49566 13354
rect 49566 13302 49568 13354
rect 49512 13300 49568 13302
rect 49616 13354 49672 13356
rect 49616 13302 49618 13354
rect 49618 13302 49670 13354
rect 49670 13302 49672 13354
rect 49616 13300 49672 13302
rect 49720 13354 49776 13356
rect 49720 13302 49722 13354
rect 49722 13302 49774 13354
rect 49774 13302 49776 13354
rect 49720 13300 49776 13302
rect 50988 13074 51044 13076
rect 50988 13022 50990 13074
rect 50990 13022 51042 13074
rect 51042 13022 51044 13074
rect 50988 13020 51044 13022
rect 49644 12962 49700 12964
rect 49644 12910 49646 12962
rect 49646 12910 49698 12962
rect 49698 12910 49700 12962
rect 49644 12908 49700 12910
rect 50092 12796 50148 12852
rect 48860 12684 48916 12740
rect 48636 12290 48692 12292
rect 48636 12238 48638 12290
rect 48638 12238 48690 12290
rect 48690 12238 48692 12290
rect 48636 12236 48692 12238
rect 49756 12236 49812 12292
rect 48412 12012 48468 12068
rect 48188 11788 48244 11844
rect 46956 11340 47012 11396
rect 47292 10668 47348 10724
rect 47516 10668 47572 10724
rect 47404 8258 47460 8260
rect 47404 8206 47406 8258
rect 47406 8206 47458 8258
rect 47458 8206 47460 8258
rect 47404 8204 47460 8206
rect 47628 8146 47684 8148
rect 47628 8094 47630 8146
rect 47630 8094 47682 8146
rect 47682 8094 47684 8146
rect 47628 8092 47684 8094
rect 46844 7756 46900 7812
rect 45388 7196 45444 7252
rect 45948 6748 46004 6804
rect 49868 12066 49924 12068
rect 49868 12014 49870 12066
rect 49870 12014 49922 12066
rect 49922 12014 49924 12066
rect 49868 12012 49924 12014
rect 50876 12908 50932 12964
rect 50652 12738 50708 12740
rect 50652 12686 50654 12738
rect 50654 12686 50706 12738
rect 50706 12686 50708 12738
rect 50652 12684 50708 12686
rect 51100 12850 51156 12852
rect 51100 12798 51102 12850
rect 51102 12798 51154 12850
rect 51154 12798 51156 12850
rect 51100 12796 51156 12798
rect 51324 12796 51380 12852
rect 50876 12236 50932 12292
rect 51324 12124 51380 12180
rect 49512 11786 49568 11788
rect 49512 11734 49514 11786
rect 49514 11734 49566 11786
rect 49566 11734 49568 11786
rect 49512 11732 49568 11734
rect 49616 11786 49672 11788
rect 49616 11734 49618 11786
rect 49618 11734 49670 11786
rect 49670 11734 49672 11786
rect 49616 11732 49672 11734
rect 49720 11786 49776 11788
rect 49720 11734 49722 11786
rect 49722 11734 49774 11786
rect 49774 11734 49776 11786
rect 49720 11732 49776 11734
rect 48860 11394 48916 11396
rect 48860 11342 48862 11394
rect 48862 11342 48914 11394
rect 48914 11342 48916 11394
rect 48860 11340 48916 11342
rect 48748 11282 48804 11284
rect 48748 11230 48750 11282
rect 48750 11230 48802 11282
rect 48802 11230 48804 11282
rect 48748 11228 48804 11230
rect 51548 11394 51604 11396
rect 51548 11342 51550 11394
rect 51550 11342 51602 11394
rect 51602 11342 51604 11394
rect 51548 11340 51604 11342
rect 50988 11170 51044 11172
rect 50988 11118 50990 11170
rect 50990 11118 51042 11170
rect 51042 11118 51044 11170
rect 50988 11116 51044 11118
rect 48636 10668 48692 10724
rect 49644 10722 49700 10724
rect 49644 10670 49646 10722
rect 49646 10670 49698 10722
rect 49698 10670 49700 10722
rect 49644 10668 49700 10670
rect 49512 10218 49568 10220
rect 49512 10166 49514 10218
rect 49514 10166 49566 10218
rect 49566 10166 49568 10218
rect 49512 10164 49568 10166
rect 49616 10218 49672 10220
rect 49616 10166 49618 10218
rect 49618 10166 49670 10218
rect 49670 10166 49672 10218
rect 49616 10164 49672 10166
rect 49720 10218 49776 10220
rect 49720 10166 49722 10218
rect 49722 10166 49774 10218
rect 49774 10166 49776 10218
rect 49720 10164 49776 10166
rect 48300 9324 48356 9380
rect 49196 9212 49252 9268
rect 48748 9154 48804 9156
rect 48748 9102 48750 9154
rect 48750 9102 48802 9154
rect 48802 9102 48804 9154
rect 48748 9100 48804 9102
rect 49420 9154 49476 9156
rect 49420 9102 49422 9154
rect 49422 9102 49474 9154
rect 49474 9102 49476 9154
rect 49420 9100 49476 9102
rect 50316 10498 50372 10500
rect 50316 10446 50318 10498
rect 50318 10446 50370 10498
rect 50370 10446 50372 10498
rect 50316 10444 50372 10446
rect 50764 10444 50820 10500
rect 50988 10332 51044 10388
rect 50764 10220 50820 10276
rect 49868 9324 49924 9380
rect 50540 9660 50596 9716
rect 49980 9266 50036 9268
rect 49980 9214 49982 9266
rect 49982 9214 50034 9266
rect 50034 9214 50036 9266
rect 49980 9212 50036 9214
rect 49756 9100 49812 9156
rect 49196 8652 49252 8708
rect 49512 8650 49568 8652
rect 49512 8598 49514 8650
rect 49514 8598 49566 8650
rect 49566 8598 49568 8650
rect 49512 8596 49568 8598
rect 49616 8650 49672 8652
rect 49616 8598 49618 8650
rect 49618 8598 49670 8650
rect 49670 8598 49672 8650
rect 49616 8596 49672 8598
rect 49720 8650 49776 8652
rect 49720 8598 49722 8650
rect 49722 8598 49774 8650
rect 49774 8598 49776 8650
rect 49720 8596 49776 8598
rect 50988 9772 51044 9828
rect 51548 9826 51604 9828
rect 51548 9774 51550 9826
rect 51550 9774 51602 9826
rect 51602 9774 51604 9826
rect 51548 9772 51604 9774
rect 50988 9548 51044 9604
rect 50876 9154 50932 9156
rect 50876 9102 50878 9154
rect 50878 9102 50930 9154
rect 50930 9102 50932 9154
rect 50876 9100 50932 9102
rect 50764 8988 50820 9044
rect 51996 14642 52052 14644
rect 51996 14590 51998 14642
rect 51998 14590 52050 14642
rect 52050 14590 52052 14642
rect 51996 14588 52052 14590
rect 51996 11116 52052 11172
rect 52444 23154 52500 23156
rect 52444 23102 52446 23154
rect 52446 23102 52498 23154
rect 52498 23102 52500 23154
rect 52444 23100 52500 23102
rect 53788 26572 53844 26628
rect 53340 25452 53396 25508
rect 54348 27132 54404 27188
rect 53900 25506 53956 25508
rect 53900 25454 53902 25506
rect 53902 25454 53954 25506
rect 53954 25454 53956 25506
rect 53900 25452 53956 25454
rect 54684 26962 54740 26964
rect 54684 26910 54686 26962
rect 54686 26910 54738 26962
rect 54738 26910 54740 26962
rect 54684 26908 54740 26910
rect 53452 23378 53508 23380
rect 53452 23326 53454 23378
rect 53454 23326 53506 23378
rect 53506 23326 53508 23378
rect 53452 23324 53508 23326
rect 53788 23660 53844 23716
rect 54348 23660 54404 23716
rect 53676 23100 53732 23156
rect 53900 22540 53956 22596
rect 55916 30156 55972 30212
rect 56364 31388 56420 31444
rect 56364 30268 56420 30324
rect 56140 30044 56196 30100
rect 56252 29820 56308 29876
rect 56028 29372 56084 29428
rect 55356 27132 55412 27188
rect 55916 26796 55972 26852
rect 55580 23154 55636 23156
rect 55580 23102 55582 23154
rect 55582 23102 55634 23154
rect 55634 23102 55636 23154
rect 55580 23100 55636 23102
rect 56252 29426 56308 29428
rect 56252 29374 56254 29426
rect 56254 29374 56306 29426
rect 56306 29374 56308 29426
rect 56252 29372 56308 29374
rect 59836 36204 59892 36260
rect 60060 36316 60116 36372
rect 59172 36090 59228 36092
rect 59172 36038 59174 36090
rect 59174 36038 59226 36090
rect 59226 36038 59228 36090
rect 59172 36036 59228 36038
rect 59276 36090 59332 36092
rect 59276 36038 59278 36090
rect 59278 36038 59330 36090
rect 59330 36038 59332 36090
rect 59276 36036 59332 36038
rect 59380 36090 59436 36092
rect 59380 36038 59382 36090
rect 59382 36038 59434 36090
rect 59434 36038 59436 36090
rect 59380 36036 59436 36038
rect 60508 36258 60564 36260
rect 60508 36206 60510 36258
rect 60510 36206 60562 36258
rect 60562 36206 60564 36258
rect 60508 36204 60564 36206
rect 58940 35586 58996 35588
rect 58940 35534 58942 35586
rect 58942 35534 58994 35586
rect 58994 35534 58996 35586
rect 58940 35532 58996 35534
rect 58268 35420 58324 35476
rect 57708 34860 57764 34916
rect 57596 34748 57652 34804
rect 57484 34018 57540 34020
rect 57484 33966 57486 34018
rect 57486 33966 57538 34018
rect 57538 33966 57540 34018
rect 57484 33964 57540 33966
rect 59164 35196 59220 35252
rect 59052 34914 59108 34916
rect 59052 34862 59054 34914
rect 59054 34862 59106 34914
rect 59106 34862 59108 34914
rect 59052 34860 59108 34862
rect 59612 35474 59668 35476
rect 59612 35422 59614 35474
rect 59614 35422 59666 35474
rect 59666 35422 59668 35474
rect 59612 35420 59668 35422
rect 59388 34636 59444 34692
rect 59172 34522 59228 34524
rect 59172 34470 59174 34522
rect 59174 34470 59226 34522
rect 59226 34470 59228 34522
rect 59172 34468 59228 34470
rect 59276 34522 59332 34524
rect 59276 34470 59278 34522
rect 59278 34470 59330 34522
rect 59330 34470 59332 34522
rect 59276 34468 59332 34470
rect 59380 34522 59436 34524
rect 59380 34470 59382 34522
rect 59382 34470 59434 34522
rect 59434 34470 59436 34522
rect 59380 34468 59436 34470
rect 57932 34188 57988 34244
rect 57596 33740 57652 33796
rect 59388 34242 59444 34244
rect 59388 34190 59390 34242
rect 59390 34190 59442 34242
rect 59442 34190 59444 34242
rect 59388 34188 59444 34190
rect 57820 33852 57876 33908
rect 57484 33292 57540 33348
rect 57708 33346 57764 33348
rect 57708 33294 57710 33346
rect 57710 33294 57762 33346
rect 57762 33294 57764 33346
rect 57708 33292 57764 33294
rect 58156 32620 58212 32676
rect 57596 31948 57652 32004
rect 59172 32954 59228 32956
rect 59172 32902 59174 32954
rect 59174 32902 59226 32954
rect 59226 32902 59228 32954
rect 59172 32900 59228 32902
rect 59276 32954 59332 32956
rect 59276 32902 59278 32954
rect 59278 32902 59330 32954
rect 59330 32902 59332 32954
rect 59276 32900 59332 32902
rect 59380 32954 59436 32956
rect 59380 32902 59382 32954
rect 59382 32902 59434 32954
rect 59434 32902 59436 32954
rect 59380 32900 59436 32902
rect 59276 32674 59332 32676
rect 59276 32622 59278 32674
rect 59278 32622 59330 32674
rect 59330 32622 59332 32674
rect 59276 32620 59332 32622
rect 59164 32002 59220 32004
rect 59164 31950 59166 32002
rect 59166 31950 59218 32002
rect 59218 31950 59220 32002
rect 59164 31948 59220 31950
rect 60732 35644 60788 35700
rect 60284 35196 60340 35252
rect 60620 35308 60676 35364
rect 60508 34130 60564 34132
rect 60508 34078 60510 34130
rect 60510 34078 60562 34130
rect 60562 34078 60564 34130
rect 60508 34076 60564 34078
rect 60732 34412 60788 34468
rect 59500 31948 59556 32004
rect 59836 32620 59892 32676
rect 58492 31724 58548 31780
rect 58268 31554 58324 31556
rect 58268 31502 58270 31554
rect 58270 31502 58322 31554
rect 58322 31502 58324 31554
rect 58268 31500 58324 31502
rect 57708 31388 57764 31444
rect 58716 31500 58772 31556
rect 57148 30156 57204 30212
rect 56700 29986 56756 29988
rect 56700 29934 56702 29986
rect 56702 29934 56754 29986
rect 56754 29934 56756 29986
rect 56700 29932 56756 29934
rect 56588 29314 56644 29316
rect 56588 29262 56590 29314
rect 56590 29262 56642 29314
rect 56642 29262 56644 29314
rect 56588 29260 56644 29262
rect 56700 28588 56756 28644
rect 56812 29372 56868 29428
rect 56588 27970 56644 27972
rect 56588 27918 56590 27970
rect 56590 27918 56642 27970
rect 56642 27918 56644 27970
rect 56588 27916 56644 27918
rect 57036 27916 57092 27972
rect 56476 27298 56532 27300
rect 56476 27246 56478 27298
rect 56478 27246 56530 27298
rect 56530 27246 56532 27298
rect 56476 27244 56532 27246
rect 56364 25676 56420 25732
rect 57372 29372 57428 29428
rect 58044 29820 58100 29876
rect 59500 31778 59556 31780
rect 59500 31726 59502 31778
rect 59502 31726 59554 31778
rect 59554 31726 59556 31778
rect 59500 31724 59556 31726
rect 59724 31666 59780 31668
rect 59724 31614 59726 31666
rect 59726 31614 59778 31666
rect 59778 31614 59780 31666
rect 59724 31612 59780 31614
rect 59172 31386 59228 31388
rect 59172 31334 59174 31386
rect 59174 31334 59226 31386
rect 59226 31334 59228 31386
rect 59172 31332 59228 31334
rect 59276 31386 59332 31388
rect 59276 31334 59278 31386
rect 59278 31334 59330 31386
rect 59330 31334 59332 31386
rect 59276 31332 59332 31334
rect 59380 31386 59436 31388
rect 59380 31334 59382 31386
rect 59382 31334 59434 31386
rect 59434 31334 59436 31386
rect 59380 31332 59436 31334
rect 59724 30604 59780 30660
rect 58940 30044 58996 30100
rect 59172 29818 59228 29820
rect 59172 29766 59174 29818
rect 59174 29766 59226 29818
rect 59226 29766 59228 29818
rect 59172 29764 59228 29766
rect 59276 29818 59332 29820
rect 59276 29766 59278 29818
rect 59278 29766 59330 29818
rect 59330 29766 59332 29818
rect 59276 29764 59332 29766
rect 59380 29818 59436 29820
rect 59380 29766 59382 29818
rect 59382 29766 59434 29818
rect 59434 29766 59436 29818
rect 59380 29764 59436 29766
rect 60060 32562 60116 32564
rect 60060 32510 60062 32562
rect 60062 32510 60114 32562
rect 60114 32510 60116 32562
rect 60060 32508 60116 32510
rect 60284 31948 60340 32004
rect 60620 33122 60676 33124
rect 60620 33070 60622 33122
rect 60622 33070 60674 33122
rect 60674 33070 60676 33122
rect 60620 33068 60676 33070
rect 60508 32508 60564 32564
rect 60284 31778 60340 31780
rect 60284 31726 60286 31778
rect 60286 31726 60338 31778
rect 60338 31726 60340 31778
rect 60284 31724 60340 31726
rect 60396 31666 60452 31668
rect 60396 31614 60398 31666
rect 60398 31614 60450 31666
rect 60450 31614 60452 31666
rect 60396 31612 60452 31614
rect 62860 36370 62916 36372
rect 62860 36318 62862 36370
rect 62862 36318 62914 36370
rect 62914 36318 62916 36370
rect 62860 36316 62916 36318
rect 63308 36540 63364 36596
rect 64652 36594 64708 36596
rect 64652 36542 64654 36594
rect 64654 36542 64706 36594
rect 64706 36542 64708 36594
rect 64652 36540 64708 36542
rect 68460 37884 68516 37940
rect 67452 37100 67508 37156
rect 63196 36370 63252 36372
rect 63196 36318 63198 36370
rect 63198 36318 63250 36370
rect 63250 36318 63252 36370
rect 63196 36316 63252 36318
rect 61404 35698 61460 35700
rect 61404 35646 61406 35698
rect 61406 35646 61458 35698
rect 61458 35646 61460 35698
rect 61404 35644 61460 35646
rect 61852 35532 61908 35588
rect 62860 35586 62916 35588
rect 62860 35534 62862 35586
rect 62862 35534 62914 35586
rect 62914 35534 62916 35586
rect 62860 35532 62916 35534
rect 62300 35196 62356 35252
rect 62524 35308 62580 35364
rect 62972 35308 63028 35364
rect 61292 34412 61348 34468
rect 61516 34188 61572 34244
rect 62524 33740 62580 33796
rect 64204 34860 64260 34916
rect 65884 36204 65940 36260
rect 63196 34802 63252 34804
rect 63196 34750 63198 34802
rect 63198 34750 63250 34802
rect 63250 34750 63252 34802
rect 63196 34748 63252 34750
rect 63980 34802 64036 34804
rect 63980 34750 63982 34802
rect 63982 34750 64034 34802
rect 64034 34750 64036 34802
rect 63980 34748 64036 34750
rect 64764 35698 64820 35700
rect 64764 35646 64766 35698
rect 64766 35646 64818 35698
rect 64818 35646 64820 35698
rect 64764 35644 64820 35646
rect 65548 35644 65604 35700
rect 64540 35586 64596 35588
rect 64540 35534 64542 35586
rect 64542 35534 64594 35586
rect 64594 35534 64596 35586
rect 64540 35532 64596 35534
rect 64988 35196 65044 35252
rect 64428 34748 64484 34804
rect 64988 34914 65044 34916
rect 64988 34862 64990 34914
rect 64990 34862 65042 34914
rect 65042 34862 65044 34914
rect 64988 34860 65044 34862
rect 64092 34690 64148 34692
rect 64092 34638 64094 34690
rect 64094 34638 64146 34690
rect 64146 34638 64148 34690
rect 64092 34636 64148 34638
rect 64764 34524 64820 34580
rect 64092 34300 64148 34356
rect 63084 34130 63140 34132
rect 63084 34078 63086 34130
rect 63086 34078 63138 34130
rect 63138 34078 63140 34130
rect 63084 34076 63140 34078
rect 63868 34188 63924 34244
rect 61516 33122 61572 33124
rect 61516 33070 61518 33122
rect 61518 33070 61570 33122
rect 61570 33070 61572 33122
rect 61516 33068 61572 33070
rect 63868 33404 63924 33460
rect 65324 34914 65380 34916
rect 65324 34862 65326 34914
rect 65326 34862 65378 34914
rect 65378 34862 65380 34914
rect 65324 34860 65380 34862
rect 65772 35586 65828 35588
rect 65772 35534 65774 35586
rect 65774 35534 65826 35586
rect 65826 35534 65828 35586
rect 65772 35532 65828 35534
rect 65660 35196 65716 35252
rect 64988 34300 65044 34356
rect 65660 34636 65716 34692
rect 65772 34354 65828 34356
rect 65772 34302 65774 34354
rect 65774 34302 65826 34354
rect 65826 34302 65828 34354
rect 65772 34300 65828 34302
rect 65100 34076 65156 34132
rect 64092 33404 64148 33460
rect 64204 33346 64260 33348
rect 64204 33294 64206 33346
rect 64206 33294 64258 33346
rect 64258 33294 64260 33346
rect 64204 33292 64260 33294
rect 65436 33346 65492 33348
rect 65436 33294 65438 33346
rect 65438 33294 65490 33346
rect 65490 33294 65492 33346
rect 65436 33292 65492 33294
rect 63196 33180 63252 33236
rect 60172 30604 60228 30660
rect 60732 30492 60788 30548
rect 60844 30044 60900 30100
rect 59836 29596 59892 29652
rect 58604 29426 58660 29428
rect 58604 29374 58606 29426
rect 58606 29374 58658 29426
rect 58658 29374 58660 29426
rect 58604 29372 58660 29374
rect 59500 29426 59556 29428
rect 59500 29374 59502 29426
rect 59502 29374 59554 29426
rect 59554 29374 59556 29426
rect 59500 29372 59556 29374
rect 58156 29314 58212 29316
rect 58156 29262 58158 29314
rect 58158 29262 58210 29314
rect 58210 29262 58212 29314
rect 58156 29260 58212 29262
rect 60620 29484 60676 29540
rect 60732 29650 60788 29652
rect 60732 29598 60734 29650
rect 60734 29598 60786 29650
rect 60786 29598 60788 29650
rect 60732 29596 60788 29598
rect 59724 29260 59780 29316
rect 60284 29314 60340 29316
rect 60284 29262 60286 29314
rect 60286 29262 60338 29314
rect 60338 29262 60340 29314
rect 60284 29260 60340 29262
rect 58268 28588 58324 28644
rect 57036 27244 57092 27300
rect 57372 27804 57428 27860
rect 58268 27804 58324 27860
rect 58940 28476 58996 28532
rect 59724 28476 59780 28532
rect 59500 28364 59556 28420
rect 59172 28250 59228 28252
rect 59172 28198 59174 28250
rect 59174 28198 59226 28250
rect 59226 28198 59228 28250
rect 59172 28196 59228 28198
rect 59276 28250 59332 28252
rect 59276 28198 59278 28250
rect 59278 28198 59330 28250
rect 59330 28198 59332 28250
rect 59276 28196 59332 28198
rect 59380 28250 59436 28252
rect 59380 28198 59382 28250
rect 59382 28198 59434 28250
rect 59434 28198 59436 28250
rect 59380 28196 59436 28198
rect 59276 27970 59332 27972
rect 59276 27918 59278 27970
rect 59278 27918 59330 27970
rect 59330 27918 59332 27970
rect 59276 27916 59332 27918
rect 58044 27692 58100 27748
rect 57372 27244 57428 27300
rect 56700 26796 56756 26852
rect 56476 25340 56532 25396
rect 56140 23436 56196 23492
rect 55916 22652 55972 22708
rect 53452 22258 53508 22260
rect 53452 22206 53454 22258
rect 53454 22206 53506 22258
rect 53506 22206 53508 22258
rect 53452 22204 53508 22206
rect 52444 22146 52500 22148
rect 52444 22094 52446 22146
rect 52446 22094 52498 22146
rect 52498 22094 52500 22146
rect 52444 22092 52500 22094
rect 52332 21644 52388 21700
rect 52444 21868 52500 21924
rect 52332 19740 52388 19796
rect 52332 18620 52388 18676
rect 55468 22146 55524 22148
rect 55468 22094 55470 22146
rect 55470 22094 55522 22146
rect 55522 22094 55524 22146
rect 55468 22092 55524 22094
rect 58492 27634 58548 27636
rect 58492 27582 58494 27634
rect 58494 27582 58546 27634
rect 58546 27582 58548 27634
rect 58492 27580 58548 27582
rect 57708 27020 57764 27076
rect 57148 25730 57204 25732
rect 57148 25678 57150 25730
rect 57150 25678 57202 25730
rect 57202 25678 57204 25730
rect 57148 25676 57204 25678
rect 57148 25452 57204 25508
rect 57036 25394 57092 25396
rect 57036 25342 57038 25394
rect 57038 25342 57090 25394
rect 57090 25342 57092 25394
rect 57036 25340 57092 25342
rect 56700 23436 56756 23492
rect 56812 23938 56868 23940
rect 56812 23886 56814 23938
rect 56814 23886 56866 23938
rect 56866 23886 56868 23938
rect 56812 23884 56868 23886
rect 56700 23154 56756 23156
rect 56700 23102 56702 23154
rect 56702 23102 56754 23154
rect 56754 23102 56756 23154
rect 56700 23100 56756 23102
rect 56476 22652 56532 22708
rect 58828 27804 58884 27860
rect 60172 28364 60228 28420
rect 60284 27916 60340 27972
rect 60620 27916 60676 27972
rect 59724 27804 59780 27860
rect 59052 27634 59108 27636
rect 59052 27582 59054 27634
rect 59054 27582 59106 27634
rect 59106 27582 59108 27634
rect 59052 27580 59108 27582
rect 59164 26962 59220 26964
rect 59164 26910 59166 26962
rect 59166 26910 59218 26962
rect 59218 26910 59220 26962
rect 59164 26908 59220 26910
rect 57932 26796 57988 26852
rect 59500 26796 59556 26852
rect 59172 26682 59228 26684
rect 59172 26630 59174 26682
rect 59174 26630 59226 26682
rect 59226 26630 59228 26682
rect 59172 26628 59228 26630
rect 59276 26682 59332 26684
rect 59276 26630 59278 26682
rect 59278 26630 59330 26682
rect 59330 26630 59332 26682
rect 59276 26628 59332 26630
rect 59380 26682 59436 26684
rect 59380 26630 59382 26682
rect 59382 26630 59434 26682
rect 59434 26630 59436 26682
rect 59380 26628 59436 26630
rect 57708 26290 57764 26292
rect 57708 26238 57710 26290
rect 57710 26238 57762 26290
rect 57762 26238 57764 26290
rect 57708 26236 57764 26238
rect 59052 26236 59108 26292
rect 57484 25340 57540 25396
rect 57708 25676 57764 25732
rect 58380 25618 58436 25620
rect 58380 25566 58382 25618
rect 58382 25566 58434 25618
rect 58434 25566 58436 25618
rect 58380 25564 58436 25566
rect 57596 23884 57652 23940
rect 58604 25452 58660 25508
rect 59052 25506 59108 25508
rect 59052 25454 59054 25506
rect 59054 25454 59106 25506
rect 59106 25454 59108 25506
rect 59052 25452 59108 25454
rect 58940 25340 58996 25396
rect 57484 23154 57540 23156
rect 57484 23102 57486 23154
rect 57486 23102 57538 23154
rect 57538 23102 57540 23154
rect 57484 23100 57540 23102
rect 57596 22930 57652 22932
rect 57596 22878 57598 22930
rect 57598 22878 57650 22930
rect 57650 22878 57652 22930
rect 57596 22876 57652 22878
rect 56476 22146 56532 22148
rect 56476 22094 56478 22146
rect 56478 22094 56530 22146
rect 56530 22094 56532 22146
rect 56476 22092 56532 22094
rect 53564 20524 53620 20580
rect 53788 21474 53844 21476
rect 53788 21422 53790 21474
rect 53790 21422 53842 21474
rect 53842 21422 53844 21474
rect 53788 21420 53844 21422
rect 55916 21586 55972 21588
rect 55916 21534 55918 21586
rect 55918 21534 55970 21586
rect 55970 21534 55972 21586
rect 55916 21532 55972 21534
rect 54236 21420 54292 21476
rect 55020 21420 55076 21476
rect 55020 20972 55076 21028
rect 54348 20802 54404 20804
rect 54348 20750 54350 20802
rect 54350 20750 54402 20802
rect 54402 20750 54404 20802
rect 54348 20748 54404 20750
rect 54348 20524 54404 20580
rect 53564 20018 53620 20020
rect 53564 19966 53566 20018
rect 53566 19966 53618 20018
rect 53618 19966 53620 20018
rect 53564 19964 53620 19966
rect 53228 19516 53284 19572
rect 53788 19404 53844 19460
rect 52444 18732 52500 18788
rect 55468 20524 55524 20580
rect 55804 21026 55860 21028
rect 55804 20974 55806 21026
rect 55806 20974 55858 21026
rect 55858 20974 55860 21026
rect 55804 20972 55860 20974
rect 56140 20914 56196 20916
rect 56140 20862 56142 20914
rect 56142 20862 56194 20914
rect 56194 20862 56196 20914
rect 56140 20860 56196 20862
rect 55580 20802 55636 20804
rect 55580 20750 55582 20802
rect 55582 20750 55634 20802
rect 55634 20750 55636 20802
rect 55580 20748 55636 20750
rect 54460 20018 54516 20020
rect 54460 19966 54462 20018
rect 54462 19966 54514 20018
rect 54514 19966 54516 20018
rect 54460 19964 54516 19966
rect 55916 20636 55972 20692
rect 56364 20690 56420 20692
rect 56364 20638 56366 20690
rect 56366 20638 56418 20690
rect 56418 20638 56420 20690
rect 56364 20636 56420 20638
rect 56140 20524 56196 20580
rect 55804 20018 55860 20020
rect 55804 19966 55806 20018
rect 55806 19966 55858 20018
rect 55858 19966 55860 20018
rect 55804 19964 55860 19966
rect 56588 19346 56644 19348
rect 56588 19294 56590 19346
rect 56590 19294 56642 19346
rect 56642 19294 56644 19346
rect 56588 19292 56644 19294
rect 55356 18674 55412 18676
rect 55356 18622 55358 18674
rect 55358 18622 55410 18674
rect 55410 18622 55412 18674
rect 55356 18620 55412 18622
rect 56252 18620 56308 18676
rect 53788 18450 53844 18452
rect 53788 18398 53790 18450
rect 53790 18398 53842 18450
rect 53842 18398 53844 18450
rect 53788 18396 53844 18398
rect 54796 18450 54852 18452
rect 54796 18398 54798 18450
rect 54798 18398 54850 18450
rect 54850 18398 54852 18450
rect 54796 18396 54852 18398
rect 54124 18338 54180 18340
rect 54124 18286 54126 18338
rect 54126 18286 54178 18338
rect 54178 18286 54180 18338
rect 54124 18284 54180 18286
rect 55020 18338 55076 18340
rect 55020 18286 55022 18338
rect 55022 18286 55074 18338
rect 55074 18286 55076 18338
rect 55020 18284 55076 18286
rect 55468 18284 55524 18340
rect 53340 17778 53396 17780
rect 53340 17726 53342 17778
rect 53342 17726 53394 17778
rect 53394 17726 53396 17778
rect 53340 17724 53396 17726
rect 52220 17442 52276 17444
rect 52220 17390 52222 17442
rect 52222 17390 52274 17442
rect 52274 17390 52276 17442
rect 52220 17388 52276 17390
rect 53676 17500 53732 17556
rect 52892 17106 52948 17108
rect 52892 17054 52894 17106
rect 52894 17054 52946 17106
rect 52946 17054 52948 17106
rect 52892 17052 52948 17054
rect 54460 17164 54516 17220
rect 53676 16828 53732 16884
rect 54236 16882 54292 16884
rect 54236 16830 54238 16882
rect 54238 16830 54290 16882
rect 54290 16830 54292 16882
rect 54236 16828 54292 16830
rect 52668 16770 52724 16772
rect 52668 16718 52670 16770
rect 52670 16718 52722 16770
rect 52722 16718 52724 16770
rect 52668 16716 52724 16718
rect 55020 17164 55076 17220
rect 55020 16940 55076 16996
rect 52332 16268 52388 16324
rect 54236 16268 54292 16324
rect 53116 16044 53172 16100
rect 52780 15820 52836 15876
rect 52444 15260 52500 15316
rect 53116 15314 53172 15316
rect 53116 15262 53118 15314
rect 53118 15262 53170 15314
rect 53170 15262 53172 15314
rect 53116 15260 53172 15262
rect 54124 15314 54180 15316
rect 54124 15262 54126 15314
rect 54126 15262 54178 15314
rect 54178 15262 54180 15314
rect 54124 15260 54180 15262
rect 52444 14588 52500 14644
rect 54572 16098 54628 16100
rect 54572 16046 54574 16098
rect 54574 16046 54626 16098
rect 54626 16046 54628 16098
rect 54572 16044 54628 16046
rect 55132 16828 55188 16884
rect 54796 15932 54852 15988
rect 54796 15260 54852 15316
rect 53116 14476 53172 14532
rect 54908 14530 54964 14532
rect 54908 14478 54910 14530
rect 54910 14478 54962 14530
rect 54962 14478 54964 14530
rect 54908 14476 54964 14478
rect 53116 13468 53172 13524
rect 52668 12460 52724 12516
rect 54012 13468 54068 13524
rect 53788 12962 53844 12964
rect 53788 12910 53790 12962
rect 53790 12910 53842 12962
rect 53842 12910 53844 12962
rect 53788 12908 53844 12910
rect 53676 12684 53732 12740
rect 53564 12290 53620 12292
rect 53564 12238 53566 12290
rect 53566 12238 53618 12290
rect 53618 12238 53620 12290
rect 53564 12236 53620 12238
rect 52220 11116 52276 11172
rect 52780 10892 52836 10948
rect 52444 10668 52500 10724
rect 52108 9772 52164 9828
rect 53788 12460 53844 12516
rect 54348 13522 54404 13524
rect 54348 13470 54350 13522
rect 54350 13470 54402 13522
rect 54402 13470 54404 13522
rect 54348 13468 54404 13470
rect 54460 13244 54516 13300
rect 54460 12236 54516 12292
rect 55916 16882 55972 16884
rect 55916 16830 55918 16882
rect 55918 16830 55970 16882
rect 55970 16830 55972 16882
rect 55916 16828 55972 16830
rect 56364 16770 56420 16772
rect 56364 16718 56366 16770
rect 56366 16718 56418 16770
rect 56418 16718 56420 16770
rect 56364 16716 56420 16718
rect 56700 16716 56756 16772
rect 55580 16098 55636 16100
rect 55580 16046 55582 16098
rect 55582 16046 55634 16098
rect 55634 16046 55636 16098
rect 55580 16044 55636 16046
rect 56364 15986 56420 15988
rect 56364 15934 56366 15986
rect 56366 15934 56418 15986
rect 56418 15934 56420 15986
rect 56364 15932 56420 15934
rect 55692 15874 55748 15876
rect 55692 15822 55694 15874
rect 55694 15822 55746 15874
rect 55746 15822 55748 15874
rect 55692 15820 55748 15822
rect 56588 15372 56644 15428
rect 56924 16098 56980 16100
rect 56924 16046 56926 16098
rect 56926 16046 56978 16098
rect 56978 16046 56980 16098
rect 56924 16044 56980 16046
rect 57484 22258 57540 22260
rect 57484 22206 57486 22258
rect 57486 22206 57538 22258
rect 57538 22206 57540 22258
rect 57484 22204 57540 22206
rect 57596 21868 57652 21924
rect 58492 24892 58548 24948
rect 58380 23938 58436 23940
rect 58380 23886 58382 23938
rect 58382 23886 58434 23938
rect 58434 23886 58436 23938
rect 58380 23884 58436 23886
rect 59164 25228 59220 25284
rect 59172 25114 59228 25116
rect 59172 25062 59174 25114
rect 59174 25062 59226 25114
rect 59226 25062 59228 25114
rect 59172 25060 59228 25062
rect 59276 25114 59332 25116
rect 59276 25062 59278 25114
rect 59278 25062 59330 25114
rect 59330 25062 59332 25114
rect 59276 25060 59332 25062
rect 59380 25114 59436 25116
rect 59380 25062 59382 25114
rect 59382 25062 59434 25114
rect 59434 25062 59436 25114
rect 59380 25060 59436 25062
rect 59052 24946 59108 24948
rect 59052 24894 59054 24946
rect 59054 24894 59106 24946
rect 59106 24894 59108 24946
rect 59052 24892 59108 24894
rect 59276 24834 59332 24836
rect 59276 24782 59278 24834
rect 59278 24782 59330 24834
rect 59330 24782 59332 24834
rect 59276 24780 59332 24782
rect 59052 23826 59108 23828
rect 59052 23774 59054 23826
rect 59054 23774 59106 23826
rect 59106 23774 59108 23826
rect 60396 27858 60452 27860
rect 60396 27806 60398 27858
rect 60398 27806 60450 27858
rect 60450 27806 60452 27858
rect 60396 27804 60452 27806
rect 59836 27746 59892 27748
rect 59836 27694 59838 27746
rect 59838 27694 59890 27746
rect 59890 27694 59892 27746
rect 59836 27692 59892 27694
rect 60060 26402 60116 26404
rect 60060 26350 60062 26402
rect 60062 26350 60114 26402
rect 60114 26350 60116 26402
rect 60060 26348 60116 26350
rect 59948 25452 60004 25508
rect 60396 25340 60452 25396
rect 60060 24780 60116 24836
rect 59724 23826 59780 23828
rect 59052 23772 59108 23774
rect 58268 23660 58324 23716
rect 59724 23774 59726 23826
rect 59726 23774 59778 23826
rect 59778 23774 59780 23826
rect 59724 23772 59780 23774
rect 59276 23714 59332 23716
rect 59276 23662 59278 23714
rect 59278 23662 59330 23714
rect 59330 23662 59332 23714
rect 59276 23660 59332 23662
rect 59172 23546 59228 23548
rect 59172 23494 59174 23546
rect 59174 23494 59226 23546
rect 59226 23494 59228 23546
rect 59172 23492 59228 23494
rect 59276 23546 59332 23548
rect 59276 23494 59278 23546
rect 59278 23494 59330 23546
rect 59330 23494 59332 23546
rect 59276 23492 59332 23494
rect 59380 23546 59436 23548
rect 59380 23494 59382 23546
rect 59382 23494 59434 23546
rect 59434 23494 59436 23546
rect 59380 23492 59436 23494
rect 58044 22876 58100 22932
rect 58156 23100 58212 23156
rect 58380 22428 58436 22484
rect 58156 21868 58212 21924
rect 58268 22092 58324 22148
rect 58604 22258 58660 22260
rect 58604 22206 58606 22258
rect 58606 22206 58658 22258
rect 58658 22206 58660 22258
rect 58604 22204 58660 22206
rect 58940 23042 58996 23044
rect 58940 22990 58942 23042
rect 58942 22990 58994 23042
rect 58994 22990 58996 23042
rect 58940 22988 58996 22990
rect 59836 23714 59892 23716
rect 59836 23662 59838 23714
rect 59838 23662 59890 23714
rect 59890 23662 59892 23714
rect 59836 23660 59892 23662
rect 59500 22988 59556 23044
rect 59164 22428 59220 22484
rect 58716 22092 58772 22148
rect 58380 21980 58436 22036
rect 59388 22146 59444 22148
rect 59388 22094 59390 22146
rect 59390 22094 59442 22146
rect 59442 22094 59444 22146
rect 59388 22092 59444 22094
rect 60732 25676 60788 25732
rect 60844 25228 60900 25284
rect 60284 23660 60340 23716
rect 60396 23772 60452 23828
rect 60060 23324 60116 23380
rect 60060 23154 60116 23156
rect 60060 23102 60062 23154
rect 60062 23102 60114 23154
rect 60114 23102 60116 23154
rect 60060 23100 60116 23102
rect 59948 22876 60004 22932
rect 59836 22482 59892 22484
rect 59836 22430 59838 22482
rect 59838 22430 59890 22482
rect 59890 22430 59892 22482
rect 59836 22428 59892 22430
rect 59724 22092 59780 22148
rect 59948 22204 60004 22260
rect 59172 21978 59228 21980
rect 59172 21926 59174 21978
rect 59174 21926 59226 21978
rect 59226 21926 59228 21978
rect 59172 21924 59228 21926
rect 59276 21978 59332 21980
rect 59276 21926 59278 21978
rect 59278 21926 59330 21978
rect 59330 21926 59332 21978
rect 59276 21924 59332 21926
rect 59380 21978 59436 21980
rect 59380 21926 59382 21978
rect 59382 21926 59434 21978
rect 59434 21926 59436 21978
rect 59380 21924 59436 21926
rect 59052 21756 59108 21812
rect 59500 21810 59556 21812
rect 59500 21758 59502 21810
rect 59502 21758 59554 21810
rect 59554 21758 59556 21810
rect 59500 21756 59556 21758
rect 59164 21644 59220 21700
rect 57820 19346 57876 19348
rect 57820 19294 57822 19346
rect 57822 19294 57874 19346
rect 57874 19294 57876 19346
rect 57820 19292 57876 19294
rect 57484 16882 57540 16884
rect 57484 16830 57486 16882
rect 57486 16830 57538 16882
rect 57538 16830 57540 16882
rect 57484 16828 57540 16830
rect 57708 16770 57764 16772
rect 57708 16718 57710 16770
rect 57710 16718 57762 16770
rect 57762 16718 57764 16770
rect 57708 16716 57764 16718
rect 57484 16044 57540 16100
rect 57372 15932 57428 15988
rect 57820 15986 57876 15988
rect 57820 15934 57822 15986
rect 57822 15934 57874 15986
rect 57874 15934 57876 15986
rect 57820 15932 57876 15934
rect 57596 15874 57652 15876
rect 57596 15822 57598 15874
rect 57598 15822 57650 15874
rect 57650 15822 57652 15874
rect 57596 15820 57652 15822
rect 57036 14642 57092 14644
rect 57036 14590 57038 14642
rect 57038 14590 57090 14642
rect 57090 14590 57092 14642
rect 57036 14588 57092 14590
rect 55356 13244 55412 13300
rect 56924 13356 56980 13412
rect 55916 13132 55972 13188
rect 55132 12962 55188 12964
rect 55132 12910 55134 12962
rect 55134 12910 55186 12962
rect 55186 12910 55188 12962
rect 55132 12908 55188 12910
rect 56140 12962 56196 12964
rect 56140 12910 56142 12962
rect 56142 12910 56194 12962
rect 56194 12910 56196 12962
rect 56140 12908 56196 12910
rect 57148 13020 57204 13076
rect 55916 12402 55972 12404
rect 55916 12350 55918 12402
rect 55918 12350 55970 12402
rect 55970 12350 55972 12402
rect 55916 12348 55972 12350
rect 55244 12290 55300 12292
rect 55244 12238 55246 12290
rect 55246 12238 55298 12290
rect 55298 12238 55300 12290
rect 56588 12402 56644 12404
rect 56588 12350 56590 12402
rect 56590 12350 56642 12402
rect 56642 12350 56644 12402
rect 56588 12348 56644 12350
rect 55244 12236 55300 12238
rect 56476 12012 56532 12068
rect 54236 11506 54292 11508
rect 54236 11454 54238 11506
rect 54238 11454 54290 11506
rect 54290 11454 54292 11506
rect 54236 11452 54292 11454
rect 53228 10722 53284 10724
rect 53228 10670 53230 10722
rect 53230 10670 53282 10722
rect 53282 10670 53284 10722
rect 53228 10668 53284 10670
rect 56364 11506 56420 11508
rect 56364 11454 56366 11506
rect 56366 11454 56418 11506
rect 56418 11454 56420 11506
rect 56364 11452 56420 11454
rect 56924 12012 56980 12068
rect 57372 12572 57428 12628
rect 57260 11506 57316 11508
rect 57260 11454 57262 11506
rect 57262 11454 57314 11506
rect 57314 11454 57316 11506
rect 57260 11452 57316 11454
rect 57036 11394 57092 11396
rect 57036 11342 57038 11394
rect 57038 11342 57090 11394
rect 57090 11342 57092 11394
rect 57036 11340 57092 11342
rect 54236 10556 54292 10612
rect 55804 10834 55860 10836
rect 55804 10782 55806 10834
rect 55806 10782 55858 10834
rect 55858 10782 55860 10834
rect 55804 10780 55860 10782
rect 56476 10834 56532 10836
rect 56476 10782 56478 10834
rect 56478 10782 56530 10834
rect 56530 10782 56532 10834
rect 56476 10780 56532 10782
rect 54796 10610 54852 10612
rect 54796 10558 54798 10610
rect 54798 10558 54850 10610
rect 54850 10558 54852 10610
rect 54796 10556 54852 10558
rect 56588 10610 56644 10612
rect 56588 10558 56590 10610
rect 56590 10558 56642 10610
rect 56642 10558 56644 10610
rect 56588 10556 56644 10558
rect 56700 10498 56756 10500
rect 56700 10446 56702 10498
rect 56702 10446 56754 10498
rect 56754 10446 56756 10498
rect 56700 10444 56756 10446
rect 60844 24556 60900 24612
rect 60732 23772 60788 23828
rect 60844 23660 60900 23716
rect 60620 23324 60676 23380
rect 60620 22482 60676 22484
rect 60620 22430 60622 22482
rect 60622 22430 60674 22482
rect 60674 22430 60676 22482
rect 60620 22428 60676 22430
rect 60396 22316 60452 22372
rect 58716 20914 58772 20916
rect 58716 20862 58718 20914
rect 58718 20862 58770 20914
rect 58770 20862 58772 20914
rect 58716 20860 58772 20862
rect 59612 20860 59668 20916
rect 58604 20802 58660 20804
rect 58604 20750 58606 20802
rect 58606 20750 58658 20802
rect 58658 20750 58660 20802
rect 58604 20748 58660 20750
rect 58044 19234 58100 19236
rect 58044 19182 58046 19234
rect 58046 19182 58098 19234
rect 58098 19182 58100 19234
rect 58044 19180 58100 19182
rect 58492 19180 58548 19236
rect 58156 18732 58212 18788
rect 58044 17554 58100 17556
rect 58044 17502 58046 17554
rect 58046 17502 58098 17554
rect 58098 17502 58100 17554
rect 58044 17500 58100 17502
rect 58044 17276 58100 17332
rect 58268 18620 58324 18676
rect 58604 17276 58660 17332
rect 58156 14588 58212 14644
rect 57484 12290 57540 12292
rect 57484 12238 57486 12290
rect 57486 12238 57538 12290
rect 57538 12238 57540 12290
rect 57484 12236 57540 12238
rect 57484 10610 57540 10612
rect 57484 10558 57486 10610
rect 57486 10558 57538 10610
rect 57538 10558 57540 10610
rect 57484 10556 57540 10558
rect 52780 9660 52836 9716
rect 52108 9212 52164 9268
rect 50316 8204 50372 8260
rect 50764 8258 50820 8260
rect 50764 8206 50766 8258
rect 50766 8206 50818 8258
rect 50818 8206 50820 8258
rect 50764 8204 50820 8206
rect 48188 7644 48244 7700
rect 48524 7980 48580 8036
rect 47292 7196 47348 7252
rect 46620 6748 46676 6804
rect 47404 6860 47460 6916
rect 46508 6466 46564 6468
rect 46508 6414 46510 6466
rect 46510 6414 46562 6466
rect 46562 6414 46564 6466
rect 46508 6412 46564 6414
rect 45948 6300 46004 6356
rect 46172 6130 46228 6132
rect 46172 6078 46174 6130
rect 46174 6078 46226 6130
rect 46226 6078 46228 6130
rect 46172 6076 46228 6078
rect 45724 5180 45780 5236
rect 44940 4956 44996 5012
rect 45612 5010 45668 5012
rect 45612 4958 45614 5010
rect 45614 4958 45666 5010
rect 45666 4958 45668 5010
rect 45612 4956 45668 4958
rect 44716 4732 44772 4788
rect 45388 3724 45444 3780
rect 44044 3554 44100 3556
rect 44044 3502 44046 3554
rect 44046 3502 44098 3554
rect 44098 3502 44100 3554
rect 44044 3500 44100 3502
rect 46060 5794 46116 5796
rect 46060 5742 46062 5794
rect 46062 5742 46114 5794
rect 46114 5742 46116 5794
rect 46060 5740 46116 5742
rect 45836 4844 45892 4900
rect 46508 5516 46564 5572
rect 46172 5404 46228 5460
rect 46396 5346 46452 5348
rect 46396 5294 46398 5346
rect 46398 5294 46450 5346
rect 46450 5294 46452 5346
rect 46396 5292 46452 5294
rect 46172 4508 46228 4564
rect 44940 3276 44996 3332
rect 45276 3388 45332 3444
rect 43932 1484 43988 1540
rect 46508 4620 46564 4676
rect 46284 3164 46340 3220
rect 45612 3052 45668 3108
rect 47068 6466 47124 6468
rect 47068 6414 47070 6466
rect 47070 6414 47122 6466
rect 47122 6414 47124 6466
rect 47068 6412 47124 6414
rect 46732 5964 46788 6020
rect 46844 5404 46900 5460
rect 46732 4844 46788 4900
rect 46844 4732 46900 4788
rect 47180 5516 47236 5572
rect 46956 4562 47012 4564
rect 46956 4510 46958 4562
rect 46958 4510 47010 4562
rect 47010 4510 47012 4562
rect 46956 4508 47012 4510
rect 47852 6748 47908 6804
rect 48412 7196 48468 7252
rect 48636 7644 48692 7700
rect 49196 8034 49252 8036
rect 49196 7982 49198 8034
rect 49198 7982 49250 8034
rect 49250 7982 49252 8034
rect 49196 7980 49252 7982
rect 49644 7644 49700 7700
rect 48860 7532 48916 7588
rect 49308 7532 49364 7588
rect 48524 7084 48580 7140
rect 49196 6972 49252 7028
rect 47852 6300 47908 6356
rect 47404 5404 47460 5460
rect 47516 6076 47572 6132
rect 47404 4508 47460 4564
rect 47292 4396 47348 4452
rect 48300 6076 48356 6132
rect 48860 6524 48916 6580
rect 48748 6300 48804 6356
rect 48636 6130 48692 6132
rect 48636 6078 48638 6130
rect 48638 6078 48690 6130
rect 48690 6078 48692 6130
rect 48636 6076 48692 6078
rect 48188 5794 48244 5796
rect 48188 5742 48190 5794
rect 48190 5742 48242 5794
rect 48242 5742 48244 5794
rect 48188 5740 48244 5742
rect 47628 5292 47684 5348
rect 47964 5292 48020 5348
rect 47404 3948 47460 4004
rect 48636 5516 48692 5572
rect 48412 5068 48468 5124
rect 48524 5292 48580 5348
rect 48748 4620 48804 4676
rect 47516 3276 47572 3332
rect 47628 3500 47684 3556
rect 47964 3442 48020 3444
rect 47964 3390 47966 3442
rect 47966 3390 48018 3442
rect 48018 3390 48020 3442
rect 47964 3388 48020 3390
rect 50652 7868 50708 7924
rect 50428 7532 50484 7588
rect 49512 7082 49568 7084
rect 49512 7030 49514 7082
rect 49514 7030 49566 7082
rect 49566 7030 49568 7082
rect 49512 7028 49568 7030
rect 49616 7082 49672 7084
rect 49616 7030 49618 7082
rect 49618 7030 49670 7082
rect 49670 7030 49672 7082
rect 49616 7028 49672 7030
rect 49720 7082 49776 7084
rect 49720 7030 49722 7082
rect 49722 7030 49774 7082
rect 49774 7030 49776 7082
rect 49720 7028 49776 7030
rect 49756 6188 49812 6244
rect 49644 6018 49700 6020
rect 49644 5966 49646 6018
rect 49646 5966 49698 6018
rect 49698 5966 49700 6018
rect 49644 5964 49700 5966
rect 50092 6914 50148 6916
rect 50092 6862 50094 6914
rect 50094 6862 50146 6914
rect 50146 6862 50148 6914
rect 50092 6860 50148 6862
rect 50876 6914 50932 6916
rect 50876 6862 50878 6914
rect 50878 6862 50930 6914
rect 50930 6862 50932 6914
rect 50876 6860 50932 6862
rect 49868 6076 49924 6132
rect 49532 5740 49588 5796
rect 49980 6578 50036 6580
rect 49980 6526 49982 6578
rect 49982 6526 50034 6578
rect 50034 6526 50036 6578
rect 49980 6524 50036 6526
rect 49980 5964 50036 6020
rect 51772 7756 51828 7812
rect 51548 7420 51604 7476
rect 51324 7250 51380 7252
rect 51324 7198 51326 7250
rect 51326 7198 51378 7250
rect 51378 7198 51380 7250
rect 51324 7196 51380 7198
rect 51212 6690 51268 6692
rect 51212 6638 51214 6690
rect 51214 6638 51266 6690
rect 51266 6638 51268 6690
rect 51212 6636 51268 6638
rect 51884 7308 51940 7364
rect 51996 6636 52052 6692
rect 51436 6578 51492 6580
rect 51436 6526 51438 6578
rect 51438 6526 51490 6578
rect 51490 6526 51492 6578
rect 51436 6524 51492 6526
rect 51100 6412 51156 6468
rect 50092 5852 50148 5908
rect 49512 5514 49568 5516
rect 49512 5462 49514 5514
rect 49514 5462 49566 5514
rect 49566 5462 49568 5514
rect 49512 5460 49568 5462
rect 49616 5514 49672 5516
rect 49616 5462 49618 5514
rect 49618 5462 49670 5514
rect 49670 5462 49672 5514
rect 49616 5460 49672 5462
rect 49720 5514 49776 5516
rect 49720 5462 49722 5514
rect 49722 5462 49774 5514
rect 49774 5462 49776 5514
rect 49720 5460 49776 5462
rect 49308 5122 49364 5124
rect 49308 5070 49310 5122
rect 49310 5070 49362 5122
rect 49362 5070 49364 5122
rect 49308 5068 49364 5070
rect 50652 5794 50708 5796
rect 50652 5742 50654 5794
rect 50654 5742 50706 5794
rect 50706 5742 50708 5794
rect 50652 5740 50708 5742
rect 50428 5234 50484 5236
rect 50428 5182 50430 5234
rect 50430 5182 50482 5234
rect 50482 5182 50484 5234
rect 50428 5180 50484 5182
rect 50204 4508 50260 4564
rect 50540 5068 50596 5124
rect 52108 6076 52164 6132
rect 51212 5740 51268 5796
rect 50988 4956 51044 5012
rect 49756 4450 49812 4452
rect 49756 4398 49758 4450
rect 49758 4398 49810 4450
rect 49810 4398 49812 4450
rect 49756 4396 49812 4398
rect 48636 3276 48692 3332
rect 48748 3164 48804 3220
rect 47180 2492 47236 2548
rect 46620 812 46676 868
rect 49512 3946 49568 3948
rect 49512 3894 49514 3946
rect 49514 3894 49566 3946
rect 49566 3894 49568 3946
rect 49512 3892 49568 3894
rect 49616 3946 49672 3948
rect 49616 3894 49618 3946
rect 49618 3894 49670 3946
rect 49670 3894 49672 3946
rect 49616 3892 49672 3894
rect 49720 3946 49776 3948
rect 49720 3894 49722 3946
rect 49722 3894 49774 3946
rect 49774 3894 49776 3946
rect 49720 3892 49776 3894
rect 50092 4284 50148 4340
rect 50764 4284 50820 4340
rect 48860 2940 48916 2996
rect 50876 3612 50932 3668
rect 50988 3500 51044 3556
rect 51436 5628 51492 5684
rect 51548 5964 51604 6020
rect 51324 5516 51380 5572
rect 51324 4732 51380 4788
rect 51996 5906 52052 5908
rect 51996 5854 51998 5906
rect 51998 5854 52050 5906
rect 52050 5854 52052 5906
rect 51996 5852 52052 5854
rect 52332 7868 52388 7924
rect 52444 7756 52500 7812
rect 52220 5628 52276 5684
rect 52332 7308 52388 7364
rect 52780 8930 52836 8932
rect 52780 8878 52782 8930
rect 52782 8878 52834 8930
rect 52834 8878 52836 8930
rect 52780 8876 52836 8878
rect 53340 7756 53396 7812
rect 52668 7308 52724 7364
rect 52332 6748 52388 6804
rect 51772 5292 51828 5348
rect 51324 4338 51380 4340
rect 51324 4286 51326 4338
rect 51326 4286 51378 4338
rect 51378 4286 51380 4338
rect 51324 4284 51380 4286
rect 51660 4620 51716 4676
rect 52108 4284 52164 4340
rect 52556 6690 52612 6692
rect 52556 6638 52558 6690
rect 52558 6638 52610 6690
rect 52610 6638 52612 6690
rect 52556 6636 52612 6638
rect 52444 6188 52500 6244
rect 52444 4620 52500 4676
rect 51548 4172 51604 4228
rect 51324 3052 51380 3108
rect 51660 3500 51716 3556
rect 51212 1148 51268 1204
rect 54460 9548 54516 9604
rect 54348 9324 54404 9380
rect 53788 7308 53844 7364
rect 54236 8092 54292 8148
rect 53004 6972 53060 7028
rect 52892 6860 52948 6916
rect 52780 6636 52836 6692
rect 52892 5628 52948 5684
rect 53004 4620 53060 4676
rect 53676 6972 53732 7028
rect 54348 6860 54404 6916
rect 53564 6412 53620 6468
rect 53340 6130 53396 6132
rect 53340 6078 53342 6130
rect 53342 6078 53394 6130
rect 53394 6078 53396 6130
rect 53340 6076 53396 6078
rect 53228 4396 53284 4452
rect 53340 5628 53396 5684
rect 53116 4172 53172 4228
rect 53900 5964 53956 6020
rect 53564 5068 53620 5124
rect 53564 4396 53620 4452
rect 52668 3500 52724 3556
rect 51772 3442 51828 3444
rect 51772 3390 51774 3442
rect 51774 3390 51826 3442
rect 51826 3390 51828 3442
rect 51772 3388 51828 3390
rect 54796 9100 54852 9156
rect 54684 8988 54740 9044
rect 54796 8876 54852 8932
rect 54572 7474 54628 7476
rect 54572 7422 54574 7474
rect 54574 7422 54626 7474
rect 54626 7422 54628 7474
rect 54572 7420 54628 7422
rect 54684 6972 54740 7028
rect 54460 6300 54516 6356
rect 53900 5180 53956 5236
rect 54012 5516 54068 5572
rect 53788 4956 53844 5012
rect 53676 4732 53732 4788
rect 53676 4284 53732 4340
rect 53900 4620 53956 4676
rect 53564 3276 53620 3332
rect 53788 2828 53844 2884
rect 54460 5516 54516 5572
rect 54124 4226 54180 4228
rect 54124 4174 54126 4226
rect 54126 4174 54178 4226
rect 54178 4174 54180 4226
rect 54124 4172 54180 4174
rect 54012 2156 54068 2212
rect 54684 5964 54740 6020
rect 54908 5906 54964 5908
rect 54908 5854 54910 5906
rect 54910 5854 54962 5906
rect 54962 5854 54964 5906
rect 54908 5852 54964 5854
rect 54796 5740 54852 5796
rect 56140 9154 56196 9156
rect 56140 9102 56142 9154
rect 56142 9102 56194 9154
rect 56194 9102 56196 9154
rect 56140 9100 56196 9102
rect 55916 9042 55972 9044
rect 55916 8990 55918 9042
rect 55918 8990 55970 9042
rect 55970 8990 55972 9042
rect 55916 8988 55972 8990
rect 56028 8930 56084 8932
rect 56028 8878 56030 8930
rect 56030 8878 56082 8930
rect 56082 8878 56084 8930
rect 56028 8876 56084 8878
rect 55580 8370 55636 8372
rect 55580 8318 55582 8370
rect 55582 8318 55634 8370
rect 55634 8318 55636 8370
rect 55580 8316 55636 8318
rect 55132 8092 55188 8148
rect 55356 6972 55412 7028
rect 55692 7308 55748 7364
rect 55580 6690 55636 6692
rect 55580 6638 55582 6690
rect 55582 6638 55634 6690
rect 55634 6638 55636 6690
rect 55580 6636 55636 6638
rect 55468 6524 55524 6580
rect 55916 6972 55972 7028
rect 55804 6690 55860 6692
rect 55804 6638 55806 6690
rect 55806 6638 55858 6690
rect 55858 6638 55860 6690
rect 55804 6636 55860 6638
rect 56028 6690 56084 6692
rect 56028 6638 56030 6690
rect 56030 6638 56082 6690
rect 56082 6638 56084 6690
rect 56028 6636 56084 6638
rect 56028 6188 56084 6244
rect 55356 5964 55412 6020
rect 54796 5010 54852 5012
rect 54796 4958 54798 5010
rect 54798 4958 54850 5010
rect 54850 4958 54852 5010
rect 54796 4956 54852 4958
rect 54684 4898 54740 4900
rect 54684 4846 54686 4898
rect 54686 4846 54738 4898
rect 54738 4846 54740 4898
rect 54684 4844 54740 4846
rect 54796 4732 54852 4788
rect 54796 4450 54852 4452
rect 54796 4398 54798 4450
rect 54798 4398 54850 4450
rect 54850 4398 54852 4450
rect 54796 4396 54852 4398
rect 56140 6076 56196 6132
rect 56028 5964 56084 6020
rect 55468 5852 55524 5908
rect 55916 5906 55972 5908
rect 55916 5854 55918 5906
rect 55918 5854 55970 5906
rect 55970 5854 55972 5906
rect 55916 5852 55972 5854
rect 55580 5516 55636 5572
rect 56140 5628 56196 5684
rect 55468 5404 55524 5460
rect 55020 4956 55076 5012
rect 55020 4620 55076 4676
rect 55244 4396 55300 4452
rect 55020 4284 55076 4340
rect 54796 4172 54852 4228
rect 55244 4060 55300 4116
rect 55132 2828 55188 2884
rect 54348 1596 54404 1652
rect 55580 4956 55636 5012
rect 55916 4898 55972 4900
rect 55916 4846 55918 4898
rect 55918 4846 55970 4898
rect 55970 4846 55972 4898
rect 55916 4844 55972 4846
rect 56140 4508 56196 4564
rect 57372 9548 57428 9604
rect 56700 9436 56756 9492
rect 57372 9324 57428 9380
rect 56700 8316 56756 8372
rect 56476 6636 56532 6692
rect 56364 5404 56420 5460
rect 57484 8258 57540 8260
rect 57484 8206 57486 8258
rect 57486 8206 57538 8258
rect 57538 8206 57540 8258
rect 57484 8204 57540 8206
rect 57372 8034 57428 8036
rect 57372 7982 57374 8034
rect 57374 7982 57426 8034
rect 57426 7982 57428 8034
rect 57372 7980 57428 7982
rect 56812 6636 56868 6692
rect 56588 6524 56644 6580
rect 56700 6300 56756 6356
rect 57036 6076 57092 6132
rect 56588 5628 56644 5684
rect 56588 5346 56644 5348
rect 56588 5294 56590 5346
rect 56590 5294 56642 5346
rect 56642 5294 56644 5346
rect 56588 5292 56644 5294
rect 56588 5068 56644 5124
rect 56700 4620 56756 4676
rect 55580 3836 55636 3892
rect 55468 3612 55524 3668
rect 55356 1036 55412 1092
rect 57148 4956 57204 5012
rect 56812 4508 56868 4564
rect 58156 13804 58212 13860
rect 58044 13020 58100 13076
rect 58044 12572 58100 12628
rect 58492 12572 58548 12628
rect 57932 11506 57988 11508
rect 57932 11454 57934 11506
rect 57934 11454 57986 11506
rect 57986 11454 57988 11506
rect 57932 11452 57988 11454
rect 58268 11394 58324 11396
rect 58268 11342 58270 11394
rect 58270 11342 58322 11394
rect 58322 11342 58324 11394
rect 58268 11340 58324 11342
rect 57708 10834 57764 10836
rect 57708 10782 57710 10834
rect 57710 10782 57762 10834
rect 57762 10782 57764 10834
rect 57708 10780 57764 10782
rect 58380 10498 58436 10500
rect 58380 10446 58382 10498
rect 58382 10446 58434 10498
rect 58434 10446 58436 10498
rect 58380 10444 58436 10446
rect 58492 9602 58548 9604
rect 58492 9550 58494 9602
rect 58494 9550 58546 9602
rect 58546 9550 58548 9602
rect 58492 9548 58548 9550
rect 58044 9436 58100 9492
rect 58380 8258 58436 8260
rect 58380 8206 58382 8258
rect 58382 8206 58434 8258
rect 58434 8206 58436 8258
rect 58380 8204 58436 8206
rect 57932 8034 57988 8036
rect 57932 7982 57934 8034
rect 57934 7982 57986 8034
rect 57986 7982 57988 8034
rect 57932 7980 57988 7982
rect 58380 7980 58436 8036
rect 58044 7420 58100 7476
rect 57372 7362 57428 7364
rect 57372 7310 57374 7362
rect 57374 7310 57426 7362
rect 57426 7310 57428 7362
rect 57372 7308 57428 7310
rect 58380 7362 58436 7364
rect 58380 7310 58382 7362
rect 58382 7310 58434 7362
rect 58434 7310 58436 7362
rect 58380 7308 58436 7310
rect 57820 6636 57876 6692
rect 57372 6466 57428 6468
rect 57372 6414 57374 6466
rect 57374 6414 57426 6466
rect 57426 6414 57428 6466
rect 57372 6412 57428 6414
rect 57932 6300 57988 6356
rect 58044 7196 58100 7252
rect 58156 6524 58212 6580
rect 57708 6018 57764 6020
rect 57708 5966 57710 6018
rect 57710 5966 57762 6018
rect 57762 5966 57764 6018
rect 57708 5964 57764 5966
rect 57596 5740 57652 5796
rect 57596 5234 57652 5236
rect 57596 5182 57598 5234
rect 57598 5182 57650 5234
rect 57650 5182 57652 5234
rect 57596 5180 57652 5182
rect 56700 4172 56756 4228
rect 57708 4844 57764 4900
rect 56812 3330 56868 3332
rect 56812 3278 56814 3330
rect 56814 3278 56866 3330
rect 56866 3278 56868 3330
rect 56812 3276 56868 3278
rect 56588 1260 56644 1316
rect 57484 3948 57540 4004
rect 58156 5964 58212 6020
rect 58044 5740 58100 5796
rect 59172 20410 59228 20412
rect 59172 20358 59174 20410
rect 59174 20358 59226 20410
rect 59226 20358 59228 20410
rect 59172 20356 59228 20358
rect 59276 20410 59332 20412
rect 59276 20358 59278 20410
rect 59278 20358 59330 20410
rect 59330 20358 59332 20410
rect 59276 20356 59332 20358
rect 59380 20410 59436 20412
rect 59380 20358 59382 20410
rect 59382 20358 59434 20410
rect 59434 20358 59436 20410
rect 59380 20356 59436 20358
rect 59948 19964 60004 20020
rect 60060 21644 60116 21700
rect 60060 20748 60116 20804
rect 59388 19234 59444 19236
rect 59388 19182 59390 19234
rect 59390 19182 59442 19234
rect 59442 19182 59444 19234
rect 59388 19180 59444 19182
rect 59172 18842 59228 18844
rect 58940 18732 58996 18788
rect 59172 18790 59174 18842
rect 59174 18790 59226 18842
rect 59226 18790 59228 18842
rect 59172 18788 59228 18790
rect 59276 18842 59332 18844
rect 59276 18790 59278 18842
rect 59278 18790 59330 18842
rect 59330 18790 59332 18842
rect 59276 18788 59332 18790
rect 59380 18842 59436 18844
rect 59380 18790 59382 18842
rect 59382 18790 59434 18842
rect 59434 18790 59436 18842
rect 59380 18788 59436 18790
rect 59164 18620 59220 18676
rect 59388 18674 59444 18676
rect 59388 18622 59390 18674
rect 59390 18622 59442 18674
rect 59442 18622 59444 18674
rect 59388 18620 59444 18622
rect 60172 19180 60228 19236
rect 60172 18620 60228 18676
rect 60508 21420 60564 21476
rect 60396 20802 60452 20804
rect 60396 20750 60398 20802
rect 60398 20750 60450 20802
rect 60450 20750 60452 20802
rect 60396 20748 60452 20750
rect 59724 18450 59780 18452
rect 59724 18398 59726 18450
rect 59726 18398 59778 18450
rect 59778 18398 59780 18450
rect 59724 18396 59780 18398
rect 59500 17500 59556 17556
rect 59172 17274 59228 17276
rect 59172 17222 59174 17274
rect 59174 17222 59226 17274
rect 59226 17222 59228 17274
rect 59172 17220 59228 17222
rect 59276 17274 59332 17276
rect 59276 17222 59278 17274
rect 59278 17222 59330 17274
rect 59330 17222 59332 17274
rect 59276 17220 59332 17222
rect 59380 17274 59436 17276
rect 59380 17222 59382 17274
rect 59382 17222 59434 17274
rect 59434 17222 59436 17274
rect 59380 17220 59436 17222
rect 59172 15706 59228 15708
rect 59172 15654 59174 15706
rect 59174 15654 59226 15706
rect 59226 15654 59228 15706
rect 59172 15652 59228 15654
rect 59276 15706 59332 15708
rect 59276 15654 59278 15706
rect 59278 15654 59330 15706
rect 59330 15654 59332 15706
rect 59276 15652 59332 15654
rect 59380 15706 59436 15708
rect 59380 15654 59382 15706
rect 59382 15654 59434 15706
rect 59434 15654 59436 15706
rect 59380 15652 59436 15654
rect 59948 16098 60004 16100
rect 59948 16046 59950 16098
rect 59950 16046 60002 16098
rect 60002 16046 60004 16098
rect 59948 16044 60004 16046
rect 59172 14138 59228 14140
rect 59172 14086 59174 14138
rect 59174 14086 59226 14138
rect 59226 14086 59228 14138
rect 59172 14084 59228 14086
rect 59276 14138 59332 14140
rect 59276 14086 59278 14138
rect 59278 14086 59330 14138
rect 59330 14086 59332 14138
rect 59276 14084 59332 14086
rect 59380 14138 59436 14140
rect 59380 14086 59382 14138
rect 59382 14086 59434 14138
rect 59434 14086 59436 14138
rect 59380 14084 59436 14086
rect 59276 13804 59332 13860
rect 60060 13804 60116 13860
rect 59836 13468 59892 13524
rect 60732 18172 60788 18228
rect 60396 17500 60452 17556
rect 60284 17106 60340 17108
rect 60284 17054 60286 17106
rect 60286 17054 60338 17106
rect 60338 17054 60340 17106
rect 60284 17052 60340 17054
rect 60732 17106 60788 17108
rect 60732 17054 60734 17106
rect 60734 17054 60786 17106
rect 60786 17054 60788 17106
rect 60732 17052 60788 17054
rect 60396 16044 60452 16100
rect 61516 32562 61572 32564
rect 61516 32510 61518 32562
rect 61518 32510 61570 32562
rect 61570 32510 61572 32562
rect 61516 32508 61572 32510
rect 61628 32396 61684 32452
rect 62188 32562 62244 32564
rect 62188 32510 62190 32562
rect 62190 32510 62242 32562
rect 62242 32510 62244 32562
rect 62188 32508 62244 32510
rect 63196 32562 63252 32564
rect 63196 32510 63198 32562
rect 63198 32510 63250 32562
rect 63250 32510 63252 32562
rect 63196 32508 63252 32510
rect 62636 32450 62692 32452
rect 62636 32398 62638 32450
rect 62638 32398 62690 32450
rect 62690 32398 62692 32450
rect 62636 32396 62692 32398
rect 61404 28530 61460 28532
rect 61404 28478 61406 28530
rect 61406 28478 61458 28530
rect 61458 28478 61460 28530
rect 61404 28476 61460 28478
rect 61852 31778 61908 31780
rect 61852 31726 61854 31778
rect 61854 31726 61906 31778
rect 61906 31726 61908 31778
rect 61852 31724 61908 31726
rect 62300 31724 62356 31780
rect 62300 30828 62356 30884
rect 61964 30604 62020 30660
rect 62076 30210 62132 30212
rect 62076 30158 62078 30210
rect 62078 30158 62130 30210
rect 62130 30158 62132 30210
rect 62076 30156 62132 30158
rect 61628 29484 61684 29540
rect 61628 28418 61684 28420
rect 61628 28366 61630 28418
rect 61630 28366 61682 28418
rect 61682 28366 61684 28418
rect 61628 28364 61684 28366
rect 61404 27970 61460 27972
rect 61404 27918 61406 27970
rect 61406 27918 61458 27970
rect 61458 27918 61460 27970
rect 61404 27916 61460 27918
rect 61852 27804 61908 27860
rect 61292 26908 61348 26964
rect 61180 26348 61236 26404
rect 61628 26962 61684 26964
rect 61628 26910 61630 26962
rect 61630 26910 61682 26962
rect 61682 26910 61684 26962
rect 61628 26908 61684 26910
rect 61964 26850 62020 26852
rect 61964 26798 61966 26850
rect 61966 26798 62018 26850
rect 62018 26798 62020 26850
rect 61964 26796 62020 26798
rect 62188 26290 62244 26292
rect 62188 26238 62190 26290
rect 62190 26238 62242 26290
rect 62242 26238 62244 26290
rect 62188 26236 62244 26238
rect 61516 25564 61572 25620
rect 61292 25452 61348 25508
rect 62188 25394 62244 25396
rect 62188 25342 62190 25394
rect 62190 25342 62242 25394
rect 62242 25342 62244 25394
rect 62188 25340 62244 25342
rect 61740 23938 61796 23940
rect 61740 23886 61742 23938
rect 61742 23886 61794 23938
rect 61794 23886 61796 23938
rect 61740 23884 61796 23886
rect 62076 23938 62132 23940
rect 62076 23886 62078 23938
rect 62078 23886 62130 23938
rect 62130 23886 62132 23938
rect 62076 23884 62132 23886
rect 61852 23548 61908 23604
rect 61292 23324 61348 23380
rect 61292 21980 61348 22036
rect 61516 21698 61572 21700
rect 61516 21646 61518 21698
rect 61518 21646 61570 21698
rect 61570 21646 61572 21698
rect 61516 21644 61572 21646
rect 61292 21586 61348 21588
rect 61292 21534 61294 21586
rect 61294 21534 61346 21586
rect 61346 21534 61348 21586
rect 61292 21532 61348 21534
rect 60956 21420 61012 21476
rect 61628 20748 61684 20804
rect 61740 21532 61796 21588
rect 63980 33234 64036 33236
rect 63980 33182 63982 33234
rect 63982 33182 64034 33234
rect 64034 33182 64036 33234
rect 63980 33180 64036 33182
rect 65660 32620 65716 32676
rect 67452 35980 67508 36036
rect 66220 35644 66276 35700
rect 67900 36204 67956 36260
rect 67564 35532 67620 35588
rect 68348 35586 68404 35588
rect 68348 35534 68350 35586
rect 68350 35534 68402 35586
rect 68402 35534 68404 35586
rect 68348 35532 68404 35534
rect 66668 35420 66724 35476
rect 67116 34860 67172 34916
rect 65996 34636 66052 34692
rect 66444 34524 66500 34580
rect 65996 34130 66052 34132
rect 65996 34078 65998 34130
rect 65998 34078 66050 34130
rect 66050 34078 66052 34130
rect 65996 34076 66052 34078
rect 66444 34076 66500 34132
rect 66668 34076 66724 34132
rect 66556 33346 66612 33348
rect 66556 33294 66558 33346
rect 66558 33294 66610 33346
rect 66610 33294 66612 33346
rect 66556 33292 66612 33294
rect 67116 33852 67172 33908
rect 70476 36988 70532 37044
rect 68832 36874 68888 36876
rect 68832 36822 68834 36874
rect 68834 36822 68886 36874
rect 68886 36822 68888 36874
rect 68832 36820 68888 36822
rect 68936 36874 68992 36876
rect 68936 36822 68938 36874
rect 68938 36822 68990 36874
rect 68990 36822 68992 36874
rect 68936 36820 68992 36822
rect 69040 36874 69096 36876
rect 69040 36822 69042 36874
rect 69042 36822 69094 36874
rect 69094 36822 69096 36874
rect 69040 36820 69096 36822
rect 68684 36316 68740 36372
rect 71148 37772 71204 37828
rect 70476 36316 70532 36372
rect 71708 36652 71764 36708
rect 71148 36092 71204 36148
rect 68832 35306 68888 35308
rect 68832 35254 68834 35306
rect 68834 35254 68886 35306
rect 68886 35254 68888 35306
rect 68832 35252 68888 35254
rect 68936 35306 68992 35308
rect 68936 35254 68938 35306
rect 68938 35254 68990 35306
rect 68990 35254 68992 35306
rect 68936 35252 68992 35254
rect 69040 35306 69096 35308
rect 69040 35254 69042 35306
rect 69042 35254 69094 35306
rect 69094 35254 69096 35306
rect 69040 35252 69096 35254
rect 68684 34860 68740 34916
rect 68832 33738 68888 33740
rect 68832 33686 68834 33738
rect 68834 33686 68886 33738
rect 68886 33686 68888 33738
rect 68832 33684 68888 33686
rect 68936 33738 68992 33740
rect 68936 33686 68938 33738
rect 68938 33686 68990 33738
rect 68990 33686 68992 33738
rect 68936 33684 68992 33686
rect 69040 33738 69096 33740
rect 69040 33686 69042 33738
rect 69042 33686 69094 33738
rect 69094 33686 69096 33738
rect 69040 33684 69096 33686
rect 68460 33292 68516 33348
rect 69468 35532 69524 35588
rect 69580 35474 69636 35476
rect 69580 35422 69582 35474
rect 69582 35422 69634 35474
rect 69634 35422 69636 35474
rect 69580 35420 69636 35422
rect 69468 34748 69524 34804
rect 69244 33180 69300 33236
rect 69692 34972 69748 35028
rect 75404 37996 75460 38052
rect 73164 36540 73220 36596
rect 73500 37212 73556 37268
rect 73164 36316 73220 36372
rect 72828 36258 72884 36260
rect 72828 36206 72830 36258
rect 72830 36206 72882 36258
rect 72882 36206 72884 36258
rect 72828 36204 72884 36206
rect 72492 35868 72548 35924
rect 71708 35756 71764 35812
rect 72268 35810 72324 35812
rect 72268 35758 72270 35810
rect 72270 35758 72322 35810
rect 72322 35758 72324 35810
rect 72268 35756 72324 35758
rect 71372 34802 71428 34804
rect 71372 34750 71374 34802
rect 71374 34750 71426 34802
rect 71426 34750 71428 34802
rect 71372 34748 71428 34750
rect 69692 34524 69748 34580
rect 70140 33906 70196 33908
rect 70140 33854 70142 33906
rect 70142 33854 70194 33906
rect 70194 33854 70196 33906
rect 70140 33852 70196 33854
rect 69580 33516 69636 33572
rect 67228 33068 67284 33124
rect 67452 32674 67508 32676
rect 67452 32622 67454 32674
rect 67454 32622 67506 32674
rect 67506 32622 67508 32674
rect 67452 32620 67508 32622
rect 69356 32620 69412 32676
rect 66780 32562 66836 32564
rect 66780 32510 66782 32562
rect 66782 32510 66834 32562
rect 66834 32510 66836 32562
rect 66780 32508 66836 32510
rect 67564 32562 67620 32564
rect 67564 32510 67566 32562
rect 67566 32510 67618 32562
rect 67618 32510 67620 32562
rect 67564 32508 67620 32510
rect 68832 32170 68888 32172
rect 68832 32118 68834 32170
rect 68834 32118 68886 32170
rect 68886 32118 68888 32170
rect 68832 32116 68888 32118
rect 68936 32170 68992 32172
rect 68936 32118 68938 32170
rect 68938 32118 68990 32170
rect 68990 32118 68992 32170
rect 68936 32116 68992 32118
rect 69040 32170 69096 32172
rect 69040 32118 69042 32170
rect 69042 32118 69094 32170
rect 69094 32118 69096 32170
rect 69040 32116 69096 32118
rect 65884 31890 65940 31892
rect 65884 31838 65886 31890
rect 65886 31838 65938 31890
rect 65938 31838 65940 31890
rect 65884 31836 65940 31838
rect 67564 31724 67620 31780
rect 63644 31554 63700 31556
rect 63644 31502 63646 31554
rect 63646 31502 63698 31554
rect 63698 31502 63700 31554
rect 63644 31500 63700 31502
rect 63308 30770 63364 30772
rect 63308 30718 63310 30770
rect 63310 30718 63362 30770
rect 63362 30718 63364 30770
rect 63308 30716 63364 30718
rect 62524 30156 62580 30212
rect 63868 30882 63924 30884
rect 63868 30830 63870 30882
rect 63870 30830 63922 30882
rect 63922 30830 63924 30882
rect 63868 30828 63924 30830
rect 64316 30828 64372 30884
rect 65436 31500 65492 31556
rect 63868 28812 63924 28868
rect 62636 27804 62692 27860
rect 62412 25506 62468 25508
rect 62412 25454 62414 25506
rect 62414 25454 62466 25506
rect 62466 25454 62468 25506
rect 62412 25452 62468 25454
rect 62860 26290 62916 26292
rect 62860 26238 62862 26290
rect 62862 26238 62914 26290
rect 62914 26238 62916 26290
rect 62860 26236 62916 26238
rect 65100 28754 65156 28756
rect 65100 28702 65102 28754
rect 65102 28702 65154 28754
rect 65154 28702 65156 28754
rect 65100 28700 65156 28702
rect 64204 27916 64260 27972
rect 64428 27692 64484 27748
rect 63084 27020 63140 27076
rect 63868 27074 63924 27076
rect 63868 27022 63870 27074
rect 63870 27022 63922 27074
rect 63922 27022 63924 27074
rect 63868 27020 63924 27022
rect 63308 26460 63364 26516
rect 63756 26908 63812 26964
rect 63980 26850 64036 26852
rect 63980 26798 63982 26850
rect 63982 26798 64034 26850
rect 64034 26798 64036 26850
rect 63980 26796 64036 26798
rect 62860 25676 62916 25732
rect 62636 25506 62692 25508
rect 62636 25454 62638 25506
rect 62638 25454 62690 25506
rect 62690 25454 62692 25506
rect 62636 25452 62692 25454
rect 64204 25618 64260 25620
rect 64204 25566 64206 25618
rect 64206 25566 64258 25618
rect 64258 25566 64260 25618
rect 64204 25564 64260 25566
rect 63308 25506 63364 25508
rect 63308 25454 63310 25506
rect 63310 25454 63362 25506
rect 63362 25454 63364 25506
rect 63308 25452 63364 25454
rect 63084 25228 63140 25284
rect 62412 24834 62468 24836
rect 62412 24782 62414 24834
rect 62414 24782 62466 24834
rect 62466 24782 62468 24834
rect 62412 24780 62468 24782
rect 62748 23154 62804 23156
rect 62748 23102 62750 23154
rect 62750 23102 62802 23154
rect 62802 23102 62804 23154
rect 62748 23100 62804 23102
rect 63868 25394 63924 25396
rect 63868 25342 63870 25394
rect 63870 25342 63922 25394
rect 63922 25342 63924 25394
rect 63868 25340 63924 25342
rect 63980 25116 64036 25172
rect 63420 24946 63476 24948
rect 63420 24894 63422 24946
rect 63422 24894 63474 24946
rect 63474 24894 63476 24946
rect 63420 24892 63476 24894
rect 63532 22540 63588 22596
rect 63756 22258 63812 22260
rect 63756 22206 63758 22258
rect 63758 22206 63810 22258
rect 63810 22206 63812 22258
rect 63756 22204 63812 22206
rect 63756 21810 63812 21812
rect 63756 21758 63758 21810
rect 63758 21758 63810 21810
rect 63810 21758 63812 21810
rect 63756 21756 63812 21758
rect 63308 21644 63364 21700
rect 61852 20748 61908 20804
rect 62972 20802 63028 20804
rect 62972 20750 62974 20802
rect 62974 20750 63026 20802
rect 63026 20750 63028 20802
rect 62972 20748 63028 20750
rect 61964 20636 62020 20692
rect 65772 31554 65828 31556
rect 65772 31502 65774 31554
rect 65774 31502 65826 31554
rect 65826 31502 65828 31554
rect 65772 31500 65828 31502
rect 66780 31388 66836 31444
rect 67228 31388 67284 31444
rect 67340 31500 67396 31556
rect 66108 30994 66164 30996
rect 66108 30942 66110 30994
rect 66110 30942 66162 30994
rect 66162 30942 66164 30994
rect 66108 30940 66164 30942
rect 68236 31612 68292 31668
rect 68460 31388 68516 31444
rect 67564 30994 67620 30996
rect 67564 30942 67566 30994
rect 67566 30942 67618 30994
rect 67618 30942 67620 30994
rect 67564 30940 67620 30942
rect 66108 30716 66164 30772
rect 66108 30210 66164 30212
rect 66108 30158 66110 30210
rect 66110 30158 66162 30210
rect 66162 30158 66164 30210
rect 66108 30156 66164 30158
rect 68572 30994 68628 30996
rect 68572 30942 68574 30994
rect 68574 30942 68626 30994
rect 68626 30942 68628 30994
rect 68572 30940 68628 30942
rect 69132 30994 69188 30996
rect 69132 30942 69134 30994
rect 69134 30942 69186 30994
rect 69186 30942 69188 30994
rect 69132 30940 69188 30942
rect 68832 30602 68888 30604
rect 68832 30550 68834 30602
rect 68834 30550 68886 30602
rect 68886 30550 68888 30602
rect 68832 30548 68888 30550
rect 68936 30602 68992 30604
rect 68936 30550 68938 30602
rect 68938 30550 68990 30602
rect 68990 30550 68992 30602
rect 68936 30548 68992 30550
rect 69040 30602 69096 30604
rect 69040 30550 69042 30602
rect 69042 30550 69094 30602
rect 69094 30550 69096 30602
rect 69040 30548 69096 30550
rect 68460 30268 68516 30324
rect 67788 30098 67844 30100
rect 67788 30046 67790 30098
rect 67790 30046 67842 30098
rect 67842 30046 67844 30098
rect 67788 30044 67844 30046
rect 67004 29932 67060 29988
rect 68460 30098 68516 30100
rect 68460 30046 68462 30098
rect 68462 30046 68514 30098
rect 68514 30046 68516 30098
rect 68460 30044 68516 30046
rect 67900 29932 67956 29988
rect 67900 29484 67956 29540
rect 68236 29538 68292 29540
rect 68236 29486 68238 29538
rect 68238 29486 68290 29538
rect 68290 29486 68292 29538
rect 68236 29484 68292 29486
rect 66780 29260 66836 29316
rect 67340 29314 67396 29316
rect 67340 29262 67342 29314
rect 67342 29262 67394 29314
rect 67394 29262 67396 29314
rect 67340 29260 67396 29262
rect 68572 29260 68628 29316
rect 68832 29034 68888 29036
rect 68832 28982 68834 29034
rect 68834 28982 68886 29034
rect 68886 28982 68888 29034
rect 68832 28980 68888 28982
rect 68936 29034 68992 29036
rect 68936 28982 68938 29034
rect 68938 28982 68990 29034
rect 68990 28982 68992 29034
rect 68936 28980 68992 28982
rect 69040 29034 69096 29036
rect 69040 28982 69042 29034
rect 69042 28982 69094 29034
rect 69094 28982 69096 29034
rect 69040 28980 69096 28982
rect 65996 28812 66052 28868
rect 65772 28754 65828 28756
rect 65772 28702 65774 28754
rect 65774 28702 65826 28754
rect 65826 28702 65828 28754
rect 65772 28700 65828 28702
rect 65884 28588 65940 28644
rect 65548 27916 65604 27972
rect 64876 27244 64932 27300
rect 65436 26514 65492 26516
rect 65436 26462 65438 26514
rect 65438 26462 65490 26514
rect 65490 26462 65492 26514
rect 65436 26460 65492 26462
rect 66668 28588 66724 28644
rect 67340 28642 67396 28644
rect 67340 28590 67342 28642
rect 67342 28590 67394 28642
rect 67394 28590 67396 28642
rect 67340 28588 67396 28590
rect 65996 27970 66052 27972
rect 65996 27918 65998 27970
rect 65998 27918 66050 27970
rect 66050 27918 66052 27970
rect 65996 27916 66052 27918
rect 66332 27916 66388 27972
rect 65996 27298 66052 27300
rect 65996 27246 65998 27298
rect 65998 27246 66050 27298
rect 66050 27246 66052 27298
rect 65996 27244 66052 27246
rect 68236 28530 68292 28532
rect 68236 28478 68238 28530
rect 68238 28478 68290 28530
rect 68290 28478 68292 28530
rect 68236 28476 68292 28478
rect 67564 27916 67620 27972
rect 71148 34242 71204 34244
rect 71148 34190 71150 34242
rect 71150 34190 71202 34242
rect 71202 34190 71204 34242
rect 71148 34188 71204 34190
rect 72268 34972 72324 35028
rect 71484 34188 71540 34244
rect 71820 33852 71876 33908
rect 72156 33852 72212 33908
rect 72604 35810 72660 35812
rect 72604 35758 72606 35810
rect 72606 35758 72658 35810
rect 72658 35758 72660 35810
rect 72604 35756 72660 35758
rect 72492 34802 72548 34804
rect 72492 34750 72494 34802
rect 72494 34750 72546 34802
rect 72546 34750 72548 34802
rect 72492 34748 72548 34750
rect 73388 36316 73444 36372
rect 73276 36092 73332 36148
rect 74060 36594 74116 36596
rect 74060 36542 74062 36594
rect 74062 36542 74114 36594
rect 74114 36542 74116 36594
rect 74060 36540 74116 36542
rect 75404 36540 75460 36596
rect 74172 36428 74228 36484
rect 77868 38444 77924 38500
rect 77084 37324 77140 37380
rect 74956 36204 75012 36260
rect 73948 34860 74004 34916
rect 73612 34188 73668 34244
rect 70588 33068 70644 33124
rect 70700 32508 70756 32564
rect 69804 31778 69860 31780
rect 69804 31726 69806 31778
rect 69806 31726 69858 31778
rect 69858 31726 69860 31778
rect 69804 31724 69860 31726
rect 69580 31666 69636 31668
rect 69580 31614 69582 31666
rect 69582 31614 69634 31666
rect 69634 31614 69636 31666
rect 69580 31612 69636 31614
rect 69580 31218 69636 31220
rect 69580 31166 69582 31218
rect 69582 31166 69634 31218
rect 69634 31166 69636 31218
rect 69580 31164 69636 31166
rect 71260 31666 71316 31668
rect 71260 31614 71262 31666
rect 71262 31614 71314 31666
rect 71314 31614 71316 31666
rect 71260 31612 71316 31614
rect 70812 31164 70868 31220
rect 69468 30268 69524 30324
rect 69468 30098 69524 30100
rect 69468 30046 69470 30098
rect 69470 30046 69522 30098
rect 69522 30046 69524 30098
rect 69468 30044 69524 30046
rect 69692 30098 69748 30100
rect 69692 30046 69694 30098
rect 69694 30046 69746 30098
rect 69746 30046 69748 30098
rect 69692 30044 69748 30046
rect 69580 29484 69636 29540
rect 71036 31500 71092 31556
rect 70812 30268 70868 30324
rect 71148 30156 71204 30212
rect 70812 29986 70868 29988
rect 70812 29934 70814 29986
rect 70814 29934 70866 29986
rect 70866 29934 70868 29986
rect 70812 29932 70868 29934
rect 71932 33068 71988 33124
rect 72380 33068 72436 33124
rect 71820 31500 71876 31556
rect 71932 31388 71988 31444
rect 71932 31218 71988 31220
rect 71932 31166 71934 31218
rect 71934 31166 71986 31218
rect 71986 31166 71988 31218
rect 71932 31164 71988 31166
rect 71708 30940 71764 30996
rect 72044 30716 72100 30772
rect 71820 29932 71876 29988
rect 71820 29708 71876 29764
rect 70812 29426 70868 29428
rect 70812 29374 70814 29426
rect 70814 29374 70866 29426
rect 70866 29374 70868 29426
rect 70812 29372 70868 29374
rect 70028 28812 70084 28868
rect 70028 28588 70084 28644
rect 69468 28530 69524 28532
rect 69468 28478 69470 28530
rect 69470 28478 69522 28530
rect 69522 28478 69524 28530
rect 69468 28476 69524 28478
rect 68832 27466 68888 27468
rect 68832 27414 68834 27466
rect 68834 27414 68886 27466
rect 68886 27414 68888 27466
rect 68832 27412 68888 27414
rect 68936 27466 68992 27468
rect 68936 27414 68938 27466
rect 68938 27414 68990 27466
rect 68990 27414 68992 27466
rect 68936 27412 68992 27414
rect 69040 27466 69096 27468
rect 69040 27414 69042 27466
rect 69042 27414 69094 27466
rect 69094 27414 69096 27466
rect 69244 27468 69300 27524
rect 70812 28588 70868 28644
rect 71372 29426 71428 29428
rect 71372 29374 71374 29426
rect 71374 29374 71426 29426
rect 71426 29374 71428 29426
rect 71372 29372 71428 29374
rect 71036 28642 71092 28644
rect 71036 28590 71038 28642
rect 71038 28590 71090 28642
rect 71090 28590 71092 28642
rect 71036 28588 71092 28590
rect 69040 27412 69096 27414
rect 68348 27074 68404 27076
rect 68348 27022 68350 27074
rect 68350 27022 68402 27074
rect 68402 27022 68404 27074
rect 68348 27020 68404 27022
rect 69468 27074 69524 27076
rect 69468 27022 69470 27074
rect 69470 27022 69522 27074
rect 69522 27022 69524 27074
rect 69468 27020 69524 27022
rect 65212 26124 65268 26180
rect 64540 24946 64596 24948
rect 64540 24894 64542 24946
rect 64542 24894 64594 24946
rect 64594 24894 64596 24946
rect 64540 24892 64596 24894
rect 64652 25676 64708 25732
rect 63980 21532 64036 21588
rect 64092 23548 64148 23604
rect 62412 20076 62468 20132
rect 61516 19234 61572 19236
rect 61516 19182 61518 19234
rect 61518 19182 61570 19234
rect 61570 19182 61572 19234
rect 61516 19180 61572 19182
rect 63084 20130 63140 20132
rect 63084 20078 63086 20130
rect 63086 20078 63138 20130
rect 63138 20078 63140 20130
rect 63084 20076 63140 20078
rect 63196 19234 63252 19236
rect 63196 19182 63198 19234
rect 63198 19182 63250 19234
rect 63250 19182 63252 19234
rect 63196 19180 63252 19182
rect 61292 18450 61348 18452
rect 61292 18398 61294 18450
rect 61294 18398 61346 18450
rect 61346 18398 61348 18450
rect 61292 18396 61348 18398
rect 60396 15314 60452 15316
rect 60396 15262 60398 15314
rect 60398 15262 60450 15314
rect 60450 15262 60452 15314
rect 60396 15260 60452 15262
rect 61180 18284 61236 18340
rect 60508 14364 60564 14420
rect 60284 14252 60340 14308
rect 59388 12796 59444 12852
rect 59172 12570 59228 12572
rect 59172 12518 59174 12570
rect 59174 12518 59226 12570
rect 59226 12518 59228 12570
rect 59172 12516 59228 12518
rect 59276 12570 59332 12572
rect 59276 12518 59278 12570
rect 59278 12518 59330 12570
rect 59330 12518 59332 12570
rect 59276 12516 59332 12518
rect 59380 12570 59436 12572
rect 59380 12518 59382 12570
rect 59382 12518 59434 12570
rect 59434 12518 59436 12570
rect 59380 12516 59436 12518
rect 58940 11282 58996 11284
rect 58940 11230 58942 11282
rect 58942 11230 58994 11282
rect 58994 11230 58996 11282
rect 58940 11228 58996 11230
rect 59500 11228 59556 11284
rect 59724 11900 59780 11956
rect 59172 11002 59228 11004
rect 59172 10950 59174 11002
rect 59174 10950 59226 11002
rect 59226 10950 59228 11002
rect 59172 10948 59228 10950
rect 59276 11002 59332 11004
rect 59276 10950 59278 11002
rect 59278 10950 59330 11002
rect 59330 10950 59332 11002
rect 59276 10948 59332 10950
rect 59380 11002 59436 11004
rect 59380 10950 59382 11002
rect 59382 10950 59434 11002
rect 59434 10950 59436 11002
rect 59380 10948 59436 10950
rect 59172 9434 59228 9436
rect 59172 9382 59174 9434
rect 59174 9382 59226 9434
rect 59226 9382 59228 9434
rect 59172 9380 59228 9382
rect 59276 9434 59332 9436
rect 59276 9382 59278 9434
rect 59278 9382 59330 9434
rect 59330 9382 59332 9434
rect 59276 9380 59332 9382
rect 59380 9434 59436 9436
rect 59380 9382 59382 9434
rect 59382 9382 59434 9434
rect 59434 9382 59436 9434
rect 59380 9380 59436 9382
rect 58828 8204 58884 8260
rect 58828 7532 58884 7588
rect 59052 8092 59108 8148
rect 59172 7866 59228 7868
rect 59172 7814 59174 7866
rect 59174 7814 59226 7866
rect 59226 7814 59228 7866
rect 59172 7812 59228 7814
rect 59276 7866 59332 7868
rect 59276 7814 59278 7866
rect 59278 7814 59330 7866
rect 59330 7814 59332 7866
rect 59276 7812 59332 7814
rect 59380 7866 59436 7868
rect 59380 7814 59382 7866
rect 59382 7814 59434 7866
rect 59434 7814 59436 7866
rect 59380 7812 59436 7814
rect 59612 8258 59668 8260
rect 59612 8206 59614 8258
rect 59614 8206 59666 8258
rect 59666 8206 59668 8258
rect 59612 8204 59668 8206
rect 59388 7196 59444 7252
rect 58940 7084 58996 7140
rect 59052 6748 59108 6804
rect 58268 5068 58324 5124
rect 58940 6130 58996 6132
rect 58940 6078 58942 6130
rect 58942 6078 58994 6130
rect 58994 6078 58996 6130
rect 58940 6076 58996 6078
rect 59164 6578 59220 6580
rect 59164 6526 59166 6578
rect 59166 6526 59218 6578
rect 59218 6526 59220 6578
rect 59164 6524 59220 6526
rect 59172 6298 59228 6300
rect 59172 6246 59174 6298
rect 59174 6246 59226 6298
rect 59226 6246 59228 6298
rect 59172 6244 59228 6246
rect 59276 6298 59332 6300
rect 59276 6246 59278 6298
rect 59278 6246 59330 6298
rect 59330 6246 59332 6298
rect 59276 6244 59332 6246
rect 59380 6298 59436 6300
rect 59380 6246 59382 6298
rect 59382 6246 59434 6298
rect 59434 6246 59436 6298
rect 59380 6244 59436 6246
rect 58380 5964 58436 6020
rect 58828 5906 58884 5908
rect 58828 5854 58830 5906
rect 58830 5854 58882 5906
rect 58882 5854 58884 5906
rect 58828 5852 58884 5854
rect 58492 5794 58548 5796
rect 58492 5742 58494 5794
rect 58494 5742 58546 5794
rect 58546 5742 58548 5794
rect 58492 5740 58548 5742
rect 58380 4732 58436 4788
rect 58604 4508 58660 4564
rect 58044 4338 58100 4340
rect 58044 4286 58046 4338
rect 58046 4286 58098 4338
rect 58098 4286 58100 4338
rect 58044 4284 58100 4286
rect 57932 4172 57988 4228
rect 57820 3948 57876 4004
rect 58716 4898 58772 4900
rect 58716 4846 58718 4898
rect 58718 4846 58770 4898
rect 58770 4846 58772 4898
rect 58716 4844 58772 4846
rect 58716 4396 58772 4452
rect 59164 5068 59220 5124
rect 58940 4898 58996 4900
rect 58940 4846 58942 4898
rect 58942 4846 58994 4898
rect 58994 4846 58996 4898
rect 58940 4844 58996 4846
rect 59172 4730 59228 4732
rect 59172 4678 59174 4730
rect 59174 4678 59226 4730
rect 59226 4678 59228 4730
rect 59172 4676 59228 4678
rect 59276 4730 59332 4732
rect 59276 4678 59278 4730
rect 59278 4678 59330 4730
rect 59330 4678 59332 4730
rect 59276 4676 59332 4678
rect 59380 4730 59436 4732
rect 59380 4678 59382 4730
rect 59382 4678 59434 4730
rect 59434 4678 59436 4730
rect 59380 4676 59436 4678
rect 58156 3948 58212 4004
rect 58044 3276 58100 3332
rect 58156 3388 58212 3444
rect 57484 2604 57540 2660
rect 58940 3442 58996 3444
rect 58940 3390 58942 3442
rect 58942 3390 58994 3442
rect 58994 3390 58996 3442
rect 58940 3388 58996 3390
rect 61068 13858 61124 13860
rect 61068 13806 61070 13858
rect 61070 13806 61122 13858
rect 61122 13806 61124 13858
rect 61068 13804 61124 13806
rect 60620 13020 60676 13076
rect 59948 12796 60004 12852
rect 60172 12962 60228 12964
rect 60172 12910 60174 12962
rect 60174 12910 60226 12962
rect 60226 12910 60228 12962
rect 60172 12908 60228 12910
rect 60956 11954 61012 11956
rect 60956 11902 60958 11954
rect 60958 11902 61010 11954
rect 61010 11902 61012 11954
rect 60956 11900 61012 11902
rect 60508 11282 60564 11284
rect 60508 11230 60510 11282
rect 60510 11230 60562 11282
rect 60562 11230 60564 11282
rect 60508 11228 60564 11230
rect 59948 9714 60004 9716
rect 59948 9662 59950 9714
rect 59950 9662 60002 9714
rect 60002 9662 60004 9714
rect 59948 9660 60004 9662
rect 60172 9436 60228 9492
rect 60844 8876 60900 8932
rect 62748 18956 62804 19012
rect 61740 17554 61796 17556
rect 61740 17502 61742 17554
rect 61742 17502 61794 17554
rect 61794 17502 61796 17554
rect 62076 17666 62132 17668
rect 62076 17614 62078 17666
rect 62078 17614 62130 17666
rect 62130 17614 62132 17666
rect 62076 17612 62132 17614
rect 61740 17500 61796 17502
rect 61292 17164 61348 17220
rect 61404 17052 61460 17108
rect 61852 16940 61908 16996
rect 61404 16828 61460 16884
rect 61628 16380 61684 16436
rect 61740 16828 61796 16884
rect 62076 16380 62132 16436
rect 61964 16210 62020 16212
rect 61964 16158 61966 16210
rect 61966 16158 62018 16210
rect 62018 16158 62020 16210
rect 61964 16156 62020 16158
rect 62636 16380 62692 16436
rect 62300 16268 62356 16324
rect 62636 16210 62692 16212
rect 62636 16158 62638 16210
rect 62638 16158 62690 16210
rect 62690 16158 62692 16210
rect 62636 16156 62692 16158
rect 61628 15874 61684 15876
rect 61628 15822 61630 15874
rect 61630 15822 61682 15874
rect 61682 15822 61684 15874
rect 61628 15820 61684 15822
rect 62076 15820 62132 15876
rect 62300 15596 62356 15652
rect 63868 20076 63924 20132
rect 63644 19964 63700 20020
rect 65212 25564 65268 25620
rect 68460 26850 68516 26852
rect 68460 26798 68462 26850
rect 68462 26798 68514 26850
rect 68514 26798 68516 26850
rect 68460 26796 68516 26798
rect 65996 26178 66052 26180
rect 65996 26126 65998 26178
rect 65998 26126 66050 26178
rect 66050 26126 66052 26178
rect 65996 26124 66052 26126
rect 65436 25340 65492 25396
rect 64764 24946 64820 24948
rect 64764 24894 64766 24946
rect 64766 24894 64818 24946
rect 64818 24894 64820 24946
rect 64764 24892 64820 24894
rect 64988 24668 65044 24724
rect 65436 24722 65492 24724
rect 65436 24670 65438 24722
rect 65438 24670 65490 24722
rect 65490 24670 65492 24722
rect 65436 24668 65492 24670
rect 65996 24892 66052 24948
rect 66332 25340 66388 25396
rect 65548 23996 65604 24052
rect 64988 23548 65044 23604
rect 65324 23548 65380 23604
rect 64876 23436 64932 23492
rect 66780 25564 66836 25620
rect 67116 26066 67172 26068
rect 67116 26014 67118 26066
rect 67118 26014 67170 26066
rect 67170 26014 67172 26066
rect 67116 26012 67172 26014
rect 67676 26066 67732 26068
rect 67676 26014 67678 26066
rect 67678 26014 67730 26066
rect 67730 26014 67732 26066
rect 67676 26012 67732 26014
rect 67788 25618 67844 25620
rect 67788 25566 67790 25618
rect 67790 25566 67842 25618
rect 67842 25566 67844 25618
rect 67788 25564 67844 25566
rect 67004 25340 67060 25396
rect 66668 25228 66724 25284
rect 66780 24946 66836 24948
rect 66780 24894 66782 24946
rect 66782 24894 66834 24946
rect 66834 24894 66836 24946
rect 66780 24892 66836 24894
rect 66780 24556 66836 24612
rect 67676 25340 67732 25396
rect 68012 26236 68068 26292
rect 71148 27468 71204 27524
rect 69804 27020 69860 27076
rect 70476 27020 70532 27076
rect 69916 26796 69972 26852
rect 69580 26290 69636 26292
rect 69580 26238 69582 26290
rect 69582 26238 69634 26290
rect 69634 26238 69636 26290
rect 69580 26236 69636 26238
rect 68832 25898 68888 25900
rect 67900 25228 67956 25284
rect 68124 25788 68180 25844
rect 68832 25846 68834 25898
rect 68834 25846 68886 25898
rect 68886 25846 68888 25898
rect 68832 25844 68888 25846
rect 68936 25898 68992 25900
rect 68936 25846 68938 25898
rect 68938 25846 68990 25898
rect 68990 25846 68992 25898
rect 68936 25844 68992 25846
rect 69040 25898 69096 25900
rect 69040 25846 69042 25898
rect 69042 25846 69094 25898
rect 69094 25846 69096 25898
rect 69040 25844 69096 25846
rect 67788 24722 67844 24724
rect 67788 24670 67790 24722
rect 67790 24670 67842 24722
rect 67842 24670 67844 24722
rect 67788 24668 67844 24670
rect 67228 24556 67284 24612
rect 67116 23996 67172 24052
rect 66332 23772 66388 23828
rect 65100 22370 65156 22372
rect 65100 22318 65102 22370
rect 65102 22318 65154 22370
rect 65154 22318 65156 22370
rect 65100 22316 65156 22318
rect 64876 22258 64932 22260
rect 64876 22206 64878 22258
rect 64878 22206 64930 22258
rect 64930 22206 64932 22258
rect 64876 22204 64932 22206
rect 65324 22204 65380 22260
rect 64540 21756 64596 21812
rect 64316 21586 64372 21588
rect 64316 21534 64318 21586
rect 64318 21534 64370 21586
rect 64370 21534 64372 21586
rect 64316 21532 64372 21534
rect 64652 21644 64708 21700
rect 63980 19740 64036 19796
rect 64204 20018 64260 20020
rect 64204 19966 64206 20018
rect 64206 19966 64258 20018
rect 64258 19966 64260 20018
rect 64204 19964 64260 19966
rect 63980 19292 64036 19348
rect 64092 19234 64148 19236
rect 64092 19182 64094 19234
rect 64094 19182 64146 19234
rect 64146 19182 64148 19234
rect 64092 19180 64148 19182
rect 64316 19180 64372 19236
rect 64204 19068 64260 19124
rect 63420 18172 63476 18228
rect 63196 17724 63252 17780
rect 62860 16210 62916 16212
rect 62860 16158 62862 16210
rect 62862 16158 62914 16210
rect 62914 16158 62916 16210
rect 62860 16156 62916 16158
rect 63084 17106 63140 17108
rect 63084 17054 63086 17106
rect 63086 17054 63138 17106
rect 63138 17054 63140 17106
rect 63084 17052 63140 17054
rect 63420 16828 63476 16884
rect 63644 16210 63700 16212
rect 63644 16158 63646 16210
rect 63646 16158 63698 16210
rect 63698 16158 63700 16210
rect 63644 16156 63700 16158
rect 62972 15932 63028 15988
rect 62972 15372 63028 15428
rect 61516 15260 61572 15316
rect 61292 14364 61348 14420
rect 61404 14306 61460 14308
rect 61404 14254 61406 14306
rect 61406 14254 61458 14306
rect 61458 14254 61460 14306
rect 61404 14252 61460 14254
rect 61516 13804 61572 13860
rect 62524 14252 62580 14308
rect 61628 13468 61684 13524
rect 61292 12962 61348 12964
rect 61292 12910 61294 12962
rect 61294 12910 61346 12962
rect 61346 12910 61348 12962
rect 61292 12908 61348 12910
rect 61740 12850 61796 12852
rect 61740 12798 61742 12850
rect 61742 12798 61794 12850
rect 61794 12798 61796 12850
rect 61740 12796 61796 12798
rect 61964 12684 62020 12740
rect 62412 12738 62468 12740
rect 62412 12686 62414 12738
rect 62414 12686 62466 12738
rect 62466 12686 62468 12738
rect 62412 12684 62468 12686
rect 62412 12460 62468 12516
rect 62076 12290 62132 12292
rect 62076 12238 62078 12290
rect 62078 12238 62130 12290
rect 62130 12238 62132 12290
rect 62076 12236 62132 12238
rect 61964 12124 62020 12180
rect 61516 10556 61572 10612
rect 61628 9996 61684 10052
rect 61964 9996 62020 10052
rect 61852 9884 61908 9940
rect 62300 11506 62356 11508
rect 62300 11454 62302 11506
rect 62302 11454 62354 11506
rect 62354 11454 62356 11506
rect 62300 11452 62356 11454
rect 62188 10780 62244 10836
rect 62524 12290 62580 12292
rect 62524 12238 62526 12290
rect 62526 12238 62578 12290
rect 62578 12238 62580 12290
rect 62524 12236 62580 12238
rect 62972 12684 63028 12740
rect 63084 12572 63140 12628
rect 63308 15036 63364 15092
rect 62860 12124 62916 12180
rect 63420 12290 63476 12292
rect 63420 12238 63422 12290
rect 63422 12238 63474 12290
rect 63474 12238 63476 12290
rect 63420 12236 63476 12238
rect 63308 11506 63364 11508
rect 63308 11454 63310 11506
rect 63310 11454 63362 11506
rect 63362 11454 63364 11506
rect 63308 11452 63364 11454
rect 63308 10892 63364 10948
rect 63196 10780 63252 10836
rect 62188 10610 62244 10612
rect 62188 10558 62190 10610
rect 62190 10558 62242 10610
rect 62242 10558 62244 10610
rect 62188 10556 62244 10558
rect 63532 11788 63588 11844
rect 65212 20860 65268 20916
rect 63868 17164 63924 17220
rect 63868 16940 63924 16996
rect 64428 17052 64484 17108
rect 63980 15596 64036 15652
rect 64092 16940 64148 16996
rect 63868 15372 63924 15428
rect 64092 15148 64148 15204
rect 64204 16044 64260 16100
rect 63980 14700 64036 14756
rect 64428 16882 64484 16884
rect 64428 16830 64430 16882
rect 64430 16830 64482 16882
rect 64482 16830 64484 16882
rect 64428 16828 64484 16830
rect 64316 15932 64372 15988
rect 64764 19906 64820 19908
rect 64764 19854 64766 19906
rect 64766 19854 64818 19906
rect 64818 19854 64820 19906
rect 64764 19852 64820 19854
rect 64764 18396 64820 18452
rect 64652 17388 64708 17444
rect 65548 22258 65604 22260
rect 65548 22206 65550 22258
rect 65550 22206 65602 22258
rect 65602 22206 65604 22258
rect 65548 22204 65604 22206
rect 66444 23714 66500 23716
rect 66444 23662 66446 23714
rect 66446 23662 66498 23714
rect 66498 23662 66500 23714
rect 66444 23660 66500 23662
rect 66108 23154 66164 23156
rect 66108 23102 66110 23154
rect 66110 23102 66162 23154
rect 66162 23102 66164 23154
rect 66108 23100 66164 23102
rect 65660 22092 65716 22148
rect 65996 22988 66052 23044
rect 65772 21868 65828 21924
rect 65548 21698 65604 21700
rect 65548 21646 65550 21698
rect 65550 21646 65602 21698
rect 65602 21646 65604 21698
rect 65548 21644 65604 21646
rect 65324 20690 65380 20692
rect 65324 20638 65326 20690
rect 65326 20638 65378 20690
rect 65378 20638 65380 20690
rect 65324 20636 65380 20638
rect 65436 21586 65492 21588
rect 65436 21534 65438 21586
rect 65438 21534 65490 21586
rect 65490 21534 65492 21586
rect 65436 21532 65492 21534
rect 65660 21532 65716 21588
rect 65548 20802 65604 20804
rect 65548 20750 65550 20802
rect 65550 20750 65602 20802
rect 65602 20750 65604 20802
rect 65548 20748 65604 20750
rect 65884 21532 65940 21588
rect 65772 20636 65828 20692
rect 65436 19068 65492 19124
rect 66668 22370 66724 22372
rect 66668 22318 66670 22370
rect 66670 22318 66722 22370
rect 66722 22318 66724 22370
rect 66668 22316 66724 22318
rect 67116 22316 67172 22372
rect 67340 23996 67396 24052
rect 67900 23772 67956 23828
rect 67452 23714 67508 23716
rect 67452 23662 67454 23714
rect 67454 23662 67506 23714
rect 67506 23662 67508 23714
rect 67452 23660 67508 23662
rect 66108 22204 66164 22260
rect 66108 21756 66164 21812
rect 66444 22092 66500 22148
rect 66332 21474 66388 21476
rect 66332 21422 66334 21474
rect 66334 21422 66386 21474
rect 66386 21422 66388 21474
rect 66332 21420 66388 21422
rect 66108 20748 66164 20804
rect 66556 21586 66612 21588
rect 66556 21534 66558 21586
rect 66558 21534 66610 21586
rect 66610 21534 66612 21586
rect 66556 21532 66612 21534
rect 67228 21980 67284 22036
rect 67900 22146 67956 22148
rect 67900 22094 67902 22146
rect 67902 22094 67954 22146
rect 67954 22094 67956 22146
rect 67900 22092 67956 22094
rect 67116 21532 67172 21588
rect 67452 21868 67508 21924
rect 66668 20748 66724 20804
rect 66332 19852 66388 19908
rect 65884 18450 65940 18452
rect 65884 18398 65886 18450
rect 65886 18398 65938 18450
rect 65938 18398 65940 18450
rect 65884 18396 65940 18398
rect 65772 18284 65828 18340
rect 66108 18620 66164 18676
rect 65324 17442 65380 17444
rect 65324 17390 65326 17442
rect 65326 17390 65378 17442
rect 65378 17390 65380 17442
rect 65324 17388 65380 17390
rect 64652 17164 64708 17220
rect 64764 16828 64820 16884
rect 64988 16322 65044 16324
rect 64988 16270 64990 16322
rect 64990 16270 65042 16322
rect 65042 16270 65044 16322
rect 64988 16268 65044 16270
rect 64652 15874 64708 15876
rect 64652 15822 64654 15874
rect 64654 15822 64706 15874
rect 64706 15822 64708 15874
rect 64652 15820 64708 15822
rect 65324 15202 65380 15204
rect 65324 15150 65326 15202
rect 65326 15150 65378 15202
rect 65378 15150 65380 15202
rect 65324 15148 65380 15150
rect 64652 14924 64708 14980
rect 65548 16268 65604 16324
rect 64652 13804 64708 13860
rect 64988 13692 65044 13748
rect 64428 13074 64484 13076
rect 64428 13022 64430 13074
rect 64430 13022 64482 13074
rect 64482 13022 64484 13074
rect 64428 13020 64484 13022
rect 65436 13858 65492 13860
rect 65436 13806 65438 13858
rect 65438 13806 65490 13858
rect 65490 13806 65492 13858
rect 65436 13804 65492 13806
rect 65548 13356 65604 13412
rect 65548 13132 65604 13188
rect 65772 16940 65828 16996
rect 65884 15820 65940 15876
rect 66220 16098 66276 16100
rect 66220 16046 66222 16098
rect 66222 16046 66274 16098
rect 66274 16046 66276 16098
rect 66220 16044 66276 16046
rect 65324 12684 65380 12740
rect 65772 15372 65828 15428
rect 66108 14418 66164 14420
rect 66108 14366 66110 14418
rect 66110 14366 66162 14418
rect 66162 14366 66164 14418
rect 66108 14364 66164 14366
rect 63756 11900 63812 11956
rect 63868 12236 63924 12292
rect 63756 11506 63812 11508
rect 63756 11454 63758 11506
rect 63758 11454 63810 11506
rect 63810 11454 63812 11506
rect 63756 11452 63812 11454
rect 63532 10892 63588 10948
rect 63420 10050 63476 10052
rect 63420 9998 63422 10050
rect 63422 9998 63474 10050
rect 63474 9998 63476 10050
rect 63420 9996 63476 9998
rect 62412 9660 62468 9716
rect 59724 6690 59780 6692
rect 59724 6638 59726 6690
rect 59726 6638 59778 6690
rect 59778 6638 59780 6690
rect 59724 6636 59780 6638
rect 60396 8370 60452 8372
rect 60396 8318 60398 8370
rect 60398 8318 60450 8370
rect 60450 8318 60452 8370
rect 60396 8316 60452 8318
rect 60284 8258 60340 8260
rect 60284 8206 60286 8258
rect 60286 8206 60338 8258
rect 60338 8206 60340 8258
rect 60284 8204 60340 8206
rect 60732 7644 60788 7700
rect 59948 6636 60004 6692
rect 60060 7196 60116 7252
rect 60284 7084 60340 7140
rect 60172 6466 60228 6468
rect 60172 6414 60174 6466
rect 60174 6414 60226 6466
rect 60226 6414 60228 6466
rect 60172 6412 60228 6414
rect 60060 6300 60116 6356
rect 59948 5794 60004 5796
rect 59948 5742 59950 5794
rect 59950 5742 60002 5794
rect 60002 5742 60004 5794
rect 59948 5740 60004 5742
rect 60060 5292 60116 5348
rect 60620 7308 60676 7364
rect 60508 6524 60564 6580
rect 60508 5180 60564 5236
rect 59612 5068 59668 5124
rect 60396 5010 60452 5012
rect 60396 4958 60398 5010
rect 60398 4958 60450 5010
rect 60450 4958 60452 5010
rect 60396 4956 60452 4958
rect 61628 8370 61684 8372
rect 61628 8318 61630 8370
rect 61630 8318 61682 8370
rect 61682 8318 61684 8370
rect 61628 8316 61684 8318
rect 61068 8204 61124 8260
rect 63420 9714 63476 9716
rect 63420 9662 63422 9714
rect 63422 9662 63474 9714
rect 63474 9662 63476 9714
rect 63420 9660 63476 9662
rect 62748 9436 62804 9492
rect 63084 9436 63140 9492
rect 62860 9324 62916 9380
rect 62748 9266 62804 9268
rect 62748 9214 62750 9266
rect 62750 9214 62802 9266
rect 62802 9214 62804 9266
rect 62748 9212 62804 9214
rect 62412 8876 62468 8932
rect 62412 8316 62468 8372
rect 62972 8316 63028 8372
rect 63532 9436 63588 9492
rect 63532 9266 63588 9268
rect 63532 9214 63534 9266
rect 63534 9214 63586 9266
rect 63586 9214 63588 9266
rect 63532 9212 63588 9214
rect 61292 7756 61348 7812
rect 63084 7698 63140 7700
rect 63084 7646 63086 7698
rect 63086 7646 63138 7698
rect 63138 7646 63140 7698
rect 63084 7644 63140 7646
rect 61292 7420 61348 7476
rect 61068 6636 61124 6692
rect 61404 7084 61460 7140
rect 62076 6972 62132 7028
rect 61852 6188 61908 6244
rect 62860 6972 62916 7028
rect 63532 7644 63588 7700
rect 63196 7362 63252 7364
rect 63196 7310 63198 7362
rect 63198 7310 63250 7362
rect 63250 7310 63252 7362
rect 63196 7308 63252 7310
rect 63420 6300 63476 6356
rect 63868 11116 63924 11172
rect 65436 12124 65492 12180
rect 64764 11170 64820 11172
rect 64764 11118 64766 11170
rect 64766 11118 64818 11170
rect 64818 11118 64820 11170
rect 64764 11116 64820 11118
rect 65548 12066 65604 12068
rect 65548 12014 65550 12066
rect 65550 12014 65602 12066
rect 65602 12014 65604 12066
rect 65548 12012 65604 12014
rect 64652 10220 64708 10276
rect 64540 9996 64596 10052
rect 65548 9938 65604 9940
rect 65548 9886 65550 9938
rect 65550 9886 65602 9938
rect 65602 9886 65604 9938
rect 65548 9884 65604 9886
rect 66108 13634 66164 13636
rect 66108 13582 66110 13634
rect 66110 13582 66162 13634
rect 66162 13582 66164 13634
rect 66108 13580 66164 13582
rect 66444 16940 66500 16996
rect 67228 20412 67284 20468
rect 67564 21532 67620 21588
rect 67452 21474 67508 21476
rect 67452 21422 67454 21474
rect 67454 21422 67506 21474
rect 67506 21422 67508 21474
rect 67452 21420 67508 21422
rect 67788 20860 67844 20916
rect 68012 20860 68068 20916
rect 71036 27074 71092 27076
rect 71036 27022 71038 27074
rect 71038 27022 71090 27074
rect 71090 27022 71092 27074
rect 71036 27020 71092 27022
rect 68572 25394 68628 25396
rect 68572 25342 68574 25394
rect 68574 25342 68626 25394
rect 68626 25342 68628 25394
rect 68572 25340 68628 25342
rect 69020 24834 69076 24836
rect 69020 24782 69022 24834
rect 69022 24782 69074 24834
rect 69074 24782 69076 24834
rect 69020 24780 69076 24782
rect 68832 24330 68888 24332
rect 68832 24278 68834 24330
rect 68834 24278 68886 24330
rect 68886 24278 68888 24330
rect 68832 24276 68888 24278
rect 68936 24330 68992 24332
rect 68936 24278 68938 24330
rect 68938 24278 68990 24330
rect 68990 24278 68992 24330
rect 68936 24276 68992 24278
rect 69040 24330 69096 24332
rect 69040 24278 69042 24330
rect 69042 24278 69094 24330
rect 69094 24278 69096 24330
rect 69040 24276 69096 24278
rect 69916 25394 69972 25396
rect 69916 25342 69918 25394
rect 69918 25342 69970 25394
rect 69970 25342 69972 25394
rect 69916 25340 69972 25342
rect 70588 25340 70644 25396
rect 69804 24834 69860 24836
rect 69804 24782 69806 24834
rect 69806 24782 69858 24834
rect 69858 24782 69860 24834
rect 69804 24780 69860 24782
rect 70700 24780 70756 24836
rect 72268 31388 72324 31444
rect 72156 30156 72212 30212
rect 73388 32508 73444 32564
rect 73500 31276 73556 31332
rect 73388 31164 73444 31220
rect 72380 29148 72436 29204
rect 72716 30044 72772 30100
rect 72716 28588 72772 28644
rect 71372 27244 71428 27300
rect 71260 26236 71316 26292
rect 71932 27074 71988 27076
rect 71932 27022 71934 27074
rect 71934 27022 71986 27074
rect 71986 27022 71988 27074
rect 71932 27020 71988 27022
rect 73052 27298 73108 27300
rect 73052 27246 73054 27298
rect 73054 27246 73106 27298
rect 73106 27246 73108 27298
rect 73052 27244 73108 27246
rect 72492 27074 72548 27076
rect 72492 27022 72494 27074
rect 72494 27022 72546 27074
rect 72546 27022 72548 27074
rect 72492 27020 72548 27022
rect 72044 26012 72100 26068
rect 72268 26908 72324 26964
rect 69244 23884 69300 23940
rect 68572 23154 68628 23156
rect 68572 23102 68574 23154
rect 68574 23102 68626 23154
rect 68626 23102 68628 23154
rect 68572 23100 68628 23102
rect 68832 22762 68888 22764
rect 68832 22710 68834 22762
rect 68834 22710 68886 22762
rect 68886 22710 68888 22762
rect 68832 22708 68888 22710
rect 68936 22762 68992 22764
rect 68936 22710 68938 22762
rect 68938 22710 68990 22762
rect 68990 22710 68992 22762
rect 68936 22708 68992 22710
rect 69040 22762 69096 22764
rect 69040 22710 69042 22762
rect 69042 22710 69094 22762
rect 69094 22710 69096 22762
rect 69040 22708 69096 22710
rect 69244 22428 69300 22484
rect 70588 23042 70644 23044
rect 70588 22990 70590 23042
rect 70590 22990 70642 23042
rect 70642 22990 70644 23042
rect 70588 22988 70644 22990
rect 71260 22988 71316 23044
rect 71148 22540 71204 22596
rect 68348 22258 68404 22260
rect 68348 22206 68350 22258
rect 68350 22206 68402 22258
rect 68402 22206 68404 22258
rect 68348 22204 68404 22206
rect 71372 22652 71428 22708
rect 71484 22540 71540 22596
rect 73500 24556 73556 24612
rect 72604 23436 72660 23492
rect 72156 23324 72212 23380
rect 72156 23154 72212 23156
rect 72156 23102 72158 23154
rect 72158 23102 72210 23154
rect 72210 23102 72212 23154
rect 72156 23100 72212 23102
rect 73612 23436 73668 23492
rect 73500 23378 73556 23380
rect 73500 23326 73502 23378
rect 73502 23326 73554 23378
rect 73554 23326 73556 23378
rect 73500 23324 73556 23326
rect 73276 22988 73332 23044
rect 72492 22482 72548 22484
rect 72492 22430 72494 22482
rect 72494 22430 72546 22482
rect 72546 22430 72548 22482
rect 72492 22428 72548 22430
rect 72940 22370 72996 22372
rect 72940 22318 72942 22370
rect 72942 22318 72994 22370
rect 72994 22318 72996 22370
rect 72940 22316 72996 22318
rect 71036 22092 71092 22148
rect 68832 21194 68888 21196
rect 68832 21142 68834 21194
rect 68834 21142 68886 21194
rect 68886 21142 68888 21194
rect 68832 21140 68888 21142
rect 68936 21194 68992 21196
rect 68936 21142 68938 21194
rect 68938 21142 68990 21194
rect 68990 21142 68992 21194
rect 68936 21140 68992 21142
rect 69040 21194 69096 21196
rect 69040 21142 69042 21194
rect 69042 21142 69094 21194
rect 69094 21142 69096 21194
rect 69040 21140 69096 21142
rect 69244 20860 69300 20916
rect 68236 20690 68292 20692
rect 68236 20638 68238 20690
rect 68238 20638 68290 20690
rect 68290 20638 68292 20690
rect 68236 20636 68292 20638
rect 67004 19852 67060 19908
rect 66780 19234 66836 19236
rect 66780 19182 66782 19234
rect 66782 19182 66834 19234
rect 66834 19182 66836 19234
rect 66780 19180 66836 19182
rect 67900 19906 67956 19908
rect 67900 19854 67902 19906
rect 67902 19854 67954 19906
rect 67954 19854 67956 19906
rect 67900 19852 67956 19854
rect 67564 19122 67620 19124
rect 67564 19070 67566 19122
rect 67566 19070 67618 19122
rect 67618 19070 67620 19122
rect 67564 19068 67620 19070
rect 66668 18338 66724 18340
rect 66668 18286 66670 18338
rect 66670 18286 66722 18338
rect 66722 18286 66724 18338
rect 66668 18284 66724 18286
rect 66332 15372 66388 15428
rect 64092 9042 64148 9044
rect 64092 8990 64094 9042
rect 64094 8990 64146 9042
rect 64146 8990 64148 9042
rect 64092 8988 64148 8990
rect 63756 8316 63812 8372
rect 63868 6860 63924 6916
rect 63756 6636 63812 6692
rect 63756 6188 63812 6244
rect 62188 6018 62244 6020
rect 62188 5966 62190 6018
rect 62190 5966 62242 6018
rect 62242 5966 62244 6018
rect 62188 5964 62244 5966
rect 61068 5740 61124 5796
rect 59500 4172 59556 4228
rect 59164 3948 59220 4004
rect 59948 4508 60004 4564
rect 59836 4450 59892 4452
rect 59836 4398 59838 4450
rect 59838 4398 59890 4450
rect 59890 4398 59892 4450
rect 59836 4396 59892 4398
rect 59724 3836 59780 3892
rect 59612 3778 59668 3780
rect 59612 3726 59614 3778
rect 59614 3726 59666 3778
rect 59666 3726 59668 3778
rect 59612 3724 59668 3726
rect 59500 3554 59556 3556
rect 59500 3502 59502 3554
rect 59502 3502 59554 3554
rect 59554 3502 59556 3554
rect 59500 3500 59556 3502
rect 60396 4450 60452 4452
rect 60396 4398 60398 4450
rect 60398 4398 60450 4450
rect 60450 4398 60452 4450
rect 60396 4396 60452 4398
rect 60396 4172 60452 4228
rect 62972 6018 63028 6020
rect 62972 5966 62974 6018
rect 62974 5966 63026 6018
rect 63026 5966 63028 6018
rect 62972 5964 63028 5966
rect 61068 4508 61124 4564
rect 60732 3836 60788 3892
rect 59948 3500 60004 3556
rect 60172 3500 60228 3556
rect 59612 3330 59668 3332
rect 59612 3278 59614 3330
rect 59614 3278 59666 3330
rect 59666 3278 59668 3330
rect 59612 3276 59668 3278
rect 59172 3162 59228 3164
rect 59172 3110 59174 3162
rect 59174 3110 59226 3162
rect 59226 3110 59228 3162
rect 59172 3108 59228 3110
rect 59276 3162 59332 3164
rect 59276 3110 59278 3162
rect 59278 3110 59330 3162
rect 59330 3110 59332 3162
rect 59276 3108 59332 3110
rect 59380 3162 59436 3164
rect 59380 3110 59382 3162
rect 59382 3110 59434 3162
rect 59434 3110 59436 3162
rect 59380 3108 59436 3110
rect 59052 2940 59108 2996
rect 56924 924 56980 980
rect 60508 3330 60564 3332
rect 60508 3278 60510 3330
rect 60510 3278 60562 3330
rect 60562 3278 60564 3330
rect 60508 3276 60564 3278
rect 62524 5852 62580 5908
rect 62076 5628 62132 5684
rect 61516 4844 61572 4900
rect 61292 4620 61348 4676
rect 61964 5234 62020 5236
rect 61964 5182 61966 5234
rect 61966 5182 62018 5234
rect 62018 5182 62020 5234
rect 61964 5180 62020 5182
rect 61964 4844 62020 4900
rect 61628 4338 61684 4340
rect 61628 4286 61630 4338
rect 61630 4286 61682 4338
rect 61682 4286 61684 4338
rect 61628 4284 61684 4286
rect 62300 4396 62356 4452
rect 61292 3724 61348 3780
rect 61404 3276 61460 3332
rect 61180 2828 61236 2884
rect 63644 5852 63700 5908
rect 63644 5682 63700 5684
rect 63644 5630 63646 5682
rect 63646 5630 63698 5682
rect 63698 5630 63700 5682
rect 63644 5628 63700 5630
rect 66332 14588 66388 14644
rect 65436 9042 65492 9044
rect 65436 8990 65438 9042
rect 65438 8990 65490 9042
rect 65490 8990 65492 9042
rect 65436 8988 65492 8990
rect 65100 8764 65156 8820
rect 65212 8876 65268 8932
rect 64988 8258 65044 8260
rect 64988 8206 64990 8258
rect 64990 8206 65042 8258
rect 65042 8206 65044 8258
rect 64988 8204 65044 8206
rect 64988 7420 65044 7476
rect 64876 7084 64932 7140
rect 64316 6188 64372 6244
rect 63196 4898 63252 4900
rect 63196 4846 63198 4898
rect 63198 4846 63250 4898
rect 63250 4846 63252 4898
rect 63196 4844 63252 4846
rect 63084 4508 63140 4564
rect 63756 4844 63812 4900
rect 63868 4732 63924 4788
rect 63532 4450 63588 4452
rect 63532 4398 63534 4450
rect 63534 4398 63586 4450
rect 63586 4398 63588 4450
rect 63532 4396 63588 4398
rect 63420 4172 63476 4228
rect 64092 4732 64148 4788
rect 64428 5964 64484 6020
rect 64204 4956 64260 5012
rect 63868 4060 63924 4116
rect 63532 3666 63588 3668
rect 63532 3614 63534 3666
rect 63534 3614 63586 3666
rect 63586 3614 63588 3666
rect 63532 3612 63588 3614
rect 64204 3612 64260 3668
rect 64540 6466 64596 6468
rect 64540 6414 64542 6466
rect 64542 6414 64594 6466
rect 64594 6414 64596 6466
rect 64540 6412 64596 6414
rect 62972 3500 63028 3556
rect 64764 6690 64820 6692
rect 64764 6638 64766 6690
rect 64766 6638 64818 6690
rect 64818 6638 64820 6690
rect 64764 6636 64820 6638
rect 64652 5794 64708 5796
rect 64652 5742 64654 5794
rect 64654 5742 64706 5794
rect 64706 5742 64708 5794
rect 64652 5740 64708 5742
rect 64540 4844 64596 4900
rect 64428 4562 64484 4564
rect 64428 4510 64430 4562
rect 64430 4510 64482 4562
rect 64482 4510 64484 4562
rect 64428 4508 64484 4510
rect 65324 8764 65380 8820
rect 65324 8428 65380 8484
rect 65548 7868 65604 7924
rect 65436 7474 65492 7476
rect 65436 7422 65438 7474
rect 65438 7422 65490 7474
rect 65490 7422 65492 7474
rect 65436 7420 65492 7422
rect 65772 8930 65828 8932
rect 65772 8878 65774 8930
rect 65774 8878 65826 8930
rect 65826 8878 65828 8930
rect 65772 8876 65828 8878
rect 65772 8428 65828 8484
rect 66220 12684 66276 12740
rect 65996 12572 66052 12628
rect 65996 10220 66052 10276
rect 67228 18620 67284 18676
rect 68012 18620 68068 18676
rect 68124 18508 68180 18564
rect 67228 17724 67284 17780
rect 66892 16882 66948 16884
rect 66892 16830 66894 16882
rect 66894 16830 66946 16882
rect 66946 16830 66948 16882
rect 66892 16828 66948 16830
rect 67004 14642 67060 14644
rect 67004 14590 67006 14642
rect 67006 14590 67058 14642
rect 67058 14590 67060 14642
rect 67004 14588 67060 14590
rect 66892 14530 66948 14532
rect 66892 14478 66894 14530
rect 66894 14478 66946 14530
rect 66946 14478 66948 14530
rect 66892 14476 66948 14478
rect 66556 13746 66612 13748
rect 66556 13694 66558 13746
rect 66558 13694 66610 13746
rect 66610 13694 66612 13746
rect 66556 13692 66612 13694
rect 66780 12962 66836 12964
rect 66780 12910 66782 12962
rect 66782 12910 66834 12962
rect 66834 12910 66836 12962
rect 66780 12908 66836 12910
rect 66668 12684 66724 12740
rect 66556 12572 66612 12628
rect 66780 12460 66836 12516
rect 66780 12290 66836 12292
rect 66780 12238 66782 12290
rect 66782 12238 66834 12290
rect 66834 12238 66836 12290
rect 66780 12236 66836 12238
rect 66780 11900 66836 11956
rect 66556 11116 66612 11172
rect 66668 11452 66724 11508
rect 66444 9884 66500 9940
rect 66668 9996 66724 10052
rect 66332 8540 66388 8596
rect 66780 9154 66836 9156
rect 66780 9102 66782 9154
rect 66782 9102 66834 9154
rect 66834 9102 66836 9154
rect 66780 9100 66836 9102
rect 66668 8428 66724 8484
rect 66780 8540 66836 8596
rect 67116 14140 67172 14196
rect 67564 16994 67620 16996
rect 67564 16942 67566 16994
rect 67566 16942 67618 16994
rect 67618 16942 67620 16994
rect 67564 16940 67620 16942
rect 67452 16882 67508 16884
rect 67452 16830 67454 16882
rect 67454 16830 67506 16882
rect 67506 16830 67508 16882
rect 67452 16828 67508 16830
rect 67340 16044 67396 16100
rect 67900 15260 67956 15316
rect 67676 14588 67732 14644
rect 68012 14530 68068 14532
rect 68012 14478 68014 14530
rect 68014 14478 68066 14530
rect 68066 14478 68068 14530
rect 68012 14476 68068 14478
rect 67228 14140 67284 14196
rect 67452 14028 67508 14084
rect 67228 13970 67284 13972
rect 67228 13918 67230 13970
rect 67230 13918 67282 13970
rect 67282 13918 67284 13970
rect 67228 13916 67284 13918
rect 67788 13970 67844 13972
rect 67788 13918 67790 13970
rect 67790 13918 67842 13970
rect 67842 13918 67844 13970
rect 67788 13916 67844 13918
rect 68012 13580 68068 13636
rect 67004 13132 67060 13188
rect 67228 13074 67284 13076
rect 67228 13022 67230 13074
rect 67230 13022 67282 13074
rect 67282 13022 67284 13074
rect 67228 13020 67284 13022
rect 67900 12962 67956 12964
rect 67900 12910 67902 12962
rect 67902 12910 67954 12962
rect 67954 12910 67956 12962
rect 67900 12908 67956 12910
rect 67004 12348 67060 12404
rect 67004 11900 67060 11956
rect 67452 11900 67508 11956
rect 67452 11116 67508 11172
rect 67340 10610 67396 10612
rect 67340 10558 67342 10610
rect 67342 10558 67394 10610
rect 67394 10558 67396 10610
rect 67340 10556 67396 10558
rect 67004 10444 67060 10500
rect 67340 10220 67396 10276
rect 66556 7868 66612 7924
rect 66108 7474 66164 7476
rect 66108 7422 66110 7474
rect 66110 7422 66162 7474
rect 66162 7422 66164 7474
rect 66108 7420 66164 7422
rect 65660 7084 65716 7140
rect 65212 6412 65268 6468
rect 64988 6188 65044 6244
rect 65436 5852 65492 5908
rect 66444 6914 66500 6916
rect 66444 6862 66446 6914
rect 66446 6862 66498 6914
rect 66498 6862 66500 6914
rect 66444 6860 66500 6862
rect 65660 6690 65716 6692
rect 65660 6638 65662 6690
rect 65662 6638 65714 6690
rect 65714 6638 65716 6690
rect 65660 6636 65716 6638
rect 65772 6412 65828 6468
rect 64316 2716 64372 2772
rect 65100 4844 65156 4900
rect 65100 1484 65156 1540
rect 65548 5180 65604 5236
rect 65660 5068 65716 5124
rect 66668 6300 66724 6356
rect 66556 6188 66612 6244
rect 66556 6018 66612 6020
rect 66556 5966 66558 6018
rect 66558 5966 66610 6018
rect 66610 5966 66612 6018
rect 66556 5964 66612 5966
rect 65884 5906 65940 5908
rect 65884 5854 65886 5906
rect 65886 5854 65938 5906
rect 65938 5854 65940 5906
rect 65884 5852 65940 5854
rect 65884 5628 65940 5684
rect 66332 5292 66388 5348
rect 66108 5180 66164 5236
rect 65660 3442 65716 3444
rect 65660 3390 65662 3442
rect 65662 3390 65714 3442
rect 65714 3390 65716 3442
rect 65660 3388 65716 3390
rect 66892 5906 66948 5908
rect 66892 5854 66894 5906
rect 66894 5854 66946 5906
rect 66946 5854 66948 5906
rect 66892 5852 66948 5854
rect 67564 10332 67620 10388
rect 69020 20018 69076 20020
rect 69020 19966 69022 20018
rect 69022 19966 69074 20018
rect 69074 19966 69076 20018
rect 69020 19964 69076 19966
rect 68684 19906 68740 19908
rect 68684 19854 68686 19906
rect 68686 19854 68738 19906
rect 68738 19854 68740 19906
rect 68684 19852 68740 19854
rect 68832 19626 68888 19628
rect 68832 19574 68834 19626
rect 68834 19574 68886 19626
rect 68886 19574 68888 19626
rect 68832 19572 68888 19574
rect 68936 19626 68992 19628
rect 68936 19574 68938 19626
rect 68938 19574 68990 19626
rect 68990 19574 68992 19626
rect 68936 19572 68992 19574
rect 69040 19626 69096 19628
rect 69040 19574 69042 19626
rect 69042 19574 69094 19626
rect 69094 19574 69096 19626
rect 69040 19572 69096 19574
rect 68684 18956 68740 19012
rect 68348 18338 68404 18340
rect 68348 18286 68350 18338
rect 68350 18286 68402 18338
rect 68402 18286 68404 18338
rect 68348 18284 68404 18286
rect 68348 17724 68404 17780
rect 68236 14364 68292 14420
rect 68236 14140 68292 14196
rect 68236 13858 68292 13860
rect 68236 13806 68238 13858
rect 68238 13806 68290 13858
rect 68290 13806 68292 13858
rect 68236 13804 68292 13806
rect 68124 13020 68180 13076
rect 68124 12236 68180 12292
rect 68236 12348 68292 12404
rect 68572 10610 68628 10612
rect 68572 10558 68574 10610
rect 68574 10558 68626 10610
rect 68626 10558 68628 10610
rect 68572 10556 68628 10558
rect 68348 10444 68404 10500
rect 68236 10386 68292 10388
rect 68236 10334 68238 10386
rect 68238 10334 68290 10386
rect 68290 10334 68292 10386
rect 68236 10332 68292 10334
rect 68572 10386 68628 10388
rect 68572 10334 68574 10386
rect 68574 10334 68626 10386
rect 68626 10334 68628 10386
rect 68572 10332 68628 10334
rect 67564 9212 67620 9268
rect 67452 9154 67508 9156
rect 67452 9102 67454 9154
rect 67454 9102 67506 9154
rect 67506 9102 67508 9154
rect 67452 9100 67508 9102
rect 67564 8370 67620 8372
rect 67564 8318 67566 8370
rect 67566 8318 67618 8370
rect 67618 8318 67620 8370
rect 67564 8316 67620 8318
rect 67452 7698 67508 7700
rect 67452 7646 67454 7698
rect 67454 7646 67506 7698
rect 67506 7646 67508 7698
rect 67452 7644 67508 7646
rect 67564 7532 67620 7588
rect 67340 7474 67396 7476
rect 67340 7422 67342 7474
rect 67342 7422 67394 7474
rect 67394 7422 67396 7474
rect 67340 7420 67396 7422
rect 67676 7474 67732 7476
rect 67676 7422 67678 7474
rect 67678 7422 67730 7474
rect 67730 7422 67732 7474
rect 67676 7420 67732 7422
rect 67676 7084 67732 7140
rect 68348 9042 68404 9044
rect 68348 8990 68350 9042
rect 68350 8990 68402 9042
rect 68402 8990 68404 9042
rect 68348 8988 68404 8990
rect 67900 7868 67956 7924
rect 68012 8876 68068 8932
rect 68908 18284 68964 18340
rect 69580 20860 69636 20916
rect 69916 21026 69972 21028
rect 69916 20974 69918 21026
rect 69918 20974 69970 21026
rect 69970 20974 69972 21026
rect 69916 20972 69972 20974
rect 70812 20972 70868 21028
rect 69804 20748 69860 20804
rect 69468 20524 69524 20580
rect 69356 19852 69412 19908
rect 69468 20300 69524 20356
rect 70364 20802 70420 20804
rect 70364 20750 70366 20802
rect 70366 20750 70418 20802
rect 70418 20750 70420 20802
rect 70364 20748 70420 20750
rect 69804 20578 69860 20580
rect 69804 20526 69806 20578
rect 69806 20526 69858 20578
rect 69858 20526 69860 20578
rect 69804 20524 69860 20526
rect 69356 19122 69412 19124
rect 69356 19070 69358 19122
rect 69358 19070 69410 19122
rect 69410 19070 69412 19122
rect 69356 19068 69412 19070
rect 69468 19010 69524 19012
rect 69468 18958 69470 19010
rect 69470 18958 69522 19010
rect 69522 18958 69524 19010
rect 69468 18956 69524 18958
rect 68832 18058 68888 18060
rect 68832 18006 68834 18058
rect 68834 18006 68886 18058
rect 68886 18006 68888 18058
rect 68832 18004 68888 18006
rect 68936 18058 68992 18060
rect 68936 18006 68938 18058
rect 68938 18006 68990 18058
rect 68990 18006 68992 18058
rect 68936 18004 68992 18006
rect 69040 18058 69096 18060
rect 69040 18006 69042 18058
rect 69042 18006 69094 18058
rect 69094 18006 69096 18058
rect 69040 18004 69096 18006
rect 68832 16490 68888 16492
rect 68832 16438 68834 16490
rect 68834 16438 68886 16490
rect 68886 16438 68888 16490
rect 68832 16436 68888 16438
rect 68936 16490 68992 16492
rect 68936 16438 68938 16490
rect 68938 16438 68990 16490
rect 68990 16438 68992 16490
rect 68936 16436 68992 16438
rect 69040 16490 69096 16492
rect 69040 16438 69042 16490
rect 69042 16438 69094 16490
rect 69094 16438 69096 16490
rect 69040 16436 69096 16438
rect 70476 20524 70532 20580
rect 69916 19964 69972 20020
rect 70028 20076 70084 20132
rect 69580 18172 69636 18228
rect 69692 19906 69748 19908
rect 69692 19854 69694 19906
rect 69694 19854 69746 19906
rect 69746 19854 69748 19906
rect 69692 19852 69748 19854
rect 70924 20578 70980 20580
rect 70924 20526 70926 20578
rect 70926 20526 70978 20578
rect 70978 20526 70980 20578
rect 70924 20524 70980 20526
rect 71148 20412 71204 20468
rect 70812 19964 70868 20020
rect 70252 19906 70308 19908
rect 70252 19854 70254 19906
rect 70254 19854 70306 19906
rect 70306 19854 70308 19906
rect 70252 19852 70308 19854
rect 70476 19068 70532 19124
rect 70364 18956 70420 19012
rect 70140 18508 70196 18564
rect 70700 18450 70756 18452
rect 70700 18398 70702 18450
rect 70702 18398 70754 18450
rect 70754 18398 70756 18450
rect 70700 18396 70756 18398
rect 69356 17666 69412 17668
rect 69356 17614 69358 17666
rect 69358 17614 69410 17666
rect 69410 17614 69412 17666
rect 69356 17612 69412 17614
rect 69468 16882 69524 16884
rect 69468 16830 69470 16882
rect 69470 16830 69522 16882
rect 69522 16830 69524 16882
rect 69468 16828 69524 16830
rect 69244 15820 69300 15876
rect 69468 16604 69524 16660
rect 68908 15596 68964 15652
rect 69468 15372 69524 15428
rect 68832 14922 68888 14924
rect 68832 14870 68834 14922
rect 68834 14870 68886 14922
rect 68886 14870 68888 14922
rect 68832 14868 68888 14870
rect 68936 14922 68992 14924
rect 68936 14870 68938 14922
rect 68938 14870 68990 14922
rect 68990 14870 68992 14922
rect 68936 14868 68992 14870
rect 69040 14922 69096 14924
rect 69040 14870 69042 14922
rect 69042 14870 69094 14922
rect 69094 14870 69096 14922
rect 69040 14868 69096 14870
rect 69356 13692 69412 13748
rect 68832 13354 68888 13356
rect 68832 13302 68834 13354
rect 68834 13302 68886 13354
rect 68886 13302 68888 13354
rect 68832 13300 68888 13302
rect 68936 13354 68992 13356
rect 68936 13302 68938 13354
rect 68938 13302 68990 13354
rect 68990 13302 68992 13354
rect 68936 13300 68992 13302
rect 69040 13354 69096 13356
rect 69040 13302 69042 13354
rect 69042 13302 69094 13354
rect 69094 13302 69096 13354
rect 69040 13300 69096 13302
rect 68796 12290 68852 12292
rect 68796 12238 68798 12290
rect 68798 12238 68850 12290
rect 68850 12238 68852 12290
rect 68796 12236 68852 12238
rect 69244 12236 69300 12292
rect 68832 11786 68888 11788
rect 68832 11734 68834 11786
rect 68834 11734 68886 11786
rect 68886 11734 68888 11786
rect 68832 11732 68888 11734
rect 68936 11786 68992 11788
rect 68936 11734 68938 11786
rect 68938 11734 68990 11786
rect 68990 11734 68992 11786
rect 68936 11732 68992 11734
rect 69040 11786 69096 11788
rect 69040 11734 69042 11786
rect 69042 11734 69094 11786
rect 69094 11734 69096 11786
rect 69040 11732 69096 11734
rect 69804 17666 69860 17668
rect 69804 17614 69806 17666
rect 69806 17614 69858 17666
rect 69858 17614 69860 17666
rect 69804 17612 69860 17614
rect 69692 17500 69748 17556
rect 70140 17500 70196 17556
rect 70364 17500 70420 17556
rect 70252 17388 70308 17444
rect 69804 16828 69860 16884
rect 69916 15372 69972 15428
rect 69692 14028 69748 14084
rect 69804 13132 69860 13188
rect 69580 12066 69636 12068
rect 69580 12014 69582 12066
rect 69582 12014 69634 12066
rect 69634 12014 69636 12066
rect 69580 12012 69636 12014
rect 70028 15314 70084 15316
rect 70028 15262 70030 15314
rect 70030 15262 70082 15314
rect 70082 15262 70084 15314
rect 70028 15260 70084 15262
rect 71260 20018 71316 20020
rect 71260 19966 71262 20018
rect 71262 19966 71314 20018
rect 71314 19966 71316 20018
rect 71260 19964 71316 19966
rect 73612 23154 73668 23156
rect 73612 23102 73614 23154
rect 73614 23102 73666 23154
rect 73666 23102 73668 23154
rect 73612 23100 73668 23102
rect 73388 22428 73444 22484
rect 73276 21980 73332 22036
rect 72156 21756 72212 21812
rect 71708 21698 71764 21700
rect 71708 21646 71710 21698
rect 71710 21646 71762 21698
rect 71762 21646 71764 21698
rect 71708 21644 71764 21646
rect 74060 34242 74116 34244
rect 74060 34190 74062 34242
rect 74062 34190 74114 34242
rect 74114 34190 74116 34242
rect 74060 34188 74116 34190
rect 73948 33346 74004 33348
rect 73948 33294 73950 33346
rect 73950 33294 74002 33346
rect 74002 33294 74004 33346
rect 73948 33292 74004 33294
rect 74956 34914 75012 34916
rect 74956 34862 74958 34914
rect 74958 34862 75010 34914
rect 75010 34862 75012 34914
rect 74956 34860 75012 34862
rect 74284 32786 74340 32788
rect 74284 32734 74286 32786
rect 74286 32734 74338 32786
rect 74338 32734 74340 32786
rect 74284 32732 74340 32734
rect 74844 33122 74900 33124
rect 74844 33070 74846 33122
rect 74846 33070 74898 33122
rect 74898 33070 74900 33122
rect 74844 33068 74900 33070
rect 74844 32562 74900 32564
rect 74844 32510 74846 32562
rect 74846 32510 74898 32562
rect 74898 32510 74900 32562
rect 74844 32508 74900 32510
rect 73836 28812 73892 28868
rect 73836 26908 73892 26964
rect 73948 26572 74004 26628
rect 74396 31500 74452 31556
rect 74620 31218 74676 31220
rect 74620 31166 74622 31218
rect 74622 31166 74674 31218
rect 74674 31166 74676 31218
rect 74620 31164 74676 31166
rect 74396 30322 74452 30324
rect 74396 30270 74398 30322
rect 74398 30270 74450 30322
rect 74450 30270 74452 30322
rect 74396 30268 74452 30270
rect 74172 29932 74228 29988
rect 74284 29820 74340 29876
rect 75068 30210 75124 30212
rect 75068 30158 75070 30210
rect 75070 30158 75122 30210
rect 75122 30158 75124 30210
rect 75068 30156 75124 30158
rect 74956 30044 75012 30100
rect 74508 28812 74564 28868
rect 74844 29820 74900 29876
rect 74508 27916 74564 27972
rect 74172 27804 74228 27860
rect 74508 27468 74564 27524
rect 75068 29708 75124 29764
rect 75740 35980 75796 36036
rect 75628 33458 75684 33460
rect 75628 33406 75630 33458
rect 75630 33406 75682 33458
rect 75682 33406 75684 33458
rect 75628 33404 75684 33406
rect 76300 35980 76356 36036
rect 76076 35868 76132 35924
rect 76748 35756 76804 35812
rect 76076 35026 76132 35028
rect 76076 34974 76078 35026
rect 76078 34974 76130 35026
rect 76130 34974 76132 35026
rect 76076 34972 76132 34974
rect 77980 36594 78036 36596
rect 77980 36542 77982 36594
rect 77982 36542 78034 36594
rect 78034 36542 78036 36594
rect 77980 36540 78036 36542
rect 77532 35196 77588 35252
rect 77084 34748 77140 34804
rect 76748 34242 76804 34244
rect 76748 34190 76750 34242
rect 76750 34190 76802 34242
rect 76802 34190 76804 34242
rect 76748 34188 76804 34190
rect 76076 33628 76132 33684
rect 76412 33404 76468 33460
rect 77980 35084 78036 35140
rect 77532 34076 77588 34132
rect 77308 33292 77364 33348
rect 75740 32732 75796 32788
rect 75404 31500 75460 31556
rect 76300 31164 76356 31220
rect 75516 31052 75572 31108
rect 75964 30716 76020 30772
rect 75404 30322 75460 30324
rect 75404 30270 75406 30322
rect 75406 30270 75458 30322
rect 75458 30270 75460 30322
rect 75404 30268 75460 30270
rect 75516 30210 75572 30212
rect 75516 30158 75518 30210
rect 75518 30158 75570 30210
rect 75570 30158 75572 30210
rect 75516 30156 75572 30158
rect 76076 30156 76132 30212
rect 76188 29820 76244 29876
rect 75516 28700 75572 28756
rect 75404 28642 75460 28644
rect 75404 28590 75406 28642
rect 75406 28590 75458 28642
rect 75458 28590 75460 28642
rect 75404 28588 75460 28590
rect 76076 28588 76132 28644
rect 76300 28700 76356 28756
rect 76636 31836 76692 31892
rect 77084 30994 77140 30996
rect 77084 30942 77086 30994
rect 77086 30942 77138 30994
rect 77138 30942 77140 30994
rect 77084 30940 77140 30942
rect 76524 30044 76580 30100
rect 76188 28140 76244 28196
rect 75740 27970 75796 27972
rect 75740 27918 75742 27970
rect 75742 27918 75794 27970
rect 75794 27918 75796 27970
rect 75740 27916 75796 27918
rect 75628 27468 75684 27524
rect 76188 27132 76244 27188
rect 74172 26572 74228 26628
rect 74284 26514 74340 26516
rect 74284 26462 74286 26514
rect 74286 26462 74338 26514
rect 74338 26462 74340 26514
rect 74284 26460 74340 26462
rect 74172 26290 74228 26292
rect 74172 26238 74174 26290
rect 74174 26238 74226 26290
rect 74226 26238 74228 26290
rect 74172 26236 74228 26238
rect 74284 26012 74340 26068
rect 74396 25900 74452 25956
rect 74060 24610 74116 24612
rect 74060 24558 74062 24610
rect 74062 24558 74114 24610
rect 74114 24558 74116 24610
rect 74060 24556 74116 24558
rect 73948 22540 74004 22596
rect 73724 21532 73780 21588
rect 72716 20914 72772 20916
rect 72716 20862 72718 20914
rect 72718 20862 72770 20914
rect 72770 20862 72772 20914
rect 72716 20860 72772 20862
rect 74396 22204 74452 22260
rect 74396 21586 74452 21588
rect 74396 21534 74398 21586
rect 74398 21534 74450 21586
rect 74450 21534 74452 21586
rect 74396 21532 74452 21534
rect 74172 20972 74228 21028
rect 73724 20802 73780 20804
rect 73724 20750 73726 20802
rect 73726 20750 73778 20802
rect 73778 20750 73780 20802
rect 73724 20748 73780 20750
rect 71596 20300 71652 20356
rect 71708 20636 71764 20692
rect 72268 20690 72324 20692
rect 72268 20638 72270 20690
rect 72270 20638 72322 20690
rect 72322 20638 72324 20690
rect 72268 20636 72324 20638
rect 72044 19964 72100 20020
rect 71932 19906 71988 19908
rect 71932 19854 71934 19906
rect 71934 19854 71986 19906
rect 71986 19854 71988 19906
rect 71932 19852 71988 19854
rect 72492 19852 72548 19908
rect 72044 19740 72100 19796
rect 71708 19010 71764 19012
rect 71708 18958 71710 19010
rect 71710 18958 71762 19010
rect 71762 18958 71764 19010
rect 71708 18956 71764 18958
rect 71372 18508 71428 18564
rect 71260 17666 71316 17668
rect 71260 17614 71262 17666
rect 71262 17614 71314 17666
rect 71314 17614 71316 17666
rect 71260 17612 71316 17614
rect 72156 18450 72212 18452
rect 72156 18398 72158 18450
rect 72158 18398 72210 18450
rect 72210 18398 72212 18450
rect 72156 18396 72212 18398
rect 71036 17554 71092 17556
rect 71036 17502 71038 17554
rect 71038 17502 71090 17554
rect 71090 17502 71092 17554
rect 71036 17500 71092 17502
rect 71484 17388 71540 17444
rect 70924 15596 70980 15652
rect 71036 15538 71092 15540
rect 71036 15486 71038 15538
rect 71038 15486 71090 15538
rect 71090 15486 71092 15538
rect 71036 15484 71092 15486
rect 71596 15426 71652 15428
rect 71596 15374 71598 15426
rect 71598 15374 71650 15426
rect 71650 15374 71652 15426
rect 71596 15372 71652 15374
rect 70364 15036 70420 15092
rect 70028 14700 70084 14756
rect 71260 14700 71316 14756
rect 71820 14700 71876 14756
rect 70476 14530 70532 14532
rect 70476 14478 70478 14530
rect 70478 14478 70530 14530
rect 70530 14478 70532 14530
rect 70476 14476 70532 14478
rect 71484 14530 71540 14532
rect 71484 14478 71486 14530
rect 71486 14478 71538 14530
rect 71538 14478 71540 14530
rect 71484 14476 71540 14478
rect 70140 13804 70196 13860
rect 70364 13634 70420 13636
rect 70364 13582 70366 13634
rect 70366 13582 70418 13634
rect 70418 13582 70420 13634
rect 70364 13580 70420 13582
rect 70812 13634 70868 13636
rect 70812 13582 70814 13634
rect 70814 13582 70866 13634
rect 70866 13582 70868 13634
rect 70812 13580 70868 13582
rect 71708 13804 71764 13860
rect 71484 13746 71540 13748
rect 71484 13694 71486 13746
rect 71486 13694 71538 13746
rect 71538 13694 71540 13746
rect 71484 13692 71540 13694
rect 71372 13634 71428 13636
rect 71372 13582 71374 13634
rect 71374 13582 71426 13634
rect 71426 13582 71428 13634
rect 71372 13580 71428 13582
rect 70140 12850 70196 12852
rect 70140 12798 70142 12850
rect 70142 12798 70194 12850
rect 70194 12798 70196 12850
rect 70140 12796 70196 12798
rect 70252 13132 70308 13188
rect 70476 12738 70532 12740
rect 70476 12686 70478 12738
rect 70478 12686 70530 12738
rect 70530 12686 70532 12738
rect 70476 12684 70532 12686
rect 71148 12684 71204 12740
rect 70028 12012 70084 12068
rect 70364 12066 70420 12068
rect 70364 12014 70366 12066
rect 70366 12014 70418 12066
rect 70418 12014 70420 12066
rect 70364 12012 70420 12014
rect 70140 11394 70196 11396
rect 70140 11342 70142 11394
rect 70142 11342 70194 11394
rect 70194 11342 70196 11394
rect 70140 11340 70196 11342
rect 69356 11004 69412 11060
rect 69356 10834 69412 10836
rect 69356 10782 69358 10834
rect 69358 10782 69410 10834
rect 69410 10782 69412 10834
rect 69356 10780 69412 10782
rect 69244 10386 69300 10388
rect 69244 10334 69246 10386
rect 69246 10334 69298 10386
rect 69298 10334 69300 10386
rect 69244 10332 69300 10334
rect 68832 10218 68888 10220
rect 68832 10166 68834 10218
rect 68834 10166 68886 10218
rect 68886 10166 68888 10218
rect 68832 10164 68888 10166
rect 68936 10218 68992 10220
rect 68936 10166 68938 10218
rect 68938 10166 68990 10218
rect 68990 10166 68992 10218
rect 68936 10164 68992 10166
rect 69040 10218 69096 10220
rect 69040 10166 69042 10218
rect 69042 10166 69094 10218
rect 69094 10166 69096 10218
rect 69040 10164 69096 10166
rect 69692 9826 69748 9828
rect 69692 9774 69694 9826
rect 69694 9774 69746 9826
rect 69746 9774 69748 9826
rect 69692 9772 69748 9774
rect 69020 9660 69076 9716
rect 68908 9436 68964 9492
rect 70140 11004 70196 11060
rect 72044 14476 72100 14532
rect 73276 19740 73332 19796
rect 73836 19740 73892 19796
rect 73836 19292 73892 19348
rect 73948 20524 74004 20580
rect 73724 18508 73780 18564
rect 73836 18284 73892 18340
rect 74060 19740 74116 19796
rect 74732 26572 74788 26628
rect 74956 25676 75012 25732
rect 75068 26236 75124 26292
rect 74844 25116 74900 25172
rect 75628 26236 75684 26292
rect 75516 26178 75572 26180
rect 75516 26126 75518 26178
rect 75518 26126 75570 26178
rect 75570 26126 75572 26178
rect 75516 26124 75572 26126
rect 75964 26962 76020 26964
rect 75964 26910 75966 26962
rect 75966 26910 76018 26962
rect 76018 26910 76020 26962
rect 75964 26908 76020 26910
rect 75852 25900 75908 25956
rect 75852 25116 75908 25172
rect 76524 28140 76580 28196
rect 76972 28924 77028 28980
rect 76748 27970 76804 27972
rect 76748 27918 76750 27970
rect 76750 27918 76802 27970
rect 76802 27918 76804 27970
rect 76748 27916 76804 27918
rect 76972 27858 77028 27860
rect 76972 27806 76974 27858
rect 76974 27806 77026 27858
rect 77026 27806 77028 27858
rect 76972 27804 77028 27806
rect 76412 27468 76468 27524
rect 76412 27298 76468 27300
rect 76412 27246 76414 27298
rect 76414 27246 76466 27298
rect 76466 27246 76468 27298
rect 76412 27244 76468 27246
rect 76972 27020 77028 27076
rect 76524 25618 76580 25620
rect 76524 25566 76526 25618
rect 76526 25566 76578 25618
rect 76578 25566 76580 25618
rect 76524 25564 76580 25566
rect 75852 24780 75908 24836
rect 75292 24722 75348 24724
rect 75292 24670 75294 24722
rect 75294 24670 75346 24722
rect 75346 24670 75348 24722
rect 75292 24668 75348 24670
rect 75180 24556 75236 24612
rect 75516 23660 75572 23716
rect 75628 23436 75684 23492
rect 75740 22988 75796 23044
rect 75628 22370 75684 22372
rect 75628 22318 75630 22370
rect 75630 22318 75682 22370
rect 75682 22318 75684 22370
rect 75628 22316 75684 22318
rect 74732 22092 74788 22148
rect 74620 21644 74676 21700
rect 75404 22258 75460 22260
rect 75404 22206 75406 22258
rect 75406 22206 75458 22258
rect 75458 22206 75460 22258
rect 75404 22204 75460 22206
rect 75852 21756 75908 21812
rect 74956 21586 75012 21588
rect 74956 21534 74958 21586
rect 74958 21534 75010 21586
rect 75010 21534 75012 21586
rect 74956 21532 75012 21534
rect 74844 20860 74900 20916
rect 75068 20972 75124 21028
rect 74620 20076 74676 20132
rect 74284 19852 74340 19908
rect 74396 19964 74452 20020
rect 74172 19628 74228 19684
rect 74396 19346 74452 19348
rect 74396 19294 74398 19346
rect 74398 19294 74450 19346
rect 74450 19294 74452 19346
rect 74396 19292 74452 19294
rect 74060 18226 74116 18228
rect 74060 18174 74062 18226
rect 74062 18174 74114 18226
rect 74114 18174 74116 18226
rect 74060 18172 74116 18174
rect 73948 17554 74004 17556
rect 73948 17502 73950 17554
rect 73950 17502 74002 17554
rect 74002 17502 74004 17554
rect 73948 17500 74004 17502
rect 72268 15372 72324 15428
rect 73276 16098 73332 16100
rect 73276 16046 73278 16098
rect 73278 16046 73330 16098
rect 73330 16046 73332 16098
rect 73276 16044 73332 16046
rect 73500 15426 73556 15428
rect 73500 15374 73502 15426
rect 73502 15374 73554 15426
rect 73554 15374 73556 15426
rect 73500 15372 73556 15374
rect 74732 19852 74788 19908
rect 74620 18450 74676 18452
rect 74620 18398 74622 18450
rect 74622 18398 74674 18450
rect 74674 18398 74676 18450
rect 74620 18396 74676 18398
rect 74620 17666 74676 17668
rect 74620 17614 74622 17666
rect 74622 17614 74674 17666
rect 74674 17614 74676 17666
rect 74620 17612 74676 17614
rect 74508 17554 74564 17556
rect 74508 17502 74510 17554
rect 74510 17502 74562 17554
rect 74562 17502 74564 17554
rect 74508 17500 74564 17502
rect 73948 16044 74004 16100
rect 74060 15426 74116 15428
rect 74060 15374 74062 15426
rect 74062 15374 74114 15426
rect 74114 15374 74116 15426
rect 74060 15372 74116 15374
rect 72380 14642 72436 14644
rect 72380 14590 72382 14642
rect 72382 14590 72434 14642
rect 72434 14590 72436 14642
rect 72380 14588 72436 14590
rect 73052 14642 73108 14644
rect 73052 14590 73054 14642
rect 73054 14590 73106 14642
rect 73106 14590 73108 14642
rect 73052 14588 73108 14590
rect 72268 13746 72324 13748
rect 72268 13694 72270 13746
rect 72270 13694 72322 13746
rect 72322 13694 72324 13746
rect 72268 13692 72324 13694
rect 72380 12796 72436 12852
rect 70812 11340 70868 11396
rect 71036 11004 71092 11060
rect 70028 9660 70084 9716
rect 69468 9436 69524 9492
rect 70028 9436 70084 9492
rect 69020 9100 69076 9156
rect 69132 9042 69188 9044
rect 69132 8990 69134 9042
rect 69134 8990 69186 9042
rect 69186 8990 69188 9042
rect 69132 8988 69188 8990
rect 68832 8650 68888 8652
rect 68832 8598 68834 8650
rect 68834 8598 68886 8650
rect 68886 8598 68888 8650
rect 68832 8596 68888 8598
rect 68936 8650 68992 8652
rect 68936 8598 68938 8650
rect 68938 8598 68990 8650
rect 68990 8598 68992 8650
rect 68936 8596 68992 8598
rect 69040 8650 69096 8652
rect 69040 8598 69042 8650
rect 69042 8598 69094 8650
rect 69094 8598 69096 8650
rect 69040 8596 69096 8598
rect 69580 9266 69636 9268
rect 69580 9214 69582 9266
rect 69582 9214 69634 9266
rect 69634 9214 69636 9266
rect 69580 9212 69636 9214
rect 68124 7586 68180 7588
rect 68124 7534 68126 7586
rect 68126 7534 68178 7586
rect 68178 7534 68180 7586
rect 68124 7532 68180 7534
rect 67900 6466 67956 6468
rect 67900 6414 67902 6466
rect 67902 6414 67954 6466
rect 67954 6414 67956 6466
rect 67900 6412 67956 6414
rect 67676 6300 67732 6356
rect 67116 5964 67172 6020
rect 67228 6076 67284 6132
rect 67452 5964 67508 6020
rect 68124 5906 68180 5908
rect 68124 5854 68126 5906
rect 68126 5854 68178 5906
rect 68178 5854 68180 5906
rect 68124 5852 68180 5854
rect 67228 5628 67284 5684
rect 67004 5292 67060 5348
rect 66668 5180 66724 5236
rect 66556 5122 66612 5124
rect 66556 5070 66558 5122
rect 66558 5070 66610 5122
rect 66610 5070 66612 5122
rect 66556 5068 66612 5070
rect 67676 4956 67732 5012
rect 66332 4898 66388 4900
rect 66332 4846 66334 4898
rect 66334 4846 66386 4898
rect 66386 4846 66388 4898
rect 66332 4844 66388 4846
rect 66556 4844 66612 4900
rect 66220 4732 66276 4788
rect 66892 4508 66948 4564
rect 67004 4732 67060 4788
rect 65436 1372 65492 1428
rect 67116 4620 67172 4676
rect 67340 4284 67396 4340
rect 67676 4114 67732 4116
rect 67676 4062 67678 4114
rect 67678 4062 67730 4114
rect 67730 4062 67732 4114
rect 67676 4060 67732 4062
rect 67340 3836 67396 3892
rect 68460 7868 68516 7924
rect 68460 7698 68516 7700
rect 68460 7646 68462 7698
rect 68462 7646 68514 7698
rect 68514 7646 68516 7698
rect 68460 7644 68516 7646
rect 69356 7474 69412 7476
rect 69356 7422 69358 7474
rect 69358 7422 69410 7474
rect 69410 7422 69412 7474
rect 69356 7420 69412 7422
rect 68348 6690 68404 6692
rect 68348 6638 68350 6690
rect 68350 6638 68402 6690
rect 68402 6638 68404 6690
rect 68348 6636 68404 6638
rect 68124 4732 68180 4788
rect 68124 4508 68180 4564
rect 68348 4732 68404 4788
rect 68236 4450 68292 4452
rect 68236 4398 68238 4450
rect 68238 4398 68290 4450
rect 68290 4398 68292 4450
rect 68236 4396 68292 4398
rect 68348 4172 68404 4228
rect 68832 7082 68888 7084
rect 68832 7030 68834 7082
rect 68834 7030 68886 7082
rect 68886 7030 68888 7082
rect 68832 7028 68888 7030
rect 68936 7082 68992 7084
rect 68936 7030 68938 7082
rect 68938 7030 68990 7082
rect 68990 7030 68992 7082
rect 68936 7028 68992 7030
rect 69040 7082 69096 7084
rect 69040 7030 69042 7082
rect 69042 7030 69094 7082
rect 69094 7030 69096 7082
rect 69040 7028 69096 7030
rect 68572 6636 68628 6692
rect 68908 6412 68964 6468
rect 70588 9826 70644 9828
rect 70588 9774 70590 9826
rect 70590 9774 70642 9826
rect 70642 9774 70644 9826
rect 70588 9772 70644 9774
rect 70252 9212 70308 9268
rect 70364 8988 70420 9044
rect 69804 8876 69860 8932
rect 69692 8204 69748 8260
rect 70476 8930 70532 8932
rect 70476 8878 70478 8930
rect 70478 8878 70530 8930
rect 70530 8878 70532 8930
rect 70476 8876 70532 8878
rect 71148 9714 71204 9716
rect 71148 9662 71150 9714
rect 71150 9662 71202 9714
rect 71202 9662 71204 9714
rect 71148 9660 71204 9662
rect 70924 8876 70980 8932
rect 72380 11900 72436 11956
rect 72268 11004 72324 11060
rect 72492 10498 72548 10500
rect 72492 10446 72494 10498
rect 72494 10446 72546 10498
rect 72546 10446 72548 10498
rect 72492 10444 72548 10446
rect 72156 9772 72212 9828
rect 69804 8146 69860 8148
rect 69804 8094 69806 8146
rect 69806 8094 69858 8146
rect 69858 8094 69860 8146
rect 69804 8092 69860 8094
rect 70364 8146 70420 8148
rect 70364 8094 70366 8146
rect 70366 8094 70418 8146
rect 70418 8094 70420 8146
rect 70364 8092 70420 8094
rect 71148 8092 71204 8148
rect 72268 9266 72324 9268
rect 72268 9214 72270 9266
rect 72270 9214 72322 9266
rect 72322 9214 72324 9266
rect 72268 9212 72324 9214
rect 71596 9042 71652 9044
rect 71596 8990 71598 9042
rect 71598 8990 71650 9042
rect 71650 8990 71652 9042
rect 71596 8988 71652 8990
rect 71932 9042 71988 9044
rect 71932 8990 71934 9042
rect 71934 8990 71986 9042
rect 71986 8990 71988 9042
rect 71932 8988 71988 8990
rect 69692 7756 69748 7812
rect 69916 7698 69972 7700
rect 69916 7646 69918 7698
rect 69918 7646 69970 7698
rect 69970 7646 69972 7698
rect 69916 7644 69972 7646
rect 72044 8258 72100 8260
rect 72044 8206 72046 8258
rect 72046 8206 72098 8258
rect 72098 8206 72100 8258
rect 72044 8204 72100 8206
rect 71372 7644 71428 7700
rect 70588 7586 70644 7588
rect 70588 7534 70590 7586
rect 70590 7534 70642 7586
rect 70642 7534 70644 7586
rect 70588 7532 70644 7534
rect 69580 7362 69636 7364
rect 69580 7310 69582 7362
rect 69582 7310 69634 7362
rect 69634 7310 69636 7362
rect 69580 7308 69636 7310
rect 69580 6860 69636 6916
rect 69468 6412 69524 6468
rect 71708 7474 71764 7476
rect 71708 7422 71710 7474
rect 71710 7422 71762 7474
rect 71762 7422 71764 7474
rect 71708 7420 71764 7422
rect 71820 7362 71876 7364
rect 71820 7310 71822 7362
rect 71822 7310 71874 7362
rect 71874 7310 71876 7362
rect 71820 7308 71876 7310
rect 70028 6690 70084 6692
rect 70028 6638 70030 6690
rect 70030 6638 70082 6690
rect 70082 6638 70084 6690
rect 70028 6636 70084 6638
rect 70924 6690 70980 6692
rect 70924 6638 70926 6690
rect 70926 6638 70978 6690
rect 70978 6638 70980 6690
rect 70924 6636 70980 6638
rect 70252 6524 70308 6580
rect 69804 6130 69860 6132
rect 69804 6078 69806 6130
rect 69806 6078 69858 6130
rect 69858 6078 69860 6130
rect 69804 6076 69860 6078
rect 70700 6300 70756 6356
rect 70588 6076 70644 6132
rect 69692 5852 69748 5908
rect 68796 5628 68852 5684
rect 69356 5794 69412 5796
rect 69356 5742 69358 5794
rect 69358 5742 69410 5794
rect 69410 5742 69412 5794
rect 69356 5740 69412 5742
rect 68832 5514 68888 5516
rect 68832 5462 68834 5514
rect 68834 5462 68886 5514
rect 68886 5462 68888 5514
rect 68832 5460 68888 5462
rect 68936 5514 68992 5516
rect 68936 5462 68938 5514
rect 68938 5462 68990 5514
rect 68990 5462 68992 5514
rect 68936 5460 68992 5462
rect 69040 5514 69096 5516
rect 69040 5462 69042 5514
rect 69042 5462 69094 5514
rect 69094 5462 69096 5514
rect 69040 5460 69096 5462
rect 69692 5234 69748 5236
rect 69692 5182 69694 5234
rect 69694 5182 69746 5234
rect 69746 5182 69748 5234
rect 69692 5180 69748 5182
rect 70924 5964 70980 6020
rect 71036 6412 71092 6468
rect 69132 4956 69188 5012
rect 69580 4620 69636 4676
rect 70252 4508 70308 4564
rect 69580 4396 69636 4452
rect 70924 4338 70980 4340
rect 70924 4286 70926 4338
rect 70926 4286 70978 4338
rect 70978 4286 70980 4338
rect 70924 4284 70980 4286
rect 68832 3946 68888 3948
rect 68832 3894 68834 3946
rect 68834 3894 68886 3946
rect 68886 3894 68888 3946
rect 68832 3892 68888 3894
rect 68936 3946 68992 3948
rect 68936 3894 68938 3946
rect 68938 3894 68990 3946
rect 68990 3894 68992 3946
rect 68936 3892 68992 3894
rect 69040 3946 69096 3948
rect 69040 3894 69042 3946
rect 69042 3894 69094 3946
rect 69094 3894 69096 3946
rect 69040 3892 69096 3894
rect 70252 3612 70308 3668
rect 68348 3554 68404 3556
rect 68348 3502 68350 3554
rect 68350 3502 68402 3554
rect 68402 3502 68404 3554
rect 68348 3500 68404 3502
rect 67004 2940 67060 2996
rect 68684 3388 68740 3444
rect 70252 3442 70308 3444
rect 70252 3390 70254 3442
rect 70254 3390 70306 3442
rect 70306 3390 70308 3442
rect 70252 3388 70308 3390
rect 70812 3388 70868 3444
rect 71484 6466 71540 6468
rect 71484 6414 71486 6466
rect 71486 6414 71538 6466
rect 71538 6414 71540 6466
rect 71484 6412 71540 6414
rect 72044 5906 72100 5908
rect 72044 5854 72046 5906
rect 72046 5854 72098 5906
rect 72098 5854 72100 5906
rect 72044 5852 72100 5854
rect 72044 5516 72100 5572
rect 71372 3442 71428 3444
rect 71372 3390 71374 3442
rect 71374 3390 71426 3442
rect 71426 3390 71428 3442
rect 71372 3388 71428 3390
rect 73500 13858 73556 13860
rect 73500 13806 73502 13858
rect 73502 13806 73554 13858
rect 73554 13806 73556 13858
rect 73500 13804 73556 13806
rect 74844 16098 74900 16100
rect 74844 16046 74846 16098
rect 74846 16046 74898 16098
rect 74898 16046 74900 16098
rect 74844 16044 74900 16046
rect 74508 15426 74564 15428
rect 74508 15374 74510 15426
rect 74510 15374 74562 15426
rect 74562 15374 74564 15426
rect 74508 15372 74564 15374
rect 75516 20914 75572 20916
rect 75516 20862 75518 20914
rect 75518 20862 75570 20914
rect 75570 20862 75572 20914
rect 75516 20860 75572 20862
rect 75180 20524 75236 20580
rect 75292 20018 75348 20020
rect 75292 19966 75294 20018
rect 75294 19966 75346 20018
rect 75346 19966 75348 20018
rect 75292 19964 75348 19966
rect 75404 19906 75460 19908
rect 75404 19854 75406 19906
rect 75406 19854 75458 19906
rect 75458 19854 75460 19906
rect 75404 19852 75460 19854
rect 75628 19794 75684 19796
rect 75628 19742 75630 19794
rect 75630 19742 75682 19794
rect 75682 19742 75684 19794
rect 75628 19740 75684 19742
rect 75516 18956 75572 19012
rect 75180 18172 75236 18228
rect 75180 17778 75236 17780
rect 75180 17726 75182 17778
rect 75182 17726 75234 17778
rect 75234 17726 75236 17778
rect 75180 17724 75236 17726
rect 75628 17500 75684 17556
rect 75180 17388 75236 17444
rect 75516 17388 75572 17444
rect 75292 16492 75348 16548
rect 75180 15260 75236 15316
rect 74620 14364 74676 14420
rect 73500 12402 73556 12404
rect 73500 12350 73502 12402
rect 73502 12350 73554 12402
rect 73554 12350 73556 12402
rect 73500 12348 73556 12350
rect 73388 11340 73444 11396
rect 73388 10498 73444 10500
rect 73388 10446 73390 10498
rect 73390 10446 73442 10498
rect 73442 10446 73444 10498
rect 73388 10444 73444 10446
rect 74060 12402 74116 12404
rect 74060 12350 74062 12402
rect 74062 12350 74114 12402
rect 74114 12350 74116 12402
rect 74060 12348 74116 12350
rect 73836 11394 73892 11396
rect 73836 11342 73838 11394
rect 73838 11342 73890 11394
rect 73890 11342 73892 11394
rect 73836 11340 73892 11342
rect 73724 10610 73780 10612
rect 73724 10558 73726 10610
rect 73726 10558 73778 10610
rect 73778 10558 73780 10610
rect 73724 10556 73780 10558
rect 73052 8876 73108 8932
rect 72716 8258 72772 8260
rect 72716 8206 72718 8258
rect 72718 8206 72770 8258
rect 72770 8206 72772 8258
rect 72716 8204 72772 8206
rect 72268 6524 72324 6580
rect 72380 6412 72436 6468
rect 72716 6466 72772 6468
rect 72716 6414 72718 6466
rect 72718 6414 72770 6466
rect 72770 6414 72772 6466
rect 72716 6412 72772 6414
rect 72492 5852 72548 5908
rect 73724 9714 73780 9716
rect 73724 9662 73726 9714
rect 73726 9662 73778 9714
rect 73778 9662 73780 9714
rect 73724 9660 73780 9662
rect 73948 9042 74004 9044
rect 73948 8990 73950 9042
rect 73950 8990 74002 9042
rect 74002 8990 74004 9042
rect 73948 8988 74004 8990
rect 74508 10332 74564 10388
rect 75404 16156 75460 16212
rect 76860 24834 76916 24836
rect 76860 24782 76862 24834
rect 76862 24782 76914 24834
rect 76914 24782 76916 24834
rect 76860 24780 76916 24782
rect 76300 24556 76356 24612
rect 76412 24668 76468 24724
rect 76188 23938 76244 23940
rect 76188 23886 76190 23938
rect 76190 23886 76242 23938
rect 76242 23886 76244 23938
rect 76188 23884 76244 23886
rect 76860 23042 76916 23044
rect 76860 22990 76862 23042
rect 76862 22990 76914 23042
rect 76914 22990 76916 23042
rect 76860 22988 76916 22990
rect 76748 22316 76804 22372
rect 77084 22092 77140 22148
rect 76860 21810 76916 21812
rect 76860 21758 76862 21810
rect 76862 21758 76914 21810
rect 76914 21758 76916 21810
rect 76860 21756 76916 21758
rect 76076 21196 76132 21252
rect 76972 20130 77028 20132
rect 76972 20078 76974 20130
rect 76974 20078 77026 20130
rect 77026 20078 77028 20130
rect 76972 20076 77028 20078
rect 77084 19740 77140 19796
rect 76636 19628 76692 19684
rect 76188 19234 76244 19236
rect 76188 19182 76190 19234
rect 76190 19182 76242 19234
rect 76242 19182 76244 19234
rect 76188 19180 76244 19182
rect 77532 32844 77588 32900
rect 77532 32674 77588 32676
rect 77532 32622 77534 32674
rect 77534 32622 77586 32674
rect 77586 32622 77588 32674
rect 77532 32620 77588 32622
rect 77308 31890 77364 31892
rect 77308 31838 77310 31890
rect 77310 31838 77362 31890
rect 77362 31838 77364 31890
rect 77308 31836 77364 31838
rect 77532 31724 77588 31780
rect 77420 31666 77476 31668
rect 77420 31614 77422 31666
rect 77422 31614 77474 31666
rect 77474 31614 77476 31666
rect 77420 31612 77476 31614
rect 77532 31554 77588 31556
rect 77532 31502 77534 31554
rect 77534 31502 77586 31554
rect 77586 31502 77588 31554
rect 77532 31500 77588 31502
rect 78492 36090 78548 36092
rect 78492 36038 78494 36090
rect 78494 36038 78546 36090
rect 78546 36038 78548 36090
rect 78492 36036 78548 36038
rect 78596 36090 78652 36092
rect 78596 36038 78598 36090
rect 78598 36038 78650 36090
rect 78650 36038 78652 36090
rect 78596 36036 78652 36038
rect 78700 36090 78756 36092
rect 78700 36038 78702 36090
rect 78702 36038 78754 36090
rect 78754 36038 78756 36090
rect 78700 36036 78756 36038
rect 78092 34972 78148 35028
rect 78092 34802 78148 34804
rect 78092 34750 78094 34802
rect 78094 34750 78146 34802
rect 78146 34750 78148 34802
rect 78092 34748 78148 34750
rect 78492 34522 78548 34524
rect 78492 34470 78494 34522
rect 78494 34470 78546 34522
rect 78546 34470 78548 34522
rect 78492 34468 78548 34470
rect 78596 34522 78652 34524
rect 78596 34470 78598 34522
rect 78598 34470 78650 34522
rect 78650 34470 78652 34522
rect 78596 34468 78652 34470
rect 78700 34522 78756 34524
rect 78700 34470 78702 34522
rect 78702 34470 78754 34522
rect 78754 34470 78756 34522
rect 78700 34468 78756 34470
rect 77980 34130 78036 34132
rect 77980 34078 77982 34130
rect 77982 34078 78034 34130
rect 78034 34078 78036 34130
rect 77980 34076 78036 34078
rect 78876 34188 78932 34244
rect 78204 34076 78260 34132
rect 78092 32844 78148 32900
rect 77980 32674 78036 32676
rect 77980 32622 77982 32674
rect 77982 32622 78034 32674
rect 78034 32622 78036 32674
rect 77980 32620 78036 32622
rect 78492 32954 78548 32956
rect 78492 32902 78494 32954
rect 78494 32902 78546 32954
rect 78546 32902 78548 32954
rect 78492 32900 78548 32902
rect 78596 32954 78652 32956
rect 78596 32902 78598 32954
rect 78598 32902 78650 32954
rect 78650 32902 78652 32954
rect 78596 32900 78652 32902
rect 78700 32954 78756 32956
rect 78700 32902 78702 32954
rect 78702 32902 78754 32954
rect 78754 32902 78756 32954
rect 78700 32900 78756 32902
rect 77308 30716 77364 30772
rect 77308 28866 77364 28868
rect 77308 28814 77310 28866
rect 77310 28814 77362 28866
rect 77362 28814 77364 28866
rect 77308 28812 77364 28814
rect 77308 27916 77364 27972
rect 77308 27074 77364 27076
rect 77308 27022 77310 27074
rect 77310 27022 77362 27074
rect 77362 27022 77364 27074
rect 77308 27020 77364 27022
rect 77644 30994 77700 30996
rect 77644 30942 77646 30994
rect 77646 30942 77698 30994
rect 77698 30942 77700 30994
rect 77644 30940 77700 30942
rect 78204 31724 78260 31780
rect 77532 29820 77588 29876
rect 77868 30156 77924 30212
rect 77756 30098 77812 30100
rect 77756 30046 77758 30098
rect 77758 30046 77810 30098
rect 77810 30046 77812 30098
rect 77756 30044 77812 30046
rect 77644 28700 77700 28756
rect 77868 28812 77924 28868
rect 77980 28700 78036 28756
rect 78092 28476 78148 28532
rect 77756 28140 77812 28196
rect 77868 28364 77924 28420
rect 77980 28252 78036 28308
rect 77532 27244 77588 27300
rect 77308 26572 77364 26628
rect 77308 25730 77364 25732
rect 77308 25678 77310 25730
rect 77310 25678 77362 25730
rect 77362 25678 77364 25730
rect 77308 25676 77364 25678
rect 77420 25618 77476 25620
rect 77420 25566 77422 25618
rect 77422 25566 77474 25618
rect 77474 25566 77476 25618
rect 77420 25564 77476 25566
rect 77644 26962 77700 26964
rect 77644 26910 77646 26962
rect 77646 26910 77698 26962
rect 77698 26910 77700 26962
rect 77644 26908 77700 26910
rect 78092 28140 78148 28196
rect 77980 27468 78036 27524
rect 77868 26572 77924 26628
rect 77756 25900 77812 25956
rect 77644 24834 77700 24836
rect 77644 24782 77646 24834
rect 77646 24782 77698 24834
rect 77698 24782 77700 24834
rect 77644 24780 77700 24782
rect 77532 24668 77588 24724
rect 77308 23884 77364 23940
rect 77420 24556 77476 24612
rect 78092 27186 78148 27188
rect 78092 27134 78094 27186
rect 78094 27134 78146 27186
rect 78146 27134 78148 27186
rect 78092 27132 78148 27134
rect 77532 22258 77588 22260
rect 77532 22206 77534 22258
rect 77534 22206 77586 22258
rect 77586 22206 77588 22258
rect 77532 22204 77588 22206
rect 77308 21644 77364 21700
rect 77532 20914 77588 20916
rect 77532 20862 77534 20914
rect 77534 20862 77586 20914
rect 77586 20862 77588 20914
rect 77532 20860 77588 20862
rect 77308 20524 77364 20580
rect 77532 20130 77588 20132
rect 77532 20078 77534 20130
rect 77534 20078 77586 20130
rect 77586 20078 77588 20130
rect 77532 20076 77588 20078
rect 77196 19180 77252 19236
rect 77756 22146 77812 22148
rect 77756 22094 77758 22146
rect 77758 22094 77810 22146
rect 77810 22094 77812 22146
rect 77756 22092 77812 22094
rect 77868 20802 77924 20804
rect 77868 20750 77870 20802
rect 77870 20750 77922 20802
rect 77922 20750 77924 20802
rect 77868 20748 77924 20750
rect 77532 18562 77588 18564
rect 77532 18510 77534 18562
rect 77534 18510 77586 18562
rect 77586 18510 77588 18562
rect 77532 18508 77588 18510
rect 76076 18284 76132 18340
rect 76076 17666 76132 17668
rect 76076 17614 76078 17666
rect 76078 17614 76130 17666
rect 76130 17614 76132 17666
rect 76076 17612 76132 17614
rect 76076 16882 76132 16884
rect 76076 16830 76078 16882
rect 76078 16830 76130 16882
rect 76130 16830 76132 16882
rect 76076 16828 76132 16830
rect 75964 16492 76020 16548
rect 76076 16604 76132 16660
rect 75964 16098 76020 16100
rect 75964 16046 75966 16098
rect 75966 16046 76018 16098
rect 76018 16046 76020 16098
rect 75964 16044 76020 16046
rect 76748 18450 76804 18452
rect 76748 18398 76750 18450
rect 76750 18398 76802 18450
rect 76802 18398 76804 18450
rect 76748 18396 76804 18398
rect 77756 18396 77812 18452
rect 77420 18284 77476 18340
rect 77308 17724 77364 17780
rect 76748 17612 76804 17668
rect 77420 17276 77476 17332
rect 76636 16604 76692 16660
rect 75404 15538 75460 15540
rect 75404 15486 75406 15538
rect 75406 15486 75458 15538
rect 75458 15486 75460 15538
rect 75404 15484 75460 15486
rect 76188 15484 76244 15540
rect 77420 16604 77476 16660
rect 77756 17276 77812 17332
rect 77084 16044 77140 16100
rect 76748 15932 76804 15988
rect 77308 15986 77364 15988
rect 77308 15934 77310 15986
rect 77310 15934 77362 15986
rect 77362 15934 77364 15986
rect 77308 15932 77364 15934
rect 77420 15484 77476 15540
rect 76748 15314 76804 15316
rect 76748 15262 76750 15314
rect 76750 15262 76802 15314
rect 76802 15262 76804 15314
rect 76748 15260 76804 15262
rect 76860 15426 76916 15428
rect 76860 15374 76862 15426
rect 76862 15374 76914 15426
rect 76914 15374 76916 15426
rect 76860 15372 76916 15374
rect 76188 15036 76244 15092
rect 74956 11394 75012 11396
rect 74956 11342 74958 11394
rect 74958 11342 75010 11394
rect 75010 11342 75012 11394
rect 74956 11340 75012 11342
rect 74732 11170 74788 11172
rect 74732 11118 74734 11170
rect 74734 11118 74786 11170
rect 74786 11118 74788 11170
rect 74732 11116 74788 11118
rect 74732 10780 74788 10836
rect 74844 10610 74900 10612
rect 74844 10558 74846 10610
rect 74846 10558 74898 10610
rect 74898 10558 74900 10610
rect 74844 10556 74900 10558
rect 74956 10498 75012 10500
rect 74956 10446 74958 10498
rect 74958 10446 75010 10498
rect 75010 10446 75012 10498
rect 74956 10444 75012 10446
rect 74956 9938 75012 9940
rect 74956 9886 74958 9938
rect 74958 9886 75010 9938
rect 75010 9886 75012 9938
rect 74956 9884 75012 9886
rect 75404 13522 75460 13524
rect 75404 13470 75406 13522
rect 75406 13470 75458 13522
rect 75458 13470 75460 13522
rect 75404 13468 75460 13470
rect 75292 13356 75348 13412
rect 76076 13804 76132 13860
rect 76412 13580 76468 13636
rect 75516 13132 75572 13188
rect 76300 13356 76356 13412
rect 76076 12962 76132 12964
rect 76076 12910 76078 12962
rect 76078 12910 76130 12962
rect 76130 12910 76132 12962
rect 76076 12908 76132 12910
rect 77532 15426 77588 15428
rect 77532 15374 77534 15426
rect 77534 15374 77586 15426
rect 77586 15374 77588 15426
rect 77532 15372 77588 15374
rect 77420 14754 77476 14756
rect 77420 14702 77422 14754
rect 77422 14702 77474 14754
rect 77474 14702 77476 14754
rect 77420 14700 77476 14702
rect 77980 16604 78036 16660
rect 78092 15538 78148 15540
rect 78092 15486 78094 15538
rect 78094 15486 78146 15538
rect 78146 15486 78148 15538
rect 78092 15484 78148 15486
rect 78492 31386 78548 31388
rect 78492 31334 78494 31386
rect 78494 31334 78546 31386
rect 78546 31334 78548 31386
rect 78492 31332 78548 31334
rect 78596 31386 78652 31388
rect 78596 31334 78598 31386
rect 78598 31334 78650 31386
rect 78650 31334 78652 31386
rect 78596 31332 78652 31334
rect 78700 31386 78756 31388
rect 78700 31334 78702 31386
rect 78702 31334 78754 31386
rect 78754 31334 78756 31386
rect 78700 31332 78756 31334
rect 78492 29818 78548 29820
rect 78492 29766 78494 29818
rect 78494 29766 78546 29818
rect 78546 29766 78548 29818
rect 78492 29764 78548 29766
rect 78596 29818 78652 29820
rect 78596 29766 78598 29818
rect 78598 29766 78650 29818
rect 78650 29766 78652 29818
rect 78596 29764 78652 29766
rect 78700 29818 78756 29820
rect 78700 29766 78702 29818
rect 78702 29766 78754 29818
rect 78754 29766 78756 29818
rect 78700 29764 78756 29766
rect 78316 28476 78372 28532
rect 78492 28250 78548 28252
rect 78492 28198 78494 28250
rect 78494 28198 78546 28250
rect 78546 28198 78548 28250
rect 78492 28196 78548 28198
rect 78596 28250 78652 28252
rect 78596 28198 78598 28250
rect 78598 28198 78650 28250
rect 78650 28198 78652 28250
rect 78596 28196 78652 28198
rect 78700 28250 78756 28252
rect 78700 28198 78702 28250
rect 78702 28198 78754 28250
rect 78754 28198 78756 28250
rect 78700 28196 78756 28198
rect 78492 26682 78548 26684
rect 78492 26630 78494 26682
rect 78494 26630 78546 26682
rect 78546 26630 78548 26682
rect 78492 26628 78548 26630
rect 78596 26682 78652 26684
rect 78596 26630 78598 26682
rect 78598 26630 78650 26682
rect 78650 26630 78652 26682
rect 78596 26628 78652 26630
rect 78700 26682 78756 26684
rect 78700 26630 78702 26682
rect 78702 26630 78754 26682
rect 78754 26630 78756 26682
rect 78700 26628 78756 26630
rect 78316 26460 78372 26516
rect 78492 25114 78548 25116
rect 78492 25062 78494 25114
rect 78494 25062 78546 25114
rect 78546 25062 78548 25114
rect 78492 25060 78548 25062
rect 78596 25114 78652 25116
rect 78596 25062 78598 25114
rect 78598 25062 78650 25114
rect 78650 25062 78652 25114
rect 78596 25060 78652 25062
rect 78700 25114 78756 25116
rect 78700 25062 78702 25114
rect 78702 25062 78754 25114
rect 78754 25062 78756 25114
rect 78700 25060 78756 25062
rect 78492 23546 78548 23548
rect 78492 23494 78494 23546
rect 78494 23494 78546 23546
rect 78546 23494 78548 23546
rect 78492 23492 78548 23494
rect 78596 23546 78652 23548
rect 78596 23494 78598 23546
rect 78598 23494 78650 23546
rect 78650 23494 78652 23546
rect 78596 23492 78652 23494
rect 78700 23546 78756 23548
rect 78700 23494 78702 23546
rect 78702 23494 78754 23546
rect 78754 23494 78756 23546
rect 78700 23492 78756 23494
rect 77756 14700 77812 14756
rect 78316 23212 78372 23268
rect 76972 13634 77028 13636
rect 76972 13582 76974 13634
rect 76974 13582 77026 13634
rect 77026 13582 77028 13634
rect 76972 13580 77028 13582
rect 77420 13468 77476 13524
rect 76188 12178 76244 12180
rect 76188 12126 76190 12178
rect 76190 12126 76242 12178
rect 76242 12126 76244 12178
rect 76188 12124 76244 12126
rect 75516 11452 75572 11508
rect 76188 11900 76244 11956
rect 75628 11394 75684 11396
rect 75628 11342 75630 11394
rect 75630 11342 75682 11394
rect 75682 11342 75684 11394
rect 75628 11340 75684 11342
rect 75852 11116 75908 11172
rect 75740 10722 75796 10724
rect 75740 10670 75742 10722
rect 75742 10670 75794 10722
rect 75794 10670 75796 10722
rect 75740 10668 75796 10670
rect 75628 10444 75684 10500
rect 75180 9212 75236 9268
rect 74956 8988 75012 9044
rect 73388 8204 73444 8260
rect 73612 8258 73668 8260
rect 73612 8206 73614 8258
rect 73614 8206 73666 8258
rect 73666 8206 73668 8258
rect 73612 8204 73668 8206
rect 73276 7756 73332 7812
rect 73164 6690 73220 6692
rect 73164 6638 73166 6690
rect 73166 6638 73218 6690
rect 73218 6638 73220 6690
rect 73164 6636 73220 6638
rect 73612 6300 73668 6356
rect 72604 5794 72660 5796
rect 72604 5742 72606 5794
rect 72606 5742 72658 5794
rect 72658 5742 72660 5794
rect 72604 5740 72660 5742
rect 72380 4844 72436 4900
rect 73052 4732 73108 4788
rect 72604 4562 72660 4564
rect 72604 4510 72606 4562
rect 72606 4510 72658 4562
rect 72658 4510 72660 4562
rect 72604 4508 72660 4510
rect 72380 4284 72436 4340
rect 71932 3276 71988 3332
rect 73500 5628 73556 5684
rect 73388 5180 73444 5236
rect 73276 4562 73332 4564
rect 73276 4510 73278 4562
rect 73278 4510 73330 4562
rect 73330 4510 73332 4562
rect 73276 4508 73332 4510
rect 74284 6748 74340 6804
rect 74060 6466 74116 6468
rect 74060 6414 74062 6466
rect 74062 6414 74114 6466
rect 74114 6414 74116 6466
rect 74060 6412 74116 6414
rect 73836 5516 73892 5572
rect 73948 5122 74004 5124
rect 73948 5070 73950 5122
rect 73950 5070 74002 5122
rect 74002 5070 74004 5122
rect 73948 5068 74004 5070
rect 74284 5292 74340 5348
rect 74620 8258 74676 8260
rect 74620 8206 74622 8258
rect 74622 8206 74674 8258
rect 74674 8206 74676 8258
rect 74620 8204 74676 8206
rect 74732 8034 74788 8036
rect 74732 7982 74734 8034
rect 74734 7982 74786 8034
rect 74786 7982 74788 8034
rect 74732 7980 74788 7982
rect 74620 6412 74676 6468
rect 74508 6130 74564 6132
rect 74508 6078 74510 6130
rect 74510 6078 74562 6130
rect 74562 6078 74564 6130
rect 74508 6076 74564 6078
rect 74172 4956 74228 5012
rect 74396 4898 74452 4900
rect 74396 4846 74398 4898
rect 74398 4846 74450 4898
rect 74450 4846 74452 4898
rect 74396 4844 74452 4846
rect 74732 4956 74788 5012
rect 74620 4508 74676 4564
rect 74172 4060 74228 4116
rect 75852 9324 75908 9380
rect 75964 9212 76020 9268
rect 75628 9100 75684 9156
rect 75516 8930 75572 8932
rect 75516 8878 75518 8930
rect 75518 8878 75570 8930
rect 75570 8878 75572 8930
rect 75516 8876 75572 8878
rect 75404 8370 75460 8372
rect 75404 8318 75406 8370
rect 75406 8318 75458 8370
rect 75458 8318 75460 8370
rect 75404 8316 75460 8318
rect 75516 8258 75572 8260
rect 75516 8206 75518 8258
rect 75518 8206 75570 8258
rect 75570 8206 75572 8258
rect 75516 8204 75572 8206
rect 75292 8092 75348 8148
rect 75964 7980 76020 8036
rect 75068 6412 75124 6468
rect 75292 6636 75348 6692
rect 76076 6748 76132 6804
rect 75068 5794 75124 5796
rect 75068 5742 75070 5794
rect 75070 5742 75122 5794
rect 75122 5742 75124 5794
rect 75068 5740 75124 5742
rect 76524 11506 76580 11508
rect 76524 11454 76526 11506
rect 76526 11454 76578 11506
rect 76578 11454 76580 11506
rect 76524 11452 76580 11454
rect 76412 10668 76468 10724
rect 76300 10498 76356 10500
rect 76300 10446 76302 10498
rect 76302 10446 76354 10498
rect 76354 10446 76356 10498
rect 76300 10444 76356 10446
rect 76524 10556 76580 10612
rect 76748 12290 76804 12292
rect 76748 12238 76750 12290
rect 76750 12238 76802 12290
rect 76802 12238 76804 12290
rect 76748 12236 76804 12238
rect 76972 11228 77028 11284
rect 76748 9324 76804 9380
rect 76860 9154 76916 9156
rect 76860 9102 76862 9154
rect 76862 9102 76914 9154
rect 76914 9102 76916 9154
rect 76860 9100 76916 9102
rect 76748 9042 76804 9044
rect 76748 8990 76750 9042
rect 76750 8990 76802 9042
rect 76802 8990 76804 9042
rect 76748 8988 76804 8990
rect 76636 8316 76692 8372
rect 76860 8204 76916 8260
rect 76300 8092 76356 8148
rect 77308 13186 77364 13188
rect 77308 13134 77310 13186
rect 77310 13134 77362 13186
rect 77362 13134 77364 13186
rect 77308 13132 77364 13134
rect 78492 21978 78548 21980
rect 78492 21926 78494 21978
rect 78494 21926 78546 21978
rect 78546 21926 78548 21978
rect 78492 21924 78548 21926
rect 78596 21978 78652 21980
rect 78596 21926 78598 21978
rect 78598 21926 78650 21978
rect 78650 21926 78652 21978
rect 78596 21924 78652 21926
rect 78700 21978 78756 21980
rect 78700 21926 78702 21978
rect 78702 21926 78754 21978
rect 78754 21926 78756 21978
rect 78700 21924 78756 21926
rect 78492 20410 78548 20412
rect 78492 20358 78494 20410
rect 78494 20358 78546 20410
rect 78546 20358 78548 20410
rect 78492 20356 78548 20358
rect 78596 20410 78652 20412
rect 78596 20358 78598 20410
rect 78598 20358 78650 20410
rect 78650 20358 78652 20410
rect 78596 20356 78652 20358
rect 78700 20410 78756 20412
rect 78700 20358 78702 20410
rect 78702 20358 78754 20410
rect 78754 20358 78756 20410
rect 78700 20356 78756 20358
rect 78492 18842 78548 18844
rect 78492 18790 78494 18842
rect 78494 18790 78546 18842
rect 78546 18790 78548 18842
rect 78492 18788 78548 18790
rect 78596 18842 78652 18844
rect 78596 18790 78598 18842
rect 78598 18790 78650 18842
rect 78650 18790 78652 18842
rect 78596 18788 78652 18790
rect 78700 18842 78756 18844
rect 78700 18790 78702 18842
rect 78702 18790 78754 18842
rect 78754 18790 78756 18842
rect 78700 18788 78756 18790
rect 79100 28028 79156 28084
rect 78988 26908 79044 26964
rect 78988 20076 79044 20132
rect 78876 17388 78932 17444
rect 78492 17274 78548 17276
rect 78492 17222 78494 17274
rect 78494 17222 78546 17274
rect 78546 17222 78548 17274
rect 78492 17220 78548 17222
rect 78596 17274 78652 17276
rect 78596 17222 78598 17274
rect 78598 17222 78650 17274
rect 78650 17222 78652 17274
rect 78596 17220 78652 17222
rect 78700 17274 78756 17276
rect 78700 17222 78702 17274
rect 78702 17222 78754 17274
rect 78754 17222 78756 17274
rect 78700 17220 78756 17222
rect 78492 15706 78548 15708
rect 78492 15654 78494 15706
rect 78494 15654 78546 15706
rect 78546 15654 78548 15706
rect 78492 15652 78548 15654
rect 78596 15706 78652 15708
rect 78596 15654 78598 15706
rect 78598 15654 78650 15706
rect 78650 15654 78652 15706
rect 78596 15652 78652 15654
rect 78700 15706 78756 15708
rect 78700 15654 78702 15706
rect 78702 15654 78754 15706
rect 78754 15654 78756 15706
rect 78700 15652 78756 15654
rect 77420 12908 77476 12964
rect 77868 12124 77924 12180
rect 77532 11452 77588 11508
rect 77196 11228 77252 11284
rect 77644 11282 77700 11284
rect 77644 11230 77646 11282
rect 77646 11230 77698 11282
rect 77698 11230 77700 11282
rect 77644 11228 77700 11230
rect 77532 10668 77588 10724
rect 77532 9324 77588 9380
rect 77420 9266 77476 9268
rect 77420 9214 77422 9266
rect 77422 9214 77474 9266
rect 77474 9214 77476 9266
rect 77420 9212 77476 9214
rect 77308 8316 77364 8372
rect 77532 8258 77588 8260
rect 77532 8206 77534 8258
rect 77534 8206 77586 8258
rect 77586 8206 77588 8258
rect 77532 8204 77588 8206
rect 77308 8092 77364 8148
rect 77532 6748 77588 6804
rect 77420 6690 77476 6692
rect 77420 6638 77422 6690
rect 77422 6638 77474 6690
rect 77474 6638 77476 6690
rect 77420 6636 77476 6638
rect 77308 6578 77364 6580
rect 77308 6526 77310 6578
rect 77310 6526 77362 6578
rect 77362 6526 77364 6578
rect 77308 6524 77364 6526
rect 76972 5906 77028 5908
rect 76972 5854 76974 5906
rect 76974 5854 77026 5906
rect 77026 5854 77028 5906
rect 76972 5852 77028 5854
rect 75516 5292 75572 5348
rect 76300 5346 76356 5348
rect 76300 5294 76302 5346
rect 76302 5294 76354 5346
rect 76354 5294 76356 5346
rect 76300 5292 76356 5294
rect 75516 5122 75572 5124
rect 75516 5070 75518 5122
rect 75518 5070 75570 5122
rect 75570 5070 75572 5122
rect 75516 5068 75572 5070
rect 75628 4956 75684 5012
rect 77532 5852 77588 5908
rect 77980 10722 78036 10724
rect 77980 10670 77982 10722
rect 77982 10670 78034 10722
rect 78034 10670 78036 10722
rect 77980 10668 78036 10670
rect 78092 10610 78148 10612
rect 78092 10558 78094 10610
rect 78094 10558 78146 10610
rect 78146 10558 78148 10610
rect 78092 10556 78148 10558
rect 77980 10386 78036 10388
rect 77980 10334 77982 10386
rect 77982 10334 78034 10386
rect 78034 10334 78036 10386
rect 77980 10332 78036 10334
rect 77868 8540 77924 8596
rect 78492 14138 78548 14140
rect 78492 14086 78494 14138
rect 78494 14086 78546 14138
rect 78546 14086 78548 14138
rect 78492 14084 78548 14086
rect 78596 14138 78652 14140
rect 78596 14086 78598 14138
rect 78598 14086 78650 14138
rect 78650 14086 78652 14138
rect 78596 14084 78652 14086
rect 78700 14138 78756 14140
rect 78700 14086 78702 14138
rect 78702 14086 78754 14138
rect 78754 14086 78756 14138
rect 78700 14084 78756 14086
rect 78492 12570 78548 12572
rect 78492 12518 78494 12570
rect 78494 12518 78546 12570
rect 78546 12518 78548 12570
rect 78492 12516 78548 12518
rect 78596 12570 78652 12572
rect 78596 12518 78598 12570
rect 78598 12518 78650 12570
rect 78650 12518 78652 12570
rect 78596 12516 78652 12518
rect 78700 12570 78756 12572
rect 78700 12518 78702 12570
rect 78702 12518 78754 12570
rect 78754 12518 78756 12570
rect 78700 12516 78756 12518
rect 78492 11002 78548 11004
rect 78492 10950 78494 11002
rect 78494 10950 78546 11002
rect 78546 10950 78548 11002
rect 78492 10948 78548 10950
rect 78596 11002 78652 11004
rect 78596 10950 78598 11002
rect 78598 10950 78650 11002
rect 78650 10950 78652 11002
rect 78596 10948 78652 10950
rect 78700 11002 78756 11004
rect 78700 10950 78702 11002
rect 78702 10950 78754 11002
rect 78754 10950 78756 11002
rect 78700 10948 78756 10950
rect 78316 9884 78372 9940
rect 77756 6076 77812 6132
rect 76972 5292 77028 5348
rect 77196 5234 77252 5236
rect 77196 5182 77198 5234
rect 77198 5182 77250 5234
rect 77250 5182 77252 5234
rect 77196 5180 77252 5182
rect 78092 5122 78148 5124
rect 78092 5070 78094 5122
rect 78094 5070 78146 5122
rect 78146 5070 78148 5122
rect 78092 5068 78148 5070
rect 77644 4956 77700 5012
rect 75516 3948 75572 4004
rect 74844 3836 74900 3892
rect 76748 3836 76804 3892
rect 75516 3554 75572 3556
rect 75516 3502 75518 3554
rect 75518 3502 75570 3554
rect 75570 3502 75572 3554
rect 75516 3500 75572 3502
rect 77196 3836 77252 3892
rect 74844 1484 74900 1540
rect 77308 3666 77364 3668
rect 77308 3614 77310 3666
rect 77310 3614 77362 3666
rect 77362 3614 77364 3666
rect 77308 3612 77364 3614
rect 78492 9434 78548 9436
rect 78492 9382 78494 9434
rect 78494 9382 78546 9434
rect 78546 9382 78548 9434
rect 78492 9380 78548 9382
rect 78596 9434 78652 9436
rect 78596 9382 78598 9434
rect 78598 9382 78650 9434
rect 78650 9382 78652 9434
rect 78596 9380 78652 9382
rect 78700 9434 78756 9436
rect 78700 9382 78702 9434
rect 78702 9382 78754 9434
rect 78754 9382 78756 9434
rect 78700 9380 78756 9382
rect 78492 7866 78548 7868
rect 78492 7814 78494 7866
rect 78494 7814 78546 7866
rect 78546 7814 78548 7866
rect 78492 7812 78548 7814
rect 78596 7866 78652 7868
rect 78596 7814 78598 7866
rect 78598 7814 78650 7866
rect 78650 7814 78652 7866
rect 78596 7812 78652 7814
rect 78700 7866 78756 7868
rect 78700 7814 78702 7866
rect 78702 7814 78754 7866
rect 78754 7814 78756 7866
rect 78700 7812 78756 7814
rect 78492 6298 78548 6300
rect 78492 6246 78494 6298
rect 78494 6246 78546 6298
rect 78546 6246 78548 6298
rect 78492 6244 78548 6246
rect 78596 6298 78652 6300
rect 78596 6246 78598 6298
rect 78598 6246 78650 6298
rect 78650 6246 78652 6298
rect 78596 6244 78652 6246
rect 78700 6298 78756 6300
rect 78700 6246 78702 6298
rect 78702 6246 78754 6298
rect 78754 6246 78756 6298
rect 78700 6244 78756 6246
rect 78492 4730 78548 4732
rect 78492 4678 78494 4730
rect 78494 4678 78546 4730
rect 78546 4678 78548 4730
rect 78492 4676 78548 4678
rect 78596 4730 78652 4732
rect 78596 4678 78598 4730
rect 78598 4678 78650 4730
rect 78650 4678 78652 4730
rect 78596 4676 78652 4678
rect 78700 4730 78756 4732
rect 78700 4678 78702 4730
rect 78702 4678 78754 4730
rect 78754 4678 78756 4730
rect 78700 4676 78756 4678
rect 77644 3500 77700 3556
rect 77756 3442 77812 3444
rect 77756 3390 77758 3442
rect 77758 3390 77810 3442
rect 77810 3390 77812 3442
rect 77756 3388 77812 3390
rect 78492 3162 78548 3164
rect 78492 3110 78494 3162
rect 78494 3110 78546 3162
rect 78546 3110 78548 3162
rect 78492 3108 78548 3110
rect 78596 3162 78652 3164
rect 78596 3110 78598 3162
rect 78598 3110 78650 3162
rect 78650 3110 78652 3162
rect 78596 3108 78652 3110
rect 78700 3162 78756 3164
rect 78700 3110 78702 3162
rect 78702 3110 78754 3162
rect 78754 3110 78756 3162
rect 78700 3108 78756 3110
<< metal3 >>
rect 0 38500 800 38528
rect 79200 38500 80000 38528
rect 0 38444 2156 38500
rect 2212 38444 2222 38500
rect 77858 38444 77868 38500
rect 77924 38444 80000 38500
rect 0 38416 800 38444
rect 79200 38416 80000 38444
rect 40226 37996 40236 38052
rect 40292 37996 75404 38052
rect 75460 37996 75470 38052
rect 33954 37884 33964 37940
rect 34020 37884 68460 37940
rect 68516 37884 68526 37940
rect 24882 37772 24892 37828
rect 24948 37772 71148 37828
rect 71204 37772 71214 37828
rect 2482 37660 2492 37716
rect 2548 37660 53676 37716
rect 53732 37660 53742 37716
rect 9986 37548 9996 37604
rect 10052 37548 63196 37604
rect 63252 37548 63262 37604
rect 2258 37436 2268 37492
rect 2324 37436 57708 37492
rect 57764 37436 57774 37492
rect 18834 37324 18844 37380
rect 18900 37324 77084 37380
rect 77140 37324 77150 37380
rect 15474 37212 15484 37268
rect 15540 37212 73500 37268
rect 73556 37212 73566 37268
rect 5058 37100 5068 37156
rect 5124 37100 67452 37156
rect 67508 37100 67518 37156
rect 7074 36988 7084 37044
rect 7140 36988 70476 37044
rect 70532 36988 70542 37044
rect 10862 36820 10872 36876
rect 10928 36820 10976 36876
rect 11032 36820 11080 36876
rect 11136 36820 11146 36876
rect 30182 36820 30192 36876
rect 30248 36820 30296 36876
rect 30352 36820 30400 36876
rect 30456 36820 30466 36876
rect 49502 36820 49512 36876
rect 49568 36820 49616 36876
rect 49672 36820 49720 36876
rect 49776 36820 49786 36876
rect 68822 36820 68832 36876
rect 68888 36820 68936 36876
rect 68992 36820 69040 36876
rect 69096 36820 69106 36876
rect 52210 36764 52220 36820
rect 52276 36764 55468 36820
rect 55412 36708 55468 36764
rect 31892 36652 33964 36708
rect 34020 36652 34030 36708
rect 55412 36652 71708 36708
rect 71764 36652 71774 36708
rect 31892 36596 31948 36652
rect 21858 36540 21868 36596
rect 21924 36540 22764 36596
rect 22820 36540 24892 36596
rect 24948 36540 24958 36596
rect 27794 36540 27804 36596
rect 27860 36540 31948 36596
rect 33506 36540 33516 36596
rect 33572 36540 35196 36596
rect 35252 36540 43876 36596
rect 48514 36540 48524 36596
rect 48580 36540 48972 36596
rect 49028 36540 49038 36596
rect 53442 36540 53452 36596
rect 53508 36540 54348 36596
rect 54404 36540 54414 36596
rect 58370 36540 58380 36596
rect 58436 36540 58828 36596
rect 58884 36540 58894 36596
rect 63298 36540 63308 36596
rect 63364 36540 64652 36596
rect 64708 36540 64718 36596
rect 73154 36540 73164 36596
rect 73220 36540 74060 36596
rect 74116 36540 74126 36596
rect 75394 36540 75404 36596
rect 75460 36540 77980 36596
rect 78036 36540 78046 36596
rect 43820 36484 43876 36540
rect 3154 36428 3164 36484
rect 3220 36428 6076 36484
rect 6132 36428 6142 36484
rect 13682 36428 13692 36484
rect 13748 36428 15484 36484
rect 15540 36428 15550 36484
rect 24546 36428 24556 36484
rect 24612 36428 25228 36484
rect 25284 36428 25294 36484
rect 34962 36428 34972 36484
rect 35028 36428 35644 36484
rect 35700 36428 35710 36484
rect 35858 36428 35868 36484
rect 35924 36428 38668 36484
rect 38724 36428 38734 36484
rect 43810 36428 43820 36484
rect 43876 36428 74172 36484
rect 74228 36428 74238 36484
rect 5282 36316 5292 36372
rect 5348 36316 9996 36372
rect 10052 36316 10062 36372
rect 15586 36316 15596 36372
rect 15652 36316 17948 36372
rect 18004 36316 18508 36372
rect 18564 36316 18574 36372
rect 23874 36316 23884 36372
rect 23940 36316 25788 36372
rect 25844 36316 27356 36372
rect 27412 36316 27422 36372
rect 28578 36316 28588 36372
rect 28644 36316 30492 36372
rect 30548 36316 31948 36372
rect 34850 36316 34860 36372
rect 34916 36316 36092 36372
rect 36148 36316 36158 36372
rect 60050 36316 60060 36372
rect 60116 36316 62860 36372
rect 62916 36316 62926 36372
rect 63186 36316 63196 36372
rect 63252 36316 68684 36372
rect 68740 36316 68750 36372
rect 70466 36316 70476 36372
rect 70532 36316 73164 36372
rect 73220 36316 73388 36372
rect 73444 36316 73454 36372
rect 31892 36260 31948 36316
rect 14354 36204 14364 36260
rect 14420 36204 16380 36260
rect 16436 36204 18844 36260
rect 18900 36204 18910 36260
rect 26114 36204 26124 36260
rect 26180 36204 29596 36260
rect 29652 36204 29662 36260
rect 31892 36204 36988 36260
rect 37044 36204 37054 36260
rect 42578 36204 42588 36260
rect 42644 36204 43036 36260
rect 43092 36204 44380 36260
rect 44436 36204 44446 36260
rect 45266 36204 45276 36260
rect 45332 36204 47180 36260
rect 47236 36204 47246 36260
rect 59826 36204 59836 36260
rect 59892 36204 60508 36260
rect 60564 36204 60574 36260
rect 65874 36204 65884 36260
rect 65940 36204 67900 36260
rect 67956 36204 67966 36260
rect 72818 36204 72828 36260
rect 72884 36204 74956 36260
rect 75012 36204 75022 36260
rect 8082 36092 8092 36148
rect 8148 36092 8540 36148
rect 8596 36092 16604 36148
rect 16660 36092 16670 36148
rect 42690 36092 42700 36148
rect 42756 36092 45500 36148
rect 45556 36092 47908 36148
rect 71138 36092 71148 36148
rect 71204 36092 73276 36148
rect 73332 36092 73342 36148
rect 0 36036 800 36064
rect 20522 36036 20532 36092
rect 20588 36036 20636 36092
rect 20692 36036 20740 36092
rect 20796 36036 20806 36092
rect 39842 36036 39852 36092
rect 39908 36036 39956 36092
rect 40012 36036 40060 36092
rect 40116 36036 40126 36092
rect 47852 36036 47908 36092
rect 59162 36036 59172 36092
rect 59228 36036 59276 36092
rect 59332 36036 59380 36092
rect 59436 36036 59446 36092
rect 78482 36036 78492 36092
rect 78548 36036 78596 36092
rect 78652 36036 78700 36092
rect 78756 36036 78766 36092
rect 79200 36036 80000 36064
rect 0 35980 1932 36036
rect 1988 35980 1998 36036
rect 47842 35980 47852 36036
rect 47908 35980 48300 36036
rect 48356 35980 49756 36036
rect 49812 35980 49822 36036
rect 67442 35980 67452 36036
rect 67508 35980 75740 36036
rect 75796 35980 76300 36036
rect 76356 35980 76366 36036
rect 78876 35980 80000 36036
rect 0 35952 800 35980
rect 78876 35924 78932 35980
rect 79200 35952 80000 35980
rect 4946 35868 4956 35924
rect 5012 35868 5628 35924
rect 5684 35868 23212 35924
rect 23268 35868 23278 35924
rect 26786 35868 26796 35924
rect 26852 35868 27468 35924
rect 27524 35868 27534 35924
rect 28466 35868 28476 35924
rect 28532 35868 31948 35924
rect 32050 35868 32060 35924
rect 32116 35868 32732 35924
rect 32788 35868 34972 35924
rect 35028 35868 35038 35924
rect 40114 35868 40124 35924
rect 40180 35868 40572 35924
rect 40628 35868 52220 35924
rect 52276 35868 52286 35924
rect 53106 35868 53116 35924
rect 53172 35868 72492 35924
rect 72548 35868 72558 35924
rect 76066 35868 76076 35924
rect 76132 35868 78932 35924
rect 31892 35812 31948 35868
rect 3042 35756 3052 35812
rect 3108 35756 3612 35812
rect 3668 35756 3678 35812
rect 4834 35756 4844 35812
rect 4900 35756 5292 35812
rect 5348 35756 5358 35812
rect 11890 35756 11900 35812
rect 11956 35756 15036 35812
rect 15092 35756 15596 35812
rect 15652 35756 15662 35812
rect 16482 35756 16492 35812
rect 16548 35756 17836 35812
rect 17892 35756 17902 35812
rect 26002 35756 26012 35812
rect 26068 35756 26460 35812
rect 26516 35756 28588 35812
rect 28644 35756 28654 35812
rect 31892 35756 32396 35812
rect 32452 35756 34860 35812
rect 34916 35756 34926 35812
rect 52098 35756 52108 35812
rect 52164 35756 52780 35812
rect 52836 35756 52846 35812
rect 71698 35756 71708 35812
rect 71764 35756 72268 35812
rect 72324 35756 72334 35812
rect 72594 35756 72604 35812
rect 72660 35756 76748 35812
rect 76804 35756 76814 35812
rect 10994 35644 11004 35700
rect 11060 35644 12012 35700
rect 12068 35644 12078 35700
rect 12226 35644 12236 35700
rect 12292 35644 12908 35700
rect 12964 35644 12974 35700
rect 16370 35644 16380 35700
rect 16436 35644 17276 35700
rect 17332 35644 17342 35700
rect 18050 35644 18060 35700
rect 18116 35644 19628 35700
rect 19684 35644 19964 35700
rect 20020 35644 20030 35700
rect 22418 35644 22428 35700
rect 22484 35644 23324 35700
rect 23380 35644 23660 35700
rect 23716 35644 23726 35700
rect 27458 35644 27468 35700
rect 27524 35644 28476 35700
rect 28532 35644 29820 35700
rect 29876 35644 29886 35700
rect 32834 35644 32844 35700
rect 32900 35644 33628 35700
rect 33684 35644 33694 35700
rect 44146 35644 44156 35700
rect 44212 35644 45612 35700
rect 45668 35644 45678 35700
rect 47170 35644 47180 35700
rect 47236 35644 48076 35700
rect 48132 35644 48524 35700
rect 48580 35644 48590 35700
rect 50652 35644 53116 35700
rect 53172 35644 53182 35700
rect 55346 35644 55356 35700
rect 55412 35644 55916 35700
rect 55972 35644 55982 35700
rect 58034 35644 58044 35700
rect 58100 35644 60732 35700
rect 60788 35644 61404 35700
rect 61460 35644 61470 35700
rect 64754 35644 64764 35700
rect 64820 35644 65548 35700
rect 65604 35644 66220 35700
rect 66276 35644 66286 35700
rect 50652 35588 50708 35644
rect 3938 35532 3948 35588
rect 4004 35532 4844 35588
rect 4900 35532 4910 35588
rect 15138 35532 15148 35588
rect 15204 35532 16044 35588
rect 16100 35532 16110 35588
rect 22978 35532 22988 35588
rect 23044 35532 25900 35588
rect 25956 35532 26236 35588
rect 26292 35532 26302 35588
rect 37650 35532 37660 35588
rect 37716 35532 38108 35588
rect 38164 35532 50708 35588
rect 51874 35532 51884 35588
rect 51940 35532 52556 35588
rect 52612 35532 52622 35588
rect 56578 35532 56588 35588
rect 56644 35532 57484 35588
rect 57540 35532 58940 35588
rect 58996 35532 59006 35588
rect 61842 35532 61852 35588
rect 61908 35532 62860 35588
rect 62916 35532 62926 35588
rect 64530 35532 64540 35588
rect 64596 35532 65772 35588
rect 65828 35532 65838 35588
rect 67554 35532 67564 35588
rect 67620 35532 68348 35588
rect 68404 35532 69468 35588
rect 69524 35532 69534 35588
rect 35522 35420 35532 35476
rect 35588 35420 46172 35476
rect 46228 35420 46238 35476
rect 57026 35420 57036 35476
rect 57092 35420 57708 35476
rect 57764 35420 57774 35476
rect 58258 35420 58268 35476
rect 58324 35420 59612 35476
rect 59668 35420 59678 35476
rect 66658 35420 66668 35476
rect 66724 35420 69580 35476
rect 69636 35420 69646 35476
rect 3042 35308 3052 35364
rect 3108 35308 4508 35364
rect 4564 35308 4574 35364
rect 60610 35308 60620 35364
rect 60676 35308 62524 35364
rect 62580 35308 62972 35364
rect 63028 35308 63038 35364
rect 10862 35252 10872 35308
rect 10928 35252 10976 35308
rect 11032 35252 11080 35308
rect 11136 35252 11146 35308
rect 30182 35252 30192 35308
rect 30248 35252 30296 35308
rect 30352 35252 30400 35308
rect 30456 35252 30466 35308
rect 49502 35252 49512 35308
rect 49568 35252 49616 35308
rect 49672 35252 49720 35308
rect 49776 35252 49786 35308
rect 68822 35252 68832 35308
rect 68888 35252 68936 35308
rect 68992 35252 69040 35308
rect 69096 35252 69106 35308
rect 12114 35196 12124 35252
rect 12180 35196 13916 35252
rect 13972 35196 13982 35252
rect 15026 35196 15036 35252
rect 15092 35196 21532 35252
rect 21588 35196 22652 35252
rect 22708 35196 22718 35252
rect 36978 35196 36988 35252
rect 37044 35196 40236 35252
rect 40292 35196 40302 35252
rect 44706 35196 44716 35252
rect 44772 35196 46508 35252
rect 46564 35196 48188 35252
rect 48244 35196 49308 35252
rect 49364 35196 49374 35252
rect 56018 35196 56028 35252
rect 56084 35196 57260 35252
rect 57316 35196 59164 35252
rect 59220 35196 60284 35252
rect 60340 35196 60350 35252
rect 62290 35196 62300 35252
rect 62356 35196 64988 35252
rect 65044 35196 65660 35252
rect 65716 35196 65726 35252
rect 69356 35196 77532 35252
rect 77588 35196 77598 35252
rect 69356 35140 69412 35196
rect 12002 35084 12012 35140
rect 12068 35084 18732 35140
rect 18788 35084 19740 35140
rect 19796 35084 19806 35140
rect 20066 35084 20076 35140
rect 20132 35084 23100 35140
rect 23156 35084 23548 35140
rect 23604 35084 23614 35140
rect 30258 35084 30268 35140
rect 30324 35084 31052 35140
rect 31108 35084 31118 35140
rect 31266 35084 31276 35140
rect 31332 35084 69412 35140
rect 69468 35084 77980 35140
rect 78036 35084 78046 35140
rect 69468 35028 69524 35084
rect 3938 34972 3948 35028
rect 4004 34972 4396 35028
rect 4452 34972 7084 35028
rect 7140 34972 7150 35028
rect 13234 34972 13244 35028
rect 13300 34972 13580 35028
rect 13636 34972 14140 35028
rect 14196 34972 14924 35028
rect 14980 34972 17724 35028
rect 17780 34972 17790 35028
rect 18620 34972 20412 35028
rect 20468 34972 69524 35028
rect 69682 34972 69692 35028
rect 69748 34972 72268 35028
rect 72324 34972 72334 35028
rect 76066 34972 76076 35028
rect 76132 34972 78092 35028
rect 78148 34972 78158 35028
rect 8978 34860 8988 34916
rect 9044 34860 11340 34916
rect 11396 34860 11406 34916
rect 13010 34860 13020 34916
rect 13076 34860 14364 34916
rect 14420 34860 16380 34916
rect 16436 34860 16446 34916
rect 18620 34804 18676 34972
rect 19730 34860 19740 34916
rect 19796 34860 20524 34916
rect 20580 34860 20590 34916
rect 25330 34860 25340 34916
rect 25396 34860 26796 34916
rect 26852 34860 27132 34916
rect 27188 34860 27198 34916
rect 28354 34860 28364 34916
rect 28420 34860 34748 34916
rect 34804 34860 35420 34916
rect 35476 34860 35486 34916
rect 35634 34860 35644 34916
rect 35700 34860 36540 34916
rect 36596 34860 37436 34916
rect 37492 34860 37502 34916
rect 40450 34860 40460 34916
rect 40516 34860 41356 34916
rect 41412 34860 42028 34916
rect 42084 34860 42094 34916
rect 44930 34860 44940 34916
rect 44996 34860 45388 34916
rect 45444 34860 45454 34916
rect 46162 34860 46172 34916
rect 46228 34860 47180 34916
rect 47236 34860 47246 34916
rect 48738 34860 48748 34916
rect 48804 34860 50876 34916
rect 50932 34860 50942 34916
rect 57698 34860 57708 34916
rect 57764 34860 59052 34916
rect 59108 34860 59118 34916
rect 64194 34860 64204 34916
rect 64260 34860 64988 34916
rect 65044 34860 65054 34916
rect 65314 34860 65324 34916
rect 65380 34860 67116 34916
rect 67172 34860 67182 34916
rect 68674 34860 68684 34916
rect 68740 34860 73948 34916
rect 74004 34860 74956 34916
rect 75012 34860 75022 34916
rect 35644 34804 35700 34860
rect 65324 34804 65380 34860
rect 12898 34748 12908 34804
rect 12964 34748 13692 34804
rect 13748 34748 13758 34804
rect 15810 34748 15820 34804
rect 15876 34748 18620 34804
rect 18676 34748 18686 34804
rect 25442 34748 25452 34804
rect 25508 34748 28476 34804
rect 28532 34748 31276 34804
rect 31332 34748 31342 34804
rect 35074 34748 35084 34804
rect 35140 34748 35700 34804
rect 36642 34748 36652 34804
rect 36708 34748 37548 34804
rect 37604 34748 37614 34804
rect 38612 34748 46620 34804
rect 46676 34748 47516 34804
rect 47572 34748 47740 34804
rect 47796 34748 47806 34804
rect 48626 34748 48636 34804
rect 48692 34748 49756 34804
rect 49812 34748 49822 34804
rect 55906 34748 55916 34804
rect 55972 34748 56812 34804
rect 56868 34748 57596 34804
rect 57652 34748 57662 34804
rect 63186 34748 63196 34804
rect 63252 34748 63980 34804
rect 64036 34748 64046 34804
rect 64418 34748 64428 34804
rect 64484 34748 65380 34804
rect 67172 34748 69468 34804
rect 69524 34748 69534 34804
rect 71362 34748 71372 34804
rect 71428 34748 72492 34804
rect 72548 34748 72558 34804
rect 77074 34748 77084 34804
rect 77140 34748 78092 34804
rect 78148 34748 78158 34804
rect 38612 34692 38668 34748
rect 67172 34692 67228 34748
rect 3042 34636 3052 34692
rect 3108 34636 3612 34692
rect 3668 34636 3678 34692
rect 9762 34636 9772 34692
rect 9828 34636 18172 34692
rect 18228 34636 18238 34692
rect 24994 34636 25004 34692
rect 25060 34636 25676 34692
rect 25732 34636 26012 34692
rect 26068 34636 26078 34692
rect 30370 34636 30380 34692
rect 30436 34636 36204 34692
rect 36260 34636 36270 34692
rect 37650 34636 37660 34692
rect 37716 34636 38668 34692
rect 43474 34636 43484 34692
rect 43540 34636 49980 34692
rect 50036 34636 50046 34692
rect 50306 34636 50316 34692
rect 50372 34636 51996 34692
rect 52052 34636 52062 34692
rect 59378 34636 59388 34692
rect 59444 34636 59668 34692
rect 64082 34636 64092 34692
rect 64148 34636 65660 34692
rect 65716 34636 65996 34692
rect 66052 34636 67228 34692
rect 59612 34580 59668 34636
rect 10434 34524 10444 34580
rect 10500 34524 15260 34580
rect 15316 34524 15326 34580
rect 59612 34524 64764 34580
rect 64820 34524 64830 34580
rect 66434 34524 66444 34580
rect 66500 34524 69692 34580
rect 69748 34524 69758 34580
rect 20522 34468 20532 34524
rect 20588 34468 20636 34524
rect 20692 34468 20740 34524
rect 20796 34468 20806 34524
rect 39842 34468 39852 34524
rect 39908 34468 39956 34524
rect 40012 34468 40060 34524
rect 40116 34468 40126 34524
rect 59162 34468 59172 34524
rect 59228 34468 59276 34524
rect 59332 34468 59380 34524
rect 59436 34468 59446 34524
rect 78482 34468 78492 34524
rect 78548 34468 78596 34524
rect 78652 34468 78700 34524
rect 78756 34468 78766 34524
rect 24770 34412 24780 34468
rect 24836 34412 29596 34468
rect 29652 34412 30716 34468
rect 30772 34412 31500 34468
rect 31556 34412 31566 34468
rect 51202 34412 51212 34468
rect 51268 34412 51278 34468
rect 60722 34412 60732 34468
rect 60788 34412 61292 34468
rect 61348 34412 61358 34468
rect 51212 34356 51268 34412
rect 16818 34300 16828 34356
rect 16884 34300 17836 34356
rect 17892 34300 17902 34356
rect 27458 34300 27468 34356
rect 27524 34300 30268 34356
rect 30324 34300 30334 34356
rect 33842 34300 33852 34356
rect 33908 34300 39676 34356
rect 39732 34300 40460 34356
rect 40516 34300 40526 34356
rect 40674 34300 40684 34356
rect 40740 34300 42812 34356
rect 42868 34300 43596 34356
rect 43652 34300 43662 34356
rect 51212 34300 64092 34356
rect 64148 34300 64158 34356
rect 64978 34300 64988 34356
rect 65044 34300 65772 34356
rect 65828 34300 65838 34356
rect 11666 34188 11676 34244
rect 11732 34188 13468 34244
rect 13524 34188 13534 34244
rect 14690 34188 14700 34244
rect 14756 34188 16940 34244
rect 16996 34188 21196 34244
rect 21252 34188 24892 34244
rect 24948 34188 24958 34244
rect 26450 34188 26460 34244
rect 26516 34188 27244 34244
rect 27300 34188 27310 34244
rect 32610 34188 32620 34244
rect 32676 34188 34244 34244
rect 35746 34188 35756 34244
rect 35812 34188 41468 34244
rect 41524 34188 41534 34244
rect 41682 34188 41692 34244
rect 41748 34188 43932 34244
rect 43988 34188 45052 34244
rect 45108 34188 45118 34244
rect 34188 34132 34244 34188
rect 51212 34132 51268 34300
rect 55122 34188 55132 34244
rect 55188 34188 57932 34244
rect 57988 34188 59388 34244
rect 59444 34188 61516 34244
rect 61572 34188 61582 34244
rect 63858 34188 63868 34244
rect 63924 34188 71148 34244
rect 71204 34188 71484 34244
rect 71540 34188 71550 34244
rect 73602 34188 73612 34244
rect 73668 34188 74060 34244
rect 74116 34188 74126 34244
rect 76738 34188 76748 34244
rect 76804 34188 78876 34244
rect 78932 34188 78942 34244
rect 23874 34076 23884 34132
rect 23940 34076 25900 34132
rect 25956 34076 26236 34132
rect 26292 34076 26302 34132
rect 31892 34076 32060 34132
rect 32116 34076 32844 34132
rect 32900 34076 33964 34132
rect 34020 34076 34030 34132
rect 34188 34076 51268 34132
rect 51874 34076 51884 34132
rect 51940 34076 52780 34132
rect 52836 34076 52846 34132
rect 60498 34076 60508 34132
rect 60564 34076 63084 34132
rect 63140 34076 65100 34132
rect 65156 34076 65166 34132
rect 65986 34076 65996 34132
rect 66052 34076 66444 34132
rect 66500 34076 66668 34132
rect 66724 34076 66734 34132
rect 77522 34076 77532 34132
rect 77588 34076 77980 34132
rect 78036 34076 78204 34132
rect 78260 34076 78270 34132
rect 31892 34020 31948 34076
rect 28690 33964 28700 34020
rect 28756 33964 31948 34020
rect 55682 33964 55692 34020
rect 55748 33964 57484 34020
rect 57540 33964 57550 34020
rect 8754 33852 8764 33908
rect 8820 33852 14364 33908
rect 14420 33852 14812 33908
rect 14868 33852 14878 33908
rect 18162 33852 18172 33908
rect 18228 33852 20188 33908
rect 20244 33852 21980 33908
rect 22036 33852 22988 33908
rect 23044 33852 23436 33908
rect 23492 33852 23502 33908
rect 23874 33852 23884 33908
rect 23940 33852 26460 33908
rect 26516 33852 26526 33908
rect 31602 33852 31612 33908
rect 31668 33852 36764 33908
rect 36820 33852 37212 33908
rect 37268 33852 37278 33908
rect 38658 33852 38668 33908
rect 38724 33852 42252 33908
rect 42308 33852 44044 33908
rect 44100 33852 44110 33908
rect 54898 33852 54908 33908
rect 54964 33852 57820 33908
rect 57876 33852 57886 33908
rect 67106 33852 67116 33908
rect 67172 33852 70140 33908
rect 70196 33852 71820 33908
rect 71876 33852 72156 33908
rect 72212 33852 72222 33908
rect 42812 33796 42868 33852
rect 17938 33740 17948 33796
rect 18004 33740 18014 33796
rect 42802 33740 42812 33796
rect 42868 33740 42878 33796
rect 57586 33740 57596 33796
rect 57652 33740 62524 33796
rect 62580 33740 62590 33796
rect 10862 33684 10872 33740
rect 10928 33684 10976 33740
rect 11032 33684 11080 33740
rect 11136 33684 11146 33740
rect 17948 33684 18004 33740
rect 30182 33684 30192 33740
rect 30248 33684 30296 33740
rect 30352 33684 30400 33740
rect 30456 33684 30466 33740
rect 49502 33684 49512 33740
rect 49568 33684 49616 33740
rect 49672 33684 49720 33740
rect 49776 33684 49786 33740
rect 68822 33684 68832 33740
rect 68888 33684 68936 33740
rect 68992 33684 69040 33740
rect 69096 33684 69106 33740
rect 13682 33628 13692 33684
rect 13748 33628 14364 33684
rect 14420 33628 15148 33684
rect 15204 33628 17276 33684
rect 17332 33628 17612 33684
rect 17668 33628 18004 33684
rect 20178 33628 20188 33684
rect 20244 33628 22764 33684
rect 22820 33628 23324 33684
rect 23380 33628 24332 33684
rect 24388 33628 24398 33684
rect 47170 33628 47180 33684
rect 47236 33628 48412 33684
rect 48468 33628 48478 33684
rect 76066 33628 76076 33684
rect 76132 33628 76142 33684
rect 0 33572 800 33600
rect 76076 33572 76132 33628
rect 79200 33572 80000 33600
rect 0 33516 1932 33572
rect 1988 33516 1998 33572
rect 3714 33516 3724 33572
rect 3780 33516 69580 33572
rect 69636 33516 69646 33572
rect 76076 33516 80000 33572
rect 0 33488 800 33516
rect 79200 33488 80000 33516
rect 3154 33404 3164 33460
rect 3220 33404 3612 33460
rect 3668 33404 63868 33460
rect 63924 33404 63934 33460
rect 64082 33404 64092 33460
rect 64148 33404 75628 33460
rect 75684 33404 76412 33460
rect 76468 33404 76478 33460
rect 8978 33292 8988 33348
rect 9044 33292 9660 33348
rect 9716 33292 10332 33348
rect 10388 33292 10398 33348
rect 11442 33292 11452 33348
rect 11508 33292 12012 33348
rect 12068 33292 13804 33348
rect 13860 33292 13870 33348
rect 28242 33292 28252 33348
rect 28308 33292 29932 33348
rect 29988 33292 29998 33348
rect 37314 33292 37324 33348
rect 37380 33292 39340 33348
rect 39396 33292 39406 33348
rect 43138 33292 43148 33348
rect 43204 33292 43484 33348
rect 43540 33292 44268 33348
rect 44324 33292 45612 33348
rect 45668 33292 45678 33348
rect 49634 33292 49644 33348
rect 49700 33292 50092 33348
rect 50148 33292 50428 33348
rect 50484 33292 50494 33348
rect 50978 33292 50988 33348
rect 51044 33292 52556 33348
rect 52612 33292 53116 33348
rect 53172 33292 53182 33348
rect 56578 33292 56588 33348
rect 56644 33292 57484 33348
rect 57540 33292 57708 33348
rect 57764 33292 57774 33348
rect 64194 33292 64204 33348
rect 64260 33292 65436 33348
rect 65492 33292 66556 33348
rect 66612 33292 66622 33348
rect 68450 33292 68460 33348
rect 68516 33292 73948 33348
rect 74004 33292 77308 33348
rect 77364 33292 77374 33348
rect 13122 33180 13132 33236
rect 13188 33180 13692 33236
rect 13748 33180 13758 33236
rect 43922 33180 43932 33236
rect 43988 33180 45500 33236
rect 45556 33180 45566 33236
rect 45826 33180 45836 33236
rect 45892 33180 46060 33236
rect 46116 33180 51548 33236
rect 51604 33180 51614 33236
rect 51762 33180 51772 33236
rect 51828 33180 52332 33236
rect 52388 33180 52398 33236
rect 53890 33180 53900 33236
rect 53956 33180 57148 33236
rect 57204 33180 57214 33236
rect 63186 33180 63196 33236
rect 63252 33180 63980 33236
rect 64036 33180 64046 33236
rect 69234 33180 69244 33236
rect 69300 33180 72436 33236
rect 72380 33124 72436 33180
rect 7634 33068 7644 33124
rect 7700 33068 9436 33124
rect 9492 33068 9502 33124
rect 12338 33068 12348 33124
rect 12404 33068 19964 33124
rect 20020 33068 21028 33124
rect 27010 33068 27020 33124
rect 27076 33068 28476 33124
rect 28532 33068 29820 33124
rect 29876 33068 29886 33124
rect 31826 33068 31836 33124
rect 31892 33068 36876 33124
rect 36932 33068 37996 33124
rect 38052 33068 38556 33124
rect 38612 33068 39228 33124
rect 39284 33068 39294 33124
rect 44706 33068 44716 33124
rect 44772 33068 50652 33124
rect 50708 33068 50988 33124
rect 51044 33068 51054 33124
rect 51650 33068 51660 33124
rect 51716 33068 52780 33124
rect 52836 33068 52846 33124
rect 60610 33068 60620 33124
rect 60676 33068 61516 33124
rect 61572 33068 61582 33124
rect 67218 33068 67228 33124
rect 67284 33068 70588 33124
rect 70644 33068 71932 33124
rect 71988 33068 71998 33124
rect 72370 33068 72380 33124
rect 72436 33068 74844 33124
rect 74900 33068 74910 33124
rect 20522 32900 20532 32956
rect 20588 32900 20636 32956
rect 20692 32900 20740 32956
rect 20796 32900 20806 32956
rect 20972 32900 21028 33068
rect 44370 32956 44380 33012
rect 44436 32956 48412 33012
rect 48468 32956 48478 33012
rect 39842 32900 39852 32956
rect 39908 32900 39956 32956
rect 40012 32900 40060 32956
rect 40116 32900 40126 32956
rect 59162 32900 59172 32956
rect 59228 32900 59276 32956
rect 59332 32900 59380 32956
rect 59436 32900 59446 32956
rect 78482 32900 78492 32956
rect 78548 32900 78596 32956
rect 78652 32900 78700 32956
rect 78756 32900 78766 32956
rect 7420 32844 8316 32900
rect 8372 32844 8382 32900
rect 20972 32844 31948 32900
rect 7420 32788 7476 32844
rect 31892 32788 31948 32844
rect 44268 32844 55468 32900
rect 44268 32788 44324 32844
rect 55412 32788 55468 32844
rect 67172 32844 77532 32900
rect 77588 32844 78092 32900
rect 78148 32844 78158 32900
rect 67172 32788 67228 32844
rect 6738 32732 6748 32788
rect 6804 32732 7420 32788
rect 7476 32732 7486 32788
rect 8194 32732 8204 32788
rect 8260 32732 9884 32788
rect 9940 32732 9950 32788
rect 31892 32732 44324 32788
rect 48066 32732 48076 32788
rect 48132 32732 50764 32788
rect 50820 32732 50830 32788
rect 55412 32732 67228 32788
rect 74274 32732 74284 32788
rect 74340 32732 75740 32788
rect 75796 32732 75806 32788
rect 7298 32620 7308 32676
rect 7364 32620 8092 32676
rect 8148 32620 8158 32676
rect 8306 32620 8316 32676
rect 8372 32620 10108 32676
rect 10164 32620 10174 32676
rect 15250 32620 15260 32676
rect 15316 32620 22652 32676
rect 22708 32620 44492 32676
rect 44548 32620 44558 32676
rect 52210 32620 52220 32676
rect 52276 32620 53788 32676
rect 53844 32620 53854 32676
rect 55412 32620 58156 32676
rect 58212 32620 59276 32676
rect 59332 32620 59836 32676
rect 59892 32620 59902 32676
rect 65650 32620 65660 32676
rect 65716 32620 67452 32676
rect 67508 32620 69356 32676
rect 69412 32620 69422 32676
rect 77522 32620 77532 32676
rect 77588 32620 77980 32676
rect 78036 32620 78046 32676
rect 7644 32564 7700 32620
rect 7634 32508 7644 32564
rect 7700 32508 7710 32564
rect 13010 32508 13020 32564
rect 13076 32508 14028 32564
rect 14084 32508 14252 32564
rect 14308 32508 14318 32564
rect 19058 32508 19068 32564
rect 19124 32508 20300 32564
rect 20356 32508 20366 32564
rect 24098 32508 24108 32564
rect 24164 32508 27468 32564
rect 27524 32508 28924 32564
rect 28980 32508 28990 32564
rect 33394 32508 33404 32564
rect 33460 32508 33852 32564
rect 33908 32508 33918 32564
rect 46498 32508 46508 32564
rect 46564 32508 49532 32564
rect 49588 32508 49598 32564
rect 55412 32452 55468 32620
rect 55682 32508 55692 32564
rect 55748 32508 56364 32564
rect 56420 32508 56430 32564
rect 60050 32508 60060 32564
rect 60116 32508 60508 32564
rect 60564 32508 61516 32564
rect 61572 32508 61582 32564
rect 62178 32508 62188 32564
rect 62244 32508 63196 32564
rect 63252 32508 63262 32564
rect 66770 32508 66780 32564
rect 66836 32508 67564 32564
rect 67620 32508 70700 32564
rect 70756 32508 70766 32564
rect 73378 32508 73388 32564
rect 73444 32508 74844 32564
rect 74900 32508 74910 32564
rect 7186 32396 7196 32452
rect 7252 32396 8540 32452
rect 8596 32396 8988 32452
rect 9044 32396 9054 32452
rect 13234 32396 13244 32452
rect 13300 32396 14140 32452
rect 14196 32396 14206 32452
rect 23426 32396 23436 32452
rect 23492 32396 23996 32452
rect 24052 32396 24062 32452
rect 31378 32396 31388 32452
rect 31444 32396 37100 32452
rect 37156 32396 37548 32452
rect 37604 32396 37614 32452
rect 53778 32396 53788 32452
rect 53844 32396 55468 32452
rect 55692 32340 55748 32508
rect 61618 32396 61628 32452
rect 61684 32396 62636 32452
rect 62692 32396 62702 32452
rect 27570 32284 27580 32340
rect 27636 32284 29148 32340
rect 29204 32284 29214 32340
rect 52322 32284 52332 32340
rect 52388 32284 55748 32340
rect 38098 32172 38108 32228
rect 38164 32172 38780 32228
rect 38836 32172 38846 32228
rect 10862 32116 10872 32172
rect 10928 32116 10976 32172
rect 11032 32116 11080 32172
rect 11136 32116 11146 32172
rect 30182 32116 30192 32172
rect 30248 32116 30296 32172
rect 30352 32116 30400 32172
rect 30456 32116 30466 32172
rect 49502 32116 49512 32172
rect 49568 32116 49616 32172
rect 49672 32116 49720 32172
rect 49776 32116 49786 32172
rect 68822 32116 68832 32172
rect 68888 32116 68936 32172
rect 68992 32116 69040 32172
rect 69096 32116 69106 32172
rect 31154 31948 31164 32004
rect 31220 31948 31612 32004
rect 31668 31948 31678 32004
rect 32162 31948 32172 32004
rect 32228 31948 33404 32004
rect 33460 31948 33470 32004
rect 37314 31948 37324 32004
rect 37380 31948 37772 32004
rect 37828 31948 37838 32004
rect 54114 31948 54124 32004
rect 54180 31948 54572 32004
rect 54628 31948 55356 32004
rect 55412 31948 55422 32004
rect 57586 31948 57596 32004
rect 57652 31948 59164 32004
rect 59220 31948 59500 32004
rect 59556 31948 60284 32004
rect 60340 31948 60350 32004
rect 4946 31836 4956 31892
rect 5012 31836 5628 31892
rect 5684 31836 5694 31892
rect 5852 31836 65884 31892
rect 65940 31836 65950 31892
rect 76626 31836 76636 31892
rect 76692 31836 77308 31892
rect 77364 31836 77374 31892
rect 5852 31668 5908 31836
rect 8754 31724 8764 31780
rect 8820 31724 9324 31780
rect 9380 31724 10444 31780
rect 10500 31724 10510 31780
rect 14130 31724 14140 31780
rect 14196 31724 14812 31780
rect 14868 31724 14878 31780
rect 20626 31724 20636 31780
rect 20692 31724 21756 31780
rect 21812 31724 21822 31780
rect 40450 31724 40460 31780
rect 40516 31724 41020 31780
rect 41076 31724 41086 31780
rect 45378 31724 45388 31780
rect 45444 31724 46620 31780
rect 46676 31724 46686 31780
rect 46946 31724 46956 31780
rect 47012 31724 47628 31780
rect 47684 31724 47694 31780
rect 49298 31724 49308 31780
rect 49364 31724 49980 31780
rect 50036 31724 50046 31780
rect 55570 31724 55580 31780
rect 55636 31724 56140 31780
rect 56196 31724 56206 31780
rect 58482 31724 58492 31780
rect 58548 31724 59500 31780
rect 59556 31724 60284 31780
rect 60340 31724 60350 31780
rect 61842 31724 61852 31780
rect 61908 31724 62300 31780
rect 62356 31724 62366 31780
rect 67554 31724 67564 31780
rect 67620 31724 69804 31780
rect 69860 31724 69870 31780
rect 77522 31724 77532 31780
rect 77588 31724 78204 31780
rect 78260 31724 78270 31780
rect 3042 31612 3052 31668
rect 3108 31612 3500 31668
rect 3556 31612 5908 31668
rect 6178 31612 6188 31668
rect 6244 31612 8428 31668
rect 15698 31612 15708 31668
rect 15764 31612 16156 31668
rect 16212 31612 16222 31668
rect 20850 31612 20860 31668
rect 20916 31612 21980 31668
rect 22036 31612 22046 31668
rect 8372 31556 8428 31612
rect 46620 31556 46676 31724
rect 46834 31612 46844 31668
rect 46900 31612 47292 31668
rect 47348 31612 47358 31668
rect 51090 31612 51100 31668
rect 51156 31612 52220 31668
rect 52276 31612 54012 31668
rect 54068 31612 54078 31668
rect 56802 31612 56812 31668
rect 56868 31612 59724 31668
rect 59780 31612 60396 31668
rect 60452 31612 60462 31668
rect 68226 31612 68236 31668
rect 68292 31612 69580 31668
rect 69636 31612 69646 31668
rect 71250 31612 71260 31668
rect 71316 31612 77420 31668
rect 77476 31612 77486 31668
rect 4162 31500 4172 31556
rect 4228 31500 6076 31556
rect 6132 31500 6142 31556
rect 8372 31500 23548 31556
rect 23604 31500 24556 31556
rect 24612 31500 24622 31556
rect 27682 31500 27692 31556
rect 27748 31500 33180 31556
rect 33236 31500 33516 31556
rect 33572 31500 33582 31556
rect 46620 31500 47516 31556
rect 47572 31500 47852 31556
rect 47908 31500 48076 31556
rect 48132 31500 48142 31556
rect 51202 31500 51212 31556
rect 51268 31500 51772 31556
rect 51828 31500 51838 31556
rect 52770 31500 52780 31556
rect 52836 31500 53900 31556
rect 53956 31500 53966 31556
rect 55906 31500 55916 31556
rect 55972 31500 57260 31556
rect 57316 31500 58268 31556
rect 58324 31500 58716 31556
rect 58772 31500 58782 31556
rect 63634 31500 63644 31556
rect 63700 31500 65436 31556
rect 65492 31500 65502 31556
rect 65762 31500 65772 31556
rect 65828 31500 67340 31556
rect 67396 31500 71036 31556
rect 71092 31500 71820 31556
rect 71876 31500 71886 31556
rect 74386 31500 74396 31556
rect 74452 31500 75404 31556
rect 75460 31500 77532 31556
rect 77588 31500 77598 31556
rect 51772 31444 51828 31500
rect 4722 31388 4732 31444
rect 4788 31388 6300 31444
rect 6356 31388 6366 31444
rect 8372 31388 20188 31444
rect 20244 31388 20254 31444
rect 43148 31388 44380 31444
rect 44436 31388 44446 31444
rect 51772 31388 53788 31444
rect 53844 31388 53854 31444
rect 56354 31388 56364 31444
rect 56420 31388 57708 31444
rect 57764 31388 57774 31444
rect 66770 31388 66780 31444
rect 66836 31388 67228 31444
rect 67284 31388 68460 31444
rect 68516 31388 68526 31444
rect 71922 31388 71932 31444
rect 71988 31388 72268 31444
rect 72324 31388 72334 31444
rect 8372 31332 8428 31388
rect 20522 31332 20532 31388
rect 20588 31332 20636 31388
rect 20692 31332 20740 31388
rect 20796 31332 20806 31388
rect 39842 31332 39852 31388
rect 39908 31332 39956 31388
rect 40012 31332 40060 31388
rect 40116 31332 40126 31388
rect 5954 31276 5964 31332
rect 6020 31276 8428 31332
rect 14354 31276 14364 31332
rect 14420 31276 14924 31332
rect 14980 31276 17052 31332
rect 17108 31276 17118 31332
rect 43148 31220 43204 31388
rect 59162 31332 59172 31388
rect 59228 31332 59276 31388
rect 59332 31332 59380 31388
rect 59436 31332 59446 31388
rect 78482 31332 78492 31388
rect 78548 31332 78596 31388
rect 78652 31332 78700 31388
rect 78756 31332 78766 31388
rect 44482 31276 44492 31332
rect 44548 31276 50428 31332
rect 73490 31276 73500 31332
rect 73556 31276 74676 31332
rect 50372 31220 50428 31276
rect 74620 31220 74676 31276
rect 1586 31164 1596 31220
rect 1652 31164 10836 31220
rect 12786 31164 12796 31220
rect 12852 31164 13468 31220
rect 13524 31164 13534 31220
rect 14690 31164 14700 31220
rect 14756 31164 15596 31220
rect 15652 31164 15662 31220
rect 16594 31164 16604 31220
rect 16660 31164 24220 31220
rect 24276 31164 24286 31220
rect 26898 31164 26908 31220
rect 26964 31164 27804 31220
rect 27860 31164 27870 31220
rect 31892 31164 43204 31220
rect 44146 31164 44156 31220
rect 44212 31164 46396 31220
rect 46452 31164 46462 31220
rect 50372 31164 67228 31220
rect 69570 31164 69580 31220
rect 69636 31164 70812 31220
rect 70868 31164 70878 31220
rect 71922 31164 71932 31220
rect 71988 31164 73388 31220
rect 73444 31164 73454 31220
rect 74610 31164 74620 31220
rect 74676 31164 76300 31220
rect 76356 31164 76366 31220
rect 0 31108 800 31136
rect 10780 31108 10836 31164
rect 31892 31108 31948 31164
rect 67172 31108 67228 31164
rect 79200 31108 80000 31136
rect 0 31052 1932 31108
rect 1988 31052 1998 31108
rect 8194 31052 8204 31108
rect 8260 31052 8652 31108
rect 8708 31052 8718 31108
rect 10780 31052 31948 31108
rect 39330 31052 39340 31108
rect 39396 31052 40460 31108
rect 40516 31052 40526 31108
rect 42018 31052 42028 31108
rect 42084 31052 43596 31108
rect 43652 31052 43662 31108
rect 49746 31052 49756 31108
rect 49812 31052 50428 31108
rect 50484 31052 50494 31108
rect 54002 31052 54012 31108
rect 54068 31052 55356 31108
rect 55412 31052 55422 31108
rect 67172 31052 74116 31108
rect 75506 31052 75516 31108
rect 75572 31052 80000 31108
rect 0 31024 800 31052
rect 74060 30996 74116 31052
rect 79200 31024 80000 31052
rect 4498 30940 4508 30996
rect 4564 30940 6972 30996
rect 7028 30940 7038 30996
rect 12450 30940 12460 30996
rect 12516 30940 13804 30996
rect 13860 30940 13870 30996
rect 14914 30940 14924 30996
rect 14980 30940 18732 30996
rect 18788 30940 19964 30996
rect 20020 30940 20030 30996
rect 26338 30940 26348 30996
rect 26404 30940 27244 30996
rect 27300 30940 27310 30996
rect 29586 30940 29596 30996
rect 29652 30940 30492 30996
rect 30548 30940 31612 30996
rect 31668 30940 31678 30996
rect 39666 30940 39676 30996
rect 39732 30940 42140 30996
rect 42196 30940 42206 30996
rect 51426 30940 51436 30996
rect 51492 30940 54236 30996
rect 54292 30940 54302 30996
rect 66098 30940 66108 30996
rect 66164 30940 67564 30996
rect 67620 30940 67630 30996
rect 68562 30940 68572 30996
rect 68628 30940 69132 30996
rect 69188 30940 71708 30996
rect 71764 30940 71774 30996
rect 74060 30940 77084 30996
rect 77140 30940 77644 30996
rect 77700 30940 77710 30996
rect 8978 30828 8988 30884
rect 9044 30828 10332 30884
rect 10388 30828 10398 30884
rect 16706 30828 16716 30884
rect 16772 30828 17612 30884
rect 17668 30828 17678 30884
rect 39106 30828 39116 30884
rect 39172 30828 40236 30884
rect 40292 30828 40302 30884
rect 46162 30828 46172 30884
rect 46228 30828 46956 30884
rect 47012 30828 47022 30884
rect 51538 30828 51548 30884
rect 51604 30828 52444 30884
rect 52500 30828 52510 30884
rect 54674 30828 54684 30884
rect 54740 30828 55580 30884
rect 55636 30828 55646 30884
rect 62290 30828 62300 30884
rect 62356 30828 63868 30884
rect 63924 30828 64316 30884
rect 64372 30828 64382 30884
rect 30594 30716 30604 30772
rect 30660 30716 32060 30772
rect 32116 30716 32126 30772
rect 37874 30716 37884 30772
rect 37940 30716 39340 30772
rect 39396 30716 39406 30772
rect 42130 30716 42140 30772
rect 42196 30716 45388 30772
rect 45444 30716 45948 30772
rect 46004 30716 46014 30772
rect 54226 30716 54236 30772
rect 54292 30716 54796 30772
rect 54852 30716 54862 30772
rect 55458 30716 55468 30772
rect 55524 30716 55916 30772
rect 55972 30716 55982 30772
rect 63298 30716 63308 30772
rect 63364 30716 66108 30772
rect 66164 30716 66174 30772
rect 72034 30716 72044 30772
rect 72100 30716 75964 30772
rect 76020 30716 77308 30772
rect 77364 30716 77374 30772
rect 19170 30604 19180 30660
rect 19236 30604 19740 30660
rect 19796 30604 19806 30660
rect 34514 30604 34524 30660
rect 34580 30604 36428 30660
rect 36484 30604 36494 30660
rect 50978 30604 50988 30660
rect 51044 30604 59724 30660
rect 59780 30604 60172 30660
rect 60228 30604 61964 30660
rect 62020 30604 62030 30660
rect 10862 30548 10872 30604
rect 10928 30548 10976 30604
rect 11032 30548 11080 30604
rect 11136 30548 11146 30604
rect 30182 30548 30192 30604
rect 30248 30548 30296 30604
rect 30352 30548 30400 30604
rect 30456 30548 30466 30604
rect 49502 30548 49512 30604
rect 49568 30548 49616 30604
rect 49672 30548 49720 30604
rect 49776 30548 49786 30604
rect 68822 30548 68832 30604
rect 68888 30548 68936 30604
rect 68992 30548 69040 30604
rect 69096 30548 69106 30604
rect 10658 30492 10668 30548
rect 10724 30492 10734 30548
rect 55346 30492 55356 30548
rect 55468 30492 55488 30548
rect 55580 30492 60732 30548
rect 60788 30492 60798 30548
rect 10668 30436 10724 30492
rect 55580 30436 55636 30492
rect 8642 30380 8652 30436
rect 8708 30380 9436 30436
rect 9492 30380 9884 30436
rect 9940 30380 11900 30436
rect 11956 30380 13692 30436
rect 13748 30380 13758 30436
rect 17602 30380 17612 30436
rect 17668 30380 18732 30436
rect 18788 30380 18798 30436
rect 20132 30380 55636 30436
rect 20132 30324 20188 30380
rect 10322 30268 10332 30324
rect 10388 30268 10668 30324
rect 10724 30268 11564 30324
rect 11620 30268 11630 30324
rect 16828 30268 20188 30324
rect 24994 30268 25004 30324
rect 25060 30268 25340 30324
rect 25396 30268 26012 30324
rect 26068 30268 26078 30324
rect 30258 30268 30268 30324
rect 30324 30268 32284 30324
rect 32340 30268 32350 30324
rect 33730 30268 33740 30324
rect 33796 30268 34524 30324
rect 34580 30268 34590 30324
rect 35410 30268 35420 30324
rect 35476 30268 39116 30324
rect 39172 30268 39182 30324
rect 48738 30268 48748 30324
rect 48804 30268 49756 30324
rect 49812 30268 49822 30324
rect 53554 30268 53564 30324
rect 53620 30268 55692 30324
rect 55748 30268 56364 30324
rect 56420 30268 56430 30324
rect 68450 30268 68460 30324
rect 68516 30268 68526 30324
rect 69458 30268 69468 30324
rect 69524 30268 70812 30324
rect 70868 30268 70878 30324
rect 74386 30268 74396 30324
rect 74452 30268 75404 30324
rect 75460 30268 75470 30324
rect 10546 30156 10556 30212
rect 10612 30156 11788 30212
rect 11844 30156 11854 30212
rect 16828 30100 16884 30268
rect 29362 30156 29372 30212
rect 29428 30156 30044 30212
rect 30100 30156 30604 30212
rect 30660 30156 30670 30212
rect 34738 30156 34748 30212
rect 34804 30156 35308 30212
rect 35364 30156 35374 30212
rect 36642 30156 36652 30212
rect 36708 30156 37436 30212
rect 37492 30156 37502 30212
rect 44706 30156 44716 30212
rect 44772 30156 46060 30212
rect 46116 30156 46126 30212
rect 54572 30100 54628 30268
rect 68460 30212 68516 30268
rect 54786 30156 54796 30212
rect 54852 30156 55916 30212
rect 55972 30156 57148 30212
rect 57204 30156 57214 30212
rect 62066 30156 62076 30212
rect 62132 30156 62524 30212
rect 62580 30156 66108 30212
rect 66164 30156 66174 30212
rect 68460 30156 69748 30212
rect 71138 30156 71148 30212
rect 71204 30156 72156 30212
rect 72212 30156 75068 30212
rect 75124 30156 75134 30212
rect 75506 30156 75516 30212
rect 75572 30156 76076 30212
rect 76132 30156 77868 30212
rect 77924 30156 77934 30212
rect 69692 30100 69748 30156
rect 75516 30100 75572 30156
rect 6626 30044 6636 30100
rect 6692 30044 6860 30100
rect 6916 30044 6926 30100
rect 8866 30044 8876 30100
rect 8932 30044 9548 30100
rect 9604 30044 10444 30100
rect 10500 30044 10510 30100
rect 14252 30044 16884 30100
rect 31602 30044 31612 30100
rect 31668 30044 32172 30100
rect 32228 30044 32238 30100
rect 33954 30044 33964 30100
rect 34020 30044 39004 30100
rect 39060 30044 41692 30100
rect 41748 30044 41758 30100
rect 47170 30044 47180 30100
rect 47236 30044 47740 30100
rect 47796 30044 47806 30100
rect 54572 30044 54684 30100
rect 54740 30044 54750 30100
rect 55682 30044 55692 30100
rect 55748 30044 56140 30100
rect 56196 30044 58940 30100
rect 58996 30044 60844 30100
rect 60900 30044 60910 30100
rect 67778 30044 67788 30100
rect 67844 30044 68460 30100
rect 68516 30044 69468 30100
rect 69524 30044 69534 30100
rect 69682 30044 69692 30100
rect 69748 30044 72716 30100
rect 72772 30044 72782 30100
rect 74946 30044 74956 30100
rect 75012 30044 75572 30100
rect 76514 30044 76524 30100
rect 76580 30044 77756 30100
rect 77812 30044 77822 30100
rect 14252 29988 14308 30044
rect 76524 29988 76580 30044
rect 2370 29932 2380 29988
rect 2436 29932 3164 29988
rect 3220 29932 14308 29988
rect 15474 29932 15484 29988
rect 15540 29932 22988 29988
rect 23044 29932 23436 29988
rect 23492 29932 24108 29988
rect 24164 29932 24174 29988
rect 25106 29932 25116 29988
rect 25172 29932 28812 29988
rect 28868 29932 30268 29988
rect 30324 29932 30334 29988
rect 34066 29932 34076 29988
rect 34132 29932 34636 29988
rect 34692 29932 36092 29988
rect 36148 29932 36540 29988
rect 36596 29932 36606 29988
rect 40898 29932 40908 29988
rect 40964 29932 41356 29988
rect 41412 29932 43148 29988
rect 43204 29932 43214 29988
rect 55570 29932 55580 29988
rect 55636 29932 56700 29988
rect 56756 29932 56766 29988
rect 66994 29932 67004 29988
rect 67060 29932 67900 29988
rect 67956 29932 67966 29988
rect 70802 29932 70812 29988
rect 70868 29932 71820 29988
rect 71876 29932 71886 29988
rect 74162 29932 74172 29988
rect 74228 29932 76580 29988
rect 5394 29820 5404 29876
rect 5460 29820 12908 29876
rect 12964 29820 13916 29876
rect 13972 29820 14812 29876
rect 14868 29820 14878 29876
rect 44482 29820 44492 29876
rect 44548 29820 53452 29876
rect 53508 29820 54012 29876
rect 54068 29820 54796 29876
rect 54852 29820 56252 29876
rect 56308 29820 58044 29876
rect 58100 29820 58110 29876
rect 74274 29820 74284 29876
rect 74340 29820 74844 29876
rect 74900 29820 76188 29876
rect 76244 29820 77532 29876
rect 77588 29820 77598 29876
rect 20522 29764 20532 29820
rect 20588 29764 20636 29820
rect 20692 29764 20740 29820
rect 20796 29764 20806 29820
rect 39842 29764 39852 29820
rect 39908 29764 39956 29820
rect 40012 29764 40060 29820
rect 40116 29764 40126 29820
rect 59162 29764 59172 29820
rect 59228 29764 59276 29820
rect 59332 29764 59380 29820
rect 59436 29764 59446 29820
rect 78482 29764 78492 29820
rect 78548 29764 78596 29820
rect 78652 29764 78700 29820
rect 78756 29764 78766 29820
rect 1474 29708 1484 29764
rect 1540 29708 20188 29764
rect 26898 29708 26908 29764
rect 26964 29708 27356 29764
rect 27412 29708 28588 29764
rect 28644 29708 29820 29764
rect 29876 29708 29886 29764
rect 71810 29708 71820 29764
rect 71876 29708 75068 29764
rect 75124 29708 75134 29764
rect 20132 29652 20188 29708
rect 6402 29596 6412 29652
rect 6468 29596 8428 29652
rect 10994 29596 11004 29652
rect 11060 29596 12124 29652
rect 12180 29596 12190 29652
rect 16034 29596 16044 29652
rect 16100 29596 16380 29652
rect 16436 29596 17164 29652
rect 17220 29596 17230 29652
rect 20132 29596 36820 29652
rect 40450 29596 40460 29652
rect 40516 29596 44604 29652
rect 44660 29596 45276 29652
rect 45332 29596 45342 29652
rect 50418 29596 50428 29652
rect 50484 29596 51100 29652
rect 51156 29596 51166 29652
rect 52434 29596 52444 29652
rect 52500 29596 52510 29652
rect 59826 29596 59836 29652
rect 59892 29596 60732 29652
rect 60788 29596 60798 29652
rect 4610 29484 4620 29540
rect 4676 29484 6972 29540
rect 7028 29484 7038 29540
rect 4162 29372 4172 29428
rect 4228 29372 4844 29428
rect 4900 29372 4910 29428
rect 8372 29204 8428 29596
rect 36764 29540 36820 29596
rect 18274 29484 18284 29540
rect 18340 29484 18844 29540
rect 18900 29484 18910 29540
rect 26898 29484 26908 29540
rect 26964 29484 27468 29540
rect 27524 29484 27534 29540
rect 33058 29484 33068 29540
rect 33124 29484 33628 29540
rect 33684 29484 33694 29540
rect 36764 29484 45500 29540
rect 45556 29484 46508 29540
rect 46564 29484 46574 29540
rect 52444 29428 52500 29596
rect 54898 29484 54908 29540
rect 54964 29484 60620 29540
rect 60676 29484 61628 29540
rect 61684 29484 61694 29540
rect 67890 29484 67900 29540
rect 67956 29484 68236 29540
rect 68292 29484 69580 29540
rect 69636 29484 69646 29540
rect 11442 29372 11452 29428
rect 11508 29372 12348 29428
rect 12404 29372 12414 29428
rect 21298 29372 21308 29428
rect 21364 29372 22428 29428
rect 22484 29372 22494 29428
rect 23090 29372 23100 29428
rect 23156 29372 23660 29428
rect 23716 29372 23726 29428
rect 23986 29372 23996 29428
rect 24052 29372 24220 29428
rect 24276 29372 26628 29428
rect 28802 29372 28812 29428
rect 28868 29372 32396 29428
rect 32452 29372 32462 29428
rect 40562 29372 40572 29428
rect 40628 29372 40796 29428
rect 40852 29372 41804 29428
rect 41860 29372 41870 29428
rect 46834 29372 46844 29428
rect 46900 29372 49644 29428
rect 49700 29372 49710 29428
rect 52444 29372 54572 29428
rect 54628 29372 56028 29428
rect 56084 29372 56094 29428
rect 56242 29372 56252 29428
rect 56308 29372 56812 29428
rect 56868 29372 57372 29428
rect 57428 29372 57438 29428
rect 58594 29372 58604 29428
rect 58660 29372 59500 29428
rect 59556 29372 59566 29428
rect 70802 29372 70812 29428
rect 70868 29372 71372 29428
rect 71428 29372 71438 29428
rect 26572 29316 26628 29372
rect 11330 29260 11340 29316
rect 11396 29260 12124 29316
rect 12180 29260 12460 29316
rect 12516 29260 12908 29316
rect 12964 29260 12974 29316
rect 21522 29260 21532 29316
rect 21588 29260 22204 29316
rect 22260 29260 22876 29316
rect 22932 29260 22942 29316
rect 24546 29260 24556 29316
rect 24612 29260 26348 29316
rect 26404 29260 26414 29316
rect 26572 29260 31948 29316
rect 32722 29260 32732 29316
rect 32788 29260 35532 29316
rect 35588 29260 35598 29316
rect 37986 29260 37996 29316
rect 38052 29260 39116 29316
rect 39172 29260 41132 29316
rect 41188 29260 41692 29316
rect 41748 29260 41758 29316
rect 56578 29260 56588 29316
rect 56644 29260 58156 29316
rect 58212 29260 58222 29316
rect 59714 29260 59724 29316
rect 59780 29260 60284 29316
rect 60340 29260 60350 29316
rect 66770 29260 66780 29316
rect 66836 29260 67340 29316
rect 67396 29260 68572 29316
rect 68628 29260 68638 29316
rect 31892 29204 31948 29260
rect 8372 29148 21756 29204
rect 21812 29148 21822 29204
rect 31892 29148 35756 29204
rect 35812 29148 35822 29204
rect 38546 29148 38556 29204
rect 38612 29148 39340 29204
rect 39396 29148 39406 29204
rect 48738 29148 48748 29204
rect 48804 29148 49868 29204
rect 49924 29148 51324 29204
rect 51380 29148 51390 29204
rect 51874 29148 51884 29204
rect 51940 29148 52668 29204
rect 52724 29148 52734 29204
rect 55412 29148 72380 29204
rect 72436 29148 72446 29204
rect 15362 29036 15372 29092
rect 15428 29036 23548 29092
rect 23604 29036 23614 29092
rect 10862 28980 10872 29036
rect 10928 28980 10976 29036
rect 11032 28980 11080 29036
rect 11136 28980 11146 29036
rect 30182 28980 30192 29036
rect 30248 28980 30296 29036
rect 30352 28980 30400 29036
rect 30456 28980 30466 29036
rect 49502 28980 49512 29036
rect 49568 28980 49616 29036
rect 49672 28980 49720 29036
rect 49776 28980 49786 29036
rect 15474 28924 15484 28980
rect 15540 28924 27356 28980
rect 27412 28924 27422 28980
rect 55412 28868 55468 29148
rect 68822 28980 68832 29036
rect 68888 28980 68936 29036
rect 68992 28980 69040 29036
rect 69096 28980 69106 29036
rect 76962 28924 76972 28980
rect 77028 28924 77924 28980
rect 77868 28868 77924 28924
rect 3602 28812 3612 28868
rect 3668 28812 55468 28868
rect 63858 28812 63868 28868
rect 63924 28812 65996 28868
rect 66052 28812 66062 28868
rect 70018 28812 70028 28868
rect 70084 28812 73836 28868
rect 73892 28812 73902 28868
rect 74498 28812 74508 28868
rect 74564 28812 77308 28868
rect 77364 28812 77374 28868
rect 77858 28812 77868 28868
rect 77924 28812 77934 28868
rect 5058 28700 5068 28756
rect 5124 28700 10388 28756
rect 17826 28700 17836 28756
rect 17892 28700 18956 28756
rect 19012 28700 19022 28756
rect 24770 28700 24780 28756
rect 24836 28700 25564 28756
rect 25620 28700 25630 28756
rect 39330 28700 39340 28756
rect 39396 28700 40012 28756
rect 40068 28700 40908 28756
rect 40964 28700 40974 28756
rect 45378 28700 45388 28756
rect 45444 28700 46620 28756
rect 46676 28700 48188 28756
rect 48244 28700 48412 28756
rect 48468 28700 48478 28756
rect 50530 28700 50540 28756
rect 50596 28700 52332 28756
rect 52388 28700 53004 28756
rect 53060 28700 53070 28756
rect 65090 28700 65100 28756
rect 65156 28700 65772 28756
rect 65828 28700 65838 28756
rect 75506 28700 75516 28756
rect 75572 28700 76300 28756
rect 76356 28700 77644 28756
rect 77700 28700 77710 28756
rect 77942 28700 77980 28756
rect 78036 28700 78046 28756
rect 0 28644 800 28672
rect 0 28588 1932 28644
rect 1988 28588 1998 28644
rect 7298 28588 7308 28644
rect 7364 28588 7756 28644
rect 7812 28588 7980 28644
rect 8036 28588 9884 28644
rect 9940 28588 9950 28644
rect 0 28560 800 28588
rect 3154 28476 3164 28532
rect 3220 28476 3612 28532
rect 3668 28476 3678 28532
rect 10332 28420 10388 28700
rect 79200 28644 80000 28672
rect 13804 28588 15372 28644
rect 15428 28588 15438 28644
rect 18610 28588 18620 28644
rect 18676 28588 19180 28644
rect 19236 28588 19246 28644
rect 28466 28588 28476 28644
rect 28532 28588 29708 28644
rect 29764 28588 29774 28644
rect 31042 28588 31052 28644
rect 31108 28588 31612 28644
rect 31668 28588 32508 28644
rect 32564 28588 33740 28644
rect 33796 28588 34300 28644
rect 34356 28588 34366 28644
rect 36866 28588 36876 28644
rect 36932 28588 37436 28644
rect 37492 28588 37502 28644
rect 46386 28588 46396 28644
rect 46452 28588 48076 28644
rect 48132 28588 48300 28644
rect 48356 28588 48366 28644
rect 48626 28588 48636 28644
rect 48692 28588 51436 28644
rect 51492 28588 51502 28644
rect 56690 28588 56700 28644
rect 56756 28588 58268 28644
rect 58324 28588 58334 28644
rect 65874 28588 65884 28644
rect 65940 28588 66668 28644
rect 66724 28588 67340 28644
rect 67396 28588 67406 28644
rect 70018 28588 70028 28644
rect 70084 28588 70812 28644
rect 70868 28588 71036 28644
rect 71092 28588 71102 28644
rect 72706 28588 72716 28644
rect 72772 28588 75404 28644
rect 75460 28588 75470 28644
rect 76066 28588 76076 28644
rect 76132 28588 80000 28644
rect 13804 28532 13860 28588
rect 79200 28560 80000 28588
rect 13234 28476 13244 28532
rect 13300 28476 13804 28532
rect 13860 28476 13870 28532
rect 17378 28476 17388 28532
rect 17444 28476 19068 28532
rect 19124 28476 19134 28532
rect 23202 28476 23212 28532
rect 23268 28476 23772 28532
rect 23828 28476 23838 28532
rect 25890 28476 25900 28532
rect 25956 28476 26796 28532
rect 26852 28476 26862 28532
rect 28130 28476 28140 28532
rect 28196 28476 28700 28532
rect 28756 28476 29932 28532
rect 29988 28476 29998 28532
rect 32386 28476 32396 28532
rect 32452 28476 33628 28532
rect 33684 28476 33694 28532
rect 40226 28476 40236 28532
rect 40292 28476 44380 28532
rect 44436 28476 45052 28532
rect 45108 28476 45118 28532
rect 53106 28476 53116 28532
rect 53172 28476 54572 28532
rect 54628 28476 54638 28532
rect 58930 28476 58940 28532
rect 58996 28476 59724 28532
rect 59780 28476 61404 28532
rect 61460 28476 61470 28532
rect 68226 28476 68236 28532
rect 68292 28476 69468 28532
rect 69524 28476 69534 28532
rect 77868 28476 78092 28532
rect 78148 28476 78316 28532
rect 78372 28476 78382 28532
rect 77868 28420 77924 28476
rect 3378 28364 3388 28420
rect 3444 28364 4844 28420
rect 4900 28364 6524 28420
rect 6580 28364 6590 28420
rect 10322 28364 10332 28420
rect 10388 28364 10398 28420
rect 12562 28364 12572 28420
rect 12628 28364 13356 28420
rect 13412 28364 17612 28420
rect 17668 28364 17678 28420
rect 17938 28364 17948 28420
rect 18004 28364 18284 28420
rect 18340 28364 20188 28420
rect 20244 28364 20254 28420
rect 24882 28364 24892 28420
rect 24948 28364 25788 28420
rect 25844 28364 27020 28420
rect 27076 28364 27086 28420
rect 27570 28364 27580 28420
rect 27636 28364 28028 28420
rect 28084 28364 28094 28420
rect 35186 28364 35196 28420
rect 35252 28364 35644 28420
rect 35700 28364 35710 28420
rect 36082 28364 36092 28420
rect 36148 28364 36652 28420
rect 36708 28364 36718 28420
rect 37090 28364 37100 28420
rect 37156 28364 38108 28420
rect 38164 28364 38174 28420
rect 54002 28364 54012 28420
rect 54068 28364 54460 28420
rect 54516 28364 55468 28420
rect 55524 28364 55534 28420
rect 59490 28364 59500 28420
rect 59556 28364 60172 28420
rect 60228 28364 61628 28420
rect 61684 28364 61694 28420
rect 77858 28364 77868 28420
rect 77924 28364 77934 28420
rect 35644 28308 35700 28364
rect 21186 28252 21196 28308
rect 21252 28252 25228 28308
rect 25284 28252 25294 28308
rect 35644 28252 36428 28308
rect 36484 28252 36494 28308
rect 77942 28252 77980 28308
rect 78036 28252 78046 28308
rect 20522 28196 20532 28252
rect 20588 28196 20636 28252
rect 20692 28196 20740 28252
rect 20796 28196 20806 28252
rect 39842 28196 39852 28252
rect 39908 28196 39956 28252
rect 40012 28196 40060 28252
rect 40116 28196 40126 28252
rect 59162 28196 59172 28252
rect 59228 28196 59276 28252
rect 59332 28196 59380 28252
rect 59436 28196 59446 28252
rect 78482 28196 78492 28252
rect 78548 28196 78596 28252
rect 78652 28196 78700 28252
rect 78756 28196 78766 28252
rect 14018 28140 14028 28196
rect 14084 28140 14588 28196
rect 14644 28140 14654 28196
rect 22764 28140 24444 28196
rect 24500 28140 24510 28196
rect 47282 28140 47292 28196
rect 47348 28140 53564 28196
rect 53620 28140 54348 28196
rect 54404 28140 54414 28196
rect 76178 28140 76188 28196
rect 76244 28140 76524 28196
rect 76580 28140 76590 28196
rect 77746 28140 77756 28196
rect 77812 28140 78092 28196
rect 78148 28140 78158 28196
rect 22764 28084 22820 28140
rect 5618 28028 5628 28084
rect 5684 28028 22820 28084
rect 22978 28028 22988 28084
rect 23044 28028 23660 28084
rect 23716 28028 23726 28084
rect 35746 28028 35756 28084
rect 35812 28028 79100 28084
rect 79156 28028 79166 28084
rect 14914 27916 14924 27972
rect 14980 27916 15260 27972
rect 15316 27916 15326 27972
rect 27906 27916 27916 27972
rect 27972 27916 28588 27972
rect 28644 27916 28654 27972
rect 30044 27916 30716 27972
rect 30772 27916 30782 27972
rect 45042 27916 45052 27972
rect 45108 27916 45724 27972
rect 45780 27916 46284 27972
rect 46340 27916 46350 27972
rect 52434 27916 52444 27972
rect 52500 27916 54572 27972
rect 54628 27916 54638 27972
rect 56578 27916 56588 27972
rect 56644 27916 56654 27972
rect 57026 27916 57036 27972
rect 57092 27916 59276 27972
rect 59332 27916 59342 27972
rect 59724 27916 60284 27972
rect 60340 27916 60350 27972
rect 60610 27916 60620 27972
rect 60676 27916 61404 27972
rect 61460 27916 64204 27972
rect 64260 27916 64270 27972
rect 65538 27916 65548 27972
rect 65604 27916 65996 27972
rect 66052 27916 66332 27972
rect 66388 27916 67564 27972
rect 67620 27916 67630 27972
rect 74498 27916 74508 27972
rect 74564 27916 75740 27972
rect 75796 27916 76748 27972
rect 76804 27916 77308 27972
rect 77364 27916 77374 27972
rect 30044 27860 30100 27916
rect 56588 27860 56644 27916
rect 59724 27860 59780 27916
rect 3154 27804 3164 27860
rect 3220 27804 4172 27860
rect 4228 27804 5516 27860
rect 5572 27804 5582 27860
rect 10546 27804 10556 27860
rect 10612 27804 13580 27860
rect 13636 27804 14140 27860
rect 14196 27804 14206 27860
rect 15026 27804 15036 27860
rect 15092 27804 15102 27860
rect 21858 27804 21868 27860
rect 21924 27804 22876 27860
rect 22932 27804 24892 27860
rect 24948 27804 24958 27860
rect 26002 27804 26012 27860
rect 26068 27804 26572 27860
rect 26628 27804 26638 27860
rect 27692 27804 30044 27860
rect 30100 27804 30110 27860
rect 30818 27804 30828 27860
rect 30884 27804 31164 27860
rect 31220 27804 31724 27860
rect 31780 27804 31790 27860
rect 45266 27804 45276 27860
rect 45332 27804 45500 27860
rect 45556 27804 46620 27860
rect 46676 27804 46686 27860
rect 46834 27804 46844 27860
rect 46900 27804 57372 27860
rect 57428 27804 57438 27860
rect 58258 27804 58268 27860
rect 58324 27804 58828 27860
rect 58884 27804 59724 27860
rect 59780 27804 59790 27860
rect 60386 27804 60396 27860
rect 60452 27804 61852 27860
rect 61908 27804 62636 27860
rect 62692 27804 62702 27860
rect 74162 27804 74172 27860
rect 74228 27804 76972 27860
rect 77028 27804 77038 27860
rect 15036 27748 15092 27804
rect 27692 27748 27748 27804
rect 4274 27692 4284 27748
rect 4340 27692 4620 27748
rect 4676 27692 4956 27748
rect 5012 27692 5740 27748
rect 5796 27692 6636 27748
rect 6692 27692 7084 27748
rect 7140 27692 12348 27748
rect 12404 27692 12414 27748
rect 13234 27692 13244 27748
rect 13300 27692 15092 27748
rect 25554 27692 25564 27748
rect 25620 27692 27356 27748
rect 27412 27692 27692 27748
rect 27748 27692 27758 27748
rect 28690 27692 28700 27748
rect 28756 27692 35532 27748
rect 35588 27692 36092 27748
rect 36148 27692 36316 27748
rect 36372 27692 36382 27748
rect 40114 27692 40124 27748
rect 40180 27692 41580 27748
rect 41636 27692 41646 27748
rect 46498 27692 46508 27748
rect 46564 27692 48748 27748
rect 48804 27692 49868 27748
rect 49924 27692 49934 27748
rect 50194 27692 50204 27748
rect 50260 27692 52892 27748
rect 52948 27692 54684 27748
rect 54740 27692 54750 27748
rect 58034 27692 58044 27748
rect 58100 27692 59836 27748
rect 59892 27692 64428 27748
rect 64484 27692 64494 27748
rect 10994 27580 11004 27636
rect 11060 27580 14028 27636
rect 14084 27580 14094 27636
rect 16482 27580 16492 27636
rect 16548 27580 17948 27636
rect 18004 27580 22820 27636
rect 30706 27580 30716 27636
rect 30772 27580 31612 27636
rect 31668 27580 31678 27636
rect 39890 27580 39900 27636
rect 39956 27580 41804 27636
rect 41860 27580 41870 27636
rect 45938 27580 45948 27636
rect 46004 27580 46844 27636
rect 46900 27580 49756 27636
rect 49812 27580 49822 27636
rect 58482 27580 58492 27636
rect 58548 27580 59052 27636
rect 59108 27580 59118 27636
rect 22764 27524 22820 27580
rect 22754 27468 22764 27524
rect 22820 27468 22830 27524
rect 41682 27468 41692 27524
rect 41748 27468 46844 27524
rect 46900 27468 46910 27524
rect 69234 27468 69244 27524
rect 69300 27468 71148 27524
rect 71204 27468 71214 27524
rect 74498 27468 74508 27524
rect 74564 27468 75628 27524
rect 75684 27468 76412 27524
rect 76468 27468 77980 27524
rect 78036 27468 78046 27524
rect 10862 27412 10872 27468
rect 10928 27412 10976 27468
rect 11032 27412 11080 27468
rect 11136 27412 11146 27468
rect 30182 27412 30192 27468
rect 30248 27412 30296 27468
rect 30352 27412 30400 27468
rect 30456 27412 30466 27468
rect 49502 27412 49512 27468
rect 49568 27412 49616 27468
rect 49672 27412 49720 27468
rect 49776 27412 49786 27468
rect 68822 27412 68832 27468
rect 68888 27412 68936 27468
rect 68992 27412 69040 27468
rect 69096 27412 69106 27468
rect 23762 27356 23772 27412
rect 23828 27356 29316 27412
rect 29260 27300 29316 27356
rect 31892 27356 42252 27412
rect 42308 27356 42318 27412
rect 31892 27300 31948 27356
rect 8754 27244 8764 27300
rect 8820 27244 10108 27300
rect 10164 27244 10174 27300
rect 14242 27244 14252 27300
rect 14308 27244 15596 27300
rect 15652 27244 20188 27300
rect 28354 27244 28364 27300
rect 28420 27244 29036 27300
rect 29092 27244 29102 27300
rect 29260 27244 31948 27300
rect 36306 27244 36316 27300
rect 36372 27244 37100 27300
rect 37156 27244 37166 27300
rect 39218 27244 39228 27300
rect 39284 27244 39676 27300
rect 39732 27244 40124 27300
rect 40180 27244 40190 27300
rect 53750 27244 53788 27300
rect 53844 27244 53854 27300
rect 56466 27244 56476 27300
rect 56532 27244 57036 27300
rect 57092 27244 57102 27300
rect 57362 27244 57372 27300
rect 57428 27244 57438 27300
rect 64866 27244 64876 27300
rect 64932 27244 65996 27300
rect 66052 27244 66062 27300
rect 71362 27244 71372 27300
rect 71428 27244 73052 27300
rect 73108 27244 73118 27300
rect 76402 27244 76412 27300
rect 76468 27244 77532 27300
rect 77588 27244 77598 27300
rect 20132 27188 20188 27244
rect 4498 27132 4508 27188
rect 4564 27132 5852 27188
rect 5908 27132 5918 27188
rect 9202 27132 9212 27188
rect 9268 27132 9548 27188
rect 9604 27132 16492 27188
rect 16548 27132 16558 27188
rect 16828 27132 17052 27188
rect 17108 27132 17118 27188
rect 20132 27132 23884 27188
rect 23940 27132 24780 27188
rect 24836 27132 24846 27188
rect 26684 27132 34468 27188
rect 34626 27132 34636 27188
rect 34692 27132 39900 27188
rect 39956 27132 39966 27188
rect 40786 27132 40796 27188
rect 40852 27132 41244 27188
rect 41300 27132 42140 27188
rect 42196 27132 44492 27188
rect 44548 27132 44558 27188
rect 44706 27132 44716 27188
rect 44772 27132 45500 27188
rect 45556 27132 45566 27188
rect 54338 27132 54348 27188
rect 54404 27132 55356 27188
rect 55412 27132 55422 27188
rect 3714 27020 3724 27076
rect 3780 27020 4396 27076
rect 4452 27020 5740 27076
rect 5796 27020 5806 27076
rect 6066 27020 6076 27076
rect 6132 27020 9996 27076
rect 10052 27020 10062 27076
rect 8306 26908 8316 26964
rect 8372 26908 8652 26964
rect 8708 26908 10668 26964
rect 10724 26908 10734 26964
rect 11666 26908 11676 26964
rect 11732 26908 12908 26964
rect 12964 26908 12974 26964
rect 13682 26908 13692 26964
rect 13748 26908 14364 26964
rect 14420 26908 15148 26964
rect 15204 26908 16156 26964
rect 16212 26908 16222 26964
rect 16828 26852 16884 27132
rect 17490 27020 17500 27076
rect 17556 27020 19068 27076
rect 19124 27020 22652 27076
rect 22708 27020 23212 27076
rect 23268 27020 24332 27076
rect 24388 27020 25228 27076
rect 25284 27020 26012 27076
rect 26068 27020 26078 27076
rect 26684 26964 26740 27132
rect 34412 27076 34468 27132
rect 57372 27076 57428 27244
rect 76178 27132 76188 27188
rect 76244 27132 78092 27188
rect 78148 27132 78158 27188
rect 31378 27020 31388 27076
rect 31444 27020 32060 27076
rect 32116 27020 32126 27076
rect 34412 27020 38556 27076
rect 38612 27020 39004 27076
rect 39060 27020 39788 27076
rect 39844 27020 39854 27076
rect 45042 27020 45052 27076
rect 45108 27020 46060 27076
rect 46116 27020 46126 27076
rect 46274 27020 46284 27076
rect 46340 27020 48524 27076
rect 48580 27020 48590 27076
rect 53554 27020 53564 27076
rect 53620 27020 53630 27076
rect 57372 27020 57708 27076
rect 57764 27020 57774 27076
rect 63074 27020 63084 27076
rect 63140 27020 63868 27076
rect 63924 27020 63934 27076
rect 67172 27020 68348 27076
rect 68404 27020 69468 27076
rect 69524 27020 69534 27076
rect 69794 27020 69804 27076
rect 69860 27020 70476 27076
rect 70532 27020 71036 27076
rect 71092 27020 71102 27076
rect 71922 27020 71932 27076
rect 71988 27020 72492 27076
rect 72548 27020 72558 27076
rect 76962 27020 76972 27076
rect 77028 27020 77308 27076
rect 77364 27020 77374 27076
rect 53564 26964 53620 27020
rect 67172 26964 67228 27020
rect 20066 26908 20076 26964
rect 20132 26908 20412 26964
rect 20468 26908 20748 26964
rect 20804 26908 21420 26964
rect 21476 26908 21486 26964
rect 22754 26908 22764 26964
rect 22820 26908 23548 26964
rect 23604 26908 24556 26964
rect 24612 26908 24622 26964
rect 24770 26908 24780 26964
rect 24836 26908 26124 26964
rect 26180 26908 26684 26964
rect 26740 26908 26750 26964
rect 28242 26908 28252 26964
rect 28308 26908 28812 26964
rect 28868 26908 28878 26964
rect 30930 26908 30940 26964
rect 30996 26908 31500 26964
rect 31556 26908 31566 26964
rect 31714 26908 31724 26964
rect 31780 26908 32396 26964
rect 32452 26908 32462 26964
rect 49298 26908 49308 26964
rect 49364 26908 54684 26964
rect 54740 26908 54750 26964
rect 59154 26908 59164 26964
rect 59220 26908 61292 26964
rect 61348 26908 61628 26964
rect 61684 26908 61694 26964
rect 63746 26908 63756 26964
rect 63812 26908 67228 26964
rect 72258 26908 72268 26964
rect 72324 26908 73836 26964
rect 73892 26908 75964 26964
rect 76020 26908 76030 26964
rect 77634 26908 77644 26964
rect 77700 26908 78988 26964
rect 79044 26908 79054 26964
rect 32396 26852 32452 26908
rect 7074 26796 7084 26852
rect 7140 26796 8204 26852
rect 8260 26796 8876 26852
rect 8932 26796 12796 26852
rect 12852 26796 12862 26852
rect 15092 26796 18172 26852
rect 18228 26796 18238 26852
rect 18834 26796 18844 26852
rect 18900 26796 19628 26852
rect 19684 26796 19694 26852
rect 19852 26796 20524 26852
rect 20580 26796 21532 26852
rect 21588 26796 22540 26852
rect 22596 26796 22606 26852
rect 26898 26796 26908 26852
rect 26964 26796 27916 26852
rect 27972 26796 28924 26852
rect 28980 26796 28990 26852
rect 32396 26796 36652 26852
rect 36708 26796 39676 26852
rect 39732 26796 39900 26852
rect 39956 26796 41692 26852
rect 41748 26796 41758 26852
rect 47394 26796 47404 26852
rect 47460 26796 52332 26852
rect 52388 26796 52398 26852
rect 55906 26796 55916 26852
rect 55972 26796 56700 26852
rect 56756 26796 57932 26852
rect 57988 26796 59500 26852
rect 59556 26796 59566 26852
rect 61954 26796 61964 26852
rect 62020 26796 63980 26852
rect 64036 26796 64046 26852
rect 68450 26796 68460 26852
rect 68516 26796 69916 26852
rect 69972 26796 69982 26852
rect 15092 26740 15148 26796
rect 19852 26740 19908 26796
rect 9538 26684 9548 26740
rect 9604 26684 11564 26740
rect 11620 26684 12012 26740
rect 12068 26684 15148 26740
rect 17042 26684 17052 26740
rect 17108 26684 18060 26740
rect 18116 26684 18956 26740
rect 19012 26684 19908 26740
rect 38658 26684 38668 26740
rect 38724 26684 39116 26740
rect 39172 26684 39182 26740
rect 43250 26684 43260 26740
rect 43316 26684 49196 26740
rect 49252 26684 49262 26740
rect 20522 26628 20532 26684
rect 20588 26628 20636 26684
rect 20692 26628 20740 26684
rect 20796 26628 20806 26684
rect 39842 26628 39852 26684
rect 39908 26628 39956 26684
rect 40012 26628 40060 26684
rect 40116 26628 40126 26684
rect 59162 26628 59172 26684
rect 59228 26628 59276 26684
rect 59332 26628 59380 26684
rect 59436 26628 59446 26684
rect 78482 26628 78492 26684
rect 78548 26628 78596 26684
rect 78652 26628 78700 26684
rect 78756 26628 78766 26684
rect 9986 26572 9996 26628
rect 10052 26572 13804 26628
rect 13860 26572 13870 26628
rect 26786 26572 26796 26628
rect 26852 26572 39564 26628
rect 39620 26572 39630 26628
rect 52770 26572 52780 26628
rect 52836 26572 53564 26628
rect 53620 26572 53630 26628
rect 53750 26572 53788 26628
rect 53844 26572 53854 26628
rect 73938 26572 73948 26628
rect 74004 26572 74172 26628
rect 74228 26572 74732 26628
rect 74788 26572 77308 26628
rect 77364 26572 77868 26628
rect 77924 26572 77934 26628
rect 12898 26460 12908 26516
rect 12964 26460 13580 26516
rect 13636 26460 13646 26516
rect 15250 26460 15260 26516
rect 15316 26460 15932 26516
rect 15988 26460 22988 26516
rect 23044 26460 25564 26516
rect 25620 26460 25630 26516
rect 27010 26460 27020 26516
rect 27076 26460 31948 26516
rect 34290 26460 34300 26516
rect 34356 26460 36540 26516
rect 36596 26460 36606 26516
rect 38612 26460 43148 26516
rect 43204 26460 43652 26516
rect 43922 26460 43932 26516
rect 43988 26460 45500 26516
rect 45556 26460 50428 26516
rect 52658 26460 52668 26516
rect 52724 26460 53452 26516
rect 53508 26460 53518 26516
rect 63298 26460 63308 26516
rect 63364 26460 65436 26516
rect 65492 26460 65502 26516
rect 74274 26460 74284 26516
rect 74340 26460 78316 26516
rect 78372 26460 78382 26516
rect 31892 26404 31948 26460
rect 38612 26404 38668 26460
rect 43596 26404 43652 26460
rect 50372 26404 50428 26460
rect 7410 26348 7420 26404
rect 7476 26348 7980 26404
rect 8036 26348 8876 26404
rect 8932 26348 8942 26404
rect 12002 26348 12012 26404
rect 12068 26348 12460 26404
rect 12516 26348 13356 26404
rect 13412 26348 13692 26404
rect 13748 26348 15148 26404
rect 15204 26348 15214 26404
rect 16146 26348 16156 26404
rect 16212 26348 16828 26404
rect 16884 26348 17500 26404
rect 17556 26348 17566 26404
rect 18162 26348 18172 26404
rect 18228 26348 18508 26404
rect 18564 26348 19852 26404
rect 19908 26348 20468 26404
rect 20626 26348 20636 26404
rect 20692 26348 21532 26404
rect 21588 26348 21598 26404
rect 21858 26348 21868 26404
rect 21924 26348 21934 26404
rect 31892 26348 38668 26404
rect 39890 26348 39900 26404
rect 39956 26348 41916 26404
rect 41972 26348 43372 26404
rect 43428 26348 43438 26404
rect 43596 26348 43820 26404
rect 43876 26348 44380 26404
rect 44436 26348 44446 26404
rect 48178 26348 48188 26404
rect 48244 26348 49756 26404
rect 49812 26348 49822 26404
rect 50372 26348 60060 26404
rect 60116 26348 61180 26404
rect 61236 26348 61246 26404
rect 20412 26292 20468 26348
rect 21868 26292 21924 26348
rect 3154 26236 3164 26292
rect 3220 26236 5292 26292
rect 5348 26236 7756 26292
rect 7812 26236 7822 26292
rect 10994 26236 11004 26292
rect 11060 26236 11676 26292
rect 11732 26236 11742 26292
rect 12460 26236 13916 26292
rect 13972 26236 16044 26292
rect 16100 26236 16110 26292
rect 17042 26236 17052 26292
rect 17108 26236 17948 26292
rect 18004 26236 18014 26292
rect 19506 26236 19516 26292
rect 19572 26236 20188 26292
rect 20244 26236 20254 26292
rect 20412 26236 21924 26292
rect 29810 26236 29820 26292
rect 29876 26236 30940 26292
rect 30996 26236 32284 26292
rect 32340 26236 32350 26292
rect 35634 26236 35644 26292
rect 35700 26236 36204 26292
rect 36260 26236 36270 26292
rect 38322 26236 38332 26292
rect 38388 26236 39788 26292
rect 39844 26236 39854 26292
rect 42018 26236 42028 26292
rect 42084 26236 44044 26292
rect 44100 26236 44492 26292
rect 44548 26236 44558 26292
rect 49186 26236 49196 26292
rect 49252 26236 50428 26292
rect 50484 26236 50494 26292
rect 50754 26236 50764 26292
rect 50820 26236 52668 26292
rect 52724 26236 52734 26292
rect 57698 26236 57708 26292
rect 57764 26236 59052 26292
rect 59108 26236 59118 26292
rect 62178 26236 62188 26292
rect 62244 26236 62860 26292
rect 62916 26236 62926 26292
rect 68002 26236 68012 26292
rect 68068 26236 69580 26292
rect 69636 26236 71260 26292
rect 71316 26236 71326 26292
rect 74162 26236 74172 26292
rect 74228 26236 75068 26292
rect 75124 26236 75628 26292
rect 75684 26236 75694 26292
rect 0 26180 800 26208
rect 12460 26180 12516 26236
rect 79200 26180 80000 26208
rect 0 26124 1932 26180
rect 1988 26124 1998 26180
rect 6850 26124 6860 26180
rect 6916 26124 7084 26180
rect 7140 26124 7308 26180
rect 7364 26124 7374 26180
rect 12450 26124 12460 26180
rect 12516 26124 12526 26180
rect 14130 26124 14140 26180
rect 14196 26124 14700 26180
rect 14756 26124 15260 26180
rect 15316 26124 15326 26180
rect 17154 26124 17164 26180
rect 17220 26124 18284 26180
rect 18340 26124 18350 26180
rect 22418 26124 22428 26180
rect 22484 26124 24108 26180
rect 24164 26124 24174 26180
rect 32386 26124 32396 26180
rect 32452 26124 35980 26180
rect 36036 26124 36046 26180
rect 39442 26124 39452 26180
rect 39508 26124 42140 26180
rect 42196 26124 42206 26180
rect 65202 26124 65212 26180
rect 65268 26124 65996 26180
rect 66052 26124 66062 26180
rect 75506 26124 75516 26180
rect 75572 26124 80000 26180
rect 0 26096 800 26124
rect 79200 26096 80000 26124
rect 8866 26012 8876 26068
rect 8932 26012 9660 26068
rect 9716 26012 11284 26068
rect 29810 26012 29820 26068
rect 29876 26012 30492 26068
rect 30548 26012 32508 26068
rect 32564 26012 32574 26068
rect 34290 26012 34300 26068
rect 34356 26012 38332 26068
rect 38388 26012 38398 26068
rect 48402 26012 48412 26068
rect 48468 26012 49532 26068
rect 49588 26012 49598 26068
rect 67106 26012 67116 26068
rect 67172 26012 67676 26068
rect 67732 26012 67742 26068
rect 72034 26012 72044 26068
rect 72100 26012 74284 26068
rect 74340 26012 74350 26068
rect 11228 25956 11284 26012
rect 3602 25900 3612 25956
rect 3668 25900 4620 25956
rect 4676 25900 7644 25956
rect 7700 25900 7710 25956
rect 11228 25900 14588 25956
rect 14644 25900 14812 25956
rect 14868 25900 15708 25956
rect 15764 25900 25676 25956
rect 25732 25900 25742 25956
rect 26898 25900 26908 25956
rect 26964 25900 27356 25956
rect 27412 25900 27692 25956
rect 27748 25900 27758 25956
rect 74386 25900 74396 25956
rect 74452 25900 75852 25956
rect 75908 25900 77756 25956
rect 77812 25900 77822 25956
rect 10862 25844 10872 25900
rect 10928 25844 10976 25900
rect 11032 25844 11080 25900
rect 11136 25844 11146 25900
rect 30182 25844 30192 25900
rect 30248 25844 30296 25900
rect 30352 25844 30400 25900
rect 30456 25844 30466 25900
rect 49502 25844 49512 25900
rect 49568 25844 49616 25900
rect 49672 25844 49720 25900
rect 49776 25844 49786 25900
rect 68822 25844 68832 25900
rect 68888 25844 68936 25900
rect 68992 25844 69040 25900
rect 69096 25844 69106 25900
rect 20514 25788 20524 25844
rect 20580 25788 21756 25844
rect 21812 25788 21822 25844
rect 38658 25788 38668 25844
rect 38724 25788 39564 25844
rect 39620 25788 40348 25844
rect 40404 25788 40414 25844
rect 50372 25788 68124 25844
rect 68180 25788 68190 25844
rect 1362 25676 1372 25732
rect 1428 25676 47404 25732
rect 47460 25676 47470 25732
rect 50372 25620 50428 25788
rect 56354 25676 56364 25732
rect 56420 25676 57148 25732
rect 57204 25676 57708 25732
rect 57764 25676 57774 25732
rect 60722 25676 60732 25732
rect 60788 25676 62860 25732
rect 62916 25676 64652 25732
rect 64708 25676 64718 25732
rect 74946 25676 74956 25732
rect 75012 25676 77308 25732
rect 77364 25676 77374 25732
rect 3266 25564 3276 25620
rect 3332 25564 3612 25620
rect 3668 25564 5516 25620
rect 5572 25564 5582 25620
rect 7410 25564 7420 25620
rect 7476 25564 7486 25620
rect 15138 25564 15148 25620
rect 15204 25564 16156 25620
rect 16212 25564 16222 25620
rect 19282 25564 19292 25620
rect 19348 25564 20300 25620
rect 20356 25564 20636 25620
rect 20692 25564 20702 25620
rect 25666 25564 25676 25620
rect 25732 25564 26796 25620
rect 26852 25564 26862 25620
rect 28018 25564 28028 25620
rect 28084 25564 29708 25620
rect 29764 25564 29774 25620
rect 31892 25564 50428 25620
rect 58370 25564 58380 25620
rect 58436 25564 61516 25620
rect 61572 25564 61582 25620
rect 62412 25564 64204 25620
rect 64260 25564 65212 25620
rect 65268 25564 66388 25620
rect 66770 25564 66780 25620
rect 66836 25564 67788 25620
rect 67844 25564 67854 25620
rect 76514 25564 76524 25620
rect 76580 25564 77420 25620
rect 77476 25564 77486 25620
rect 7420 25172 7476 25564
rect 31892 25508 31948 25564
rect 62412 25508 62468 25564
rect 12114 25452 12124 25508
rect 12180 25452 12190 25508
rect 18386 25452 18396 25508
rect 18452 25452 21980 25508
rect 22036 25452 22046 25508
rect 24882 25452 24892 25508
rect 24948 25452 27412 25508
rect 27570 25452 27580 25508
rect 27636 25452 27916 25508
rect 27972 25452 27982 25508
rect 28140 25452 31948 25508
rect 33058 25452 33068 25508
rect 33124 25452 34300 25508
rect 34356 25452 34366 25508
rect 39106 25452 39116 25508
rect 39172 25452 39340 25508
rect 39396 25452 39900 25508
rect 39956 25452 39966 25508
rect 40114 25452 40124 25508
rect 40180 25452 40796 25508
rect 40852 25452 40862 25508
rect 44370 25452 44380 25508
rect 44436 25452 44940 25508
rect 44996 25452 45006 25508
rect 53330 25452 53340 25508
rect 53396 25452 53900 25508
rect 53956 25452 53966 25508
rect 57138 25452 57148 25508
rect 57204 25452 58604 25508
rect 58660 25452 59052 25508
rect 59108 25452 59948 25508
rect 60004 25452 60014 25508
rect 61282 25452 61292 25508
rect 61348 25452 62412 25508
rect 62468 25452 62478 25508
rect 62626 25452 62636 25508
rect 62692 25452 63308 25508
rect 63364 25452 63374 25508
rect 12124 25396 12180 25452
rect 27356 25396 27412 25452
rect 28140 25396 28196 25452
rect 66332 25396 66388 25564
rect 12124 25340 20132 25396
rect 21858 25340 21868 25396
rect 21924 25340 25228 25396
rect 25284 25340 25294 25396
rect 26226 25340 26236 25396
rect 26292 25340 26684 25396
rect 26740 25340 27132 25396
rect 27188 25340 27198 25396
rect 27356 25340 28196 25396
rect 30930 25340 30940 25396
rect 30996 25340 33180 25396
rect 33236 25340 33852 25396
rect 33908 25340 33918 25396
rect 39666 25340 39676 25396
rect 39732 25340 41244 25396
rect 41300 25340 41310 25396
rect 44594 25340 44604 25396
rect 44660 25340 45500 25396
rect 45556 25340 45566 25396
rect 56466 25340 56476 25396
rect 56532 25340 57036 25396
rect 57092 25340 57484 25396
rect 57540 25340 58940 25396
rect 58996 25340 60396 25396
rect 60452 25340 60462 25396
rect 62178 25340 62188 25396
rect 62244 25340 63868 25396
rect 63924 25340 65436 25396
rect 65492 25340 65502 25396
rect 66322 25340 66332 25396
rect 66388 25340 66398 25396
rect 66994 25340 67004 25396
rect 67060 25340 67676 25396
rect 67732 25340 67742 25396
rect 68562 25340 68572 25396
rect 68628 25340 69916 25396
rect 69972 25340 70588 25396
rect 70644 25340 70654 25396
rect 20076 25284 20132 25340
rect 9874 25228 9884 25284
rect 9940 25228 15932 25284
rect 15988 25228 15998 25284
rect 20066 25228 20076 25284
rect 20132 25228 20142 25284
rect 20514 25228 20524 25284
rect 20580 25228 20860 25284
rect 20916 25228 22092 25284
rect 22148 25228 22428 25284
rect 22484 25228 22652 25284
rect 22708 25228 23548 25284
rect 23604 25228 23614 25284
rect 39218 25228 39228 25284
rect 39284 25228 41468 25284
rect 41524 25228 41534 25284
rect 42018 25228 42028 25284
rect 42084 25228 45612 25284
rect 45668 25228 45678 25284
rect 59154 25228 59164 25284
rect 59220 25228 60564 25284
rect 60834 25228 60844 25284
rect 60900 25228 63084 25284
rect 63140 25228 63150 25284
rect 66658 25228 66668 25284
rect 66724 25228 67900 25284
rect 67956 25228 67966 25284
rect 60508 25172 60564 25228
rect 5282 25116 5292 25172
rect 5348 25116 7476 25172
rect 9986 25116 9996 25172
rect 10052 25116 11900 25172
rect 11956 25116 12572 25172
rect 12628 25116 12908 25172
rect 12964 25116 12974 25172
rect 60508 25116 63980 25172
rect 64036 25116 64046 25172
rect 74834 25116 74844 25172
rect 74900 25116 75852 25172
rect 75908 25116 75918 25172
rect 20522 25060 20532 25116
rect 20588 25060 20636 25116
rect 20692 25060 20740 25116
rect 20796 25060 20806 25116
rect 39842 25060 39852 25116
rect 39908 25060 39956 25116
rect 40012 25060 40060 25116
rect 40116 25060 40126 25116
rect 59162 25060 59172 25116
rect 59228 25060 59276 25116
rect 59332 25060 59380 25116
rect 59436 25060 59446 25116
rect 78482 25060 78492 25116
rect 78548 25060 78596 25116
rect 78652 25060 78700 25116
rect 78756 25060 78766 25116
rect 10770 25004 10780 25060
rect 10836 25004 12124 25060
rect 12180 25004 13300 25060
rect 22306 25004 22316 25060
rect 22372 25004 23100 25060
rect 23156 25004 23166 25060
rect 13244 24948 13300 25004
rect 4386 24892 4396 24948
rect 4452 24892 12460 24948
rect 12516 24892 12526 24948
rect 13234 24892 13244 24948
rect 13300 24892 21868 24948
rect 21924 24892 49308 24948
rect 49364 24892 49374 24948
rect 58482 24892 58492 24948
rect 58548 24892 59052 24948
rect 59108 24892 59118 24948
rect 63410 24892 63420 24948
rect 63476 24892 64540 24948
rect 64596 24892 64606 24948
rect 64754 24892 64764 24948
rect 64820 24892 65996 24948
rect 66052 24892 66780 24948
rect 66836 24892 66846 24948
rect 12002 24780 12012 24836
rect 12068 24780 16268 24836
rect 16324 24780 23324 24836
rect 23380 24780 24444 24836
rect 24500 24780 24510 24836
rect 24882 24780 24892 24836
rect 24948 24780 26124 24836
rect 26180 24780 26190 24836
rect 30594 24780 30604 24836
rect 30660 24780 32732 24836
rect 32788 24780 32798 24836
rect 33852 24780 35420 24836
rect 35476 24780 35486 24836
rect 43474 24780 43484 24836
rect 43540 24780 44044 24836
rect 44100 24780 44110 24836
rect 59266 24780 59276 24836
rect 59332 24780 60060 24836
rect 60116 24780 60126 24836
rect 62402 24780 62412 24836
rect 62468 24780 69020 24836
rect 69076 24780 69804 24836
rect 69860 24780 70700 24836
rect 70756 24780 70766 24836
rect 75842 24780 75852 24836
rect 75908 24780 76692 24836
rect 76850 24780 76860 24836
rect 76916 24780 77644 24836
rect 77700 24780 77710 24836
rect 33852 24724 33908 24780
rect 76636 24724 76692 24780
rect 7074 24668 7084 24724
rect 7140 24668 9660 24724
rect 9716 24668 9726 24724
rect 11218 24668 11228 24724
rect 11284 24668 13020 24724
rect 13076 24668 13086 24724
rect 13682 24668 13692 24724
rect 13748 24668 14364 24724
rect 14420 24668 15820 24724
rect 15876 24668 15886 24724
rect 25666 24668 25676 24724
rect 25732 24668 26348 24724
rect 26404 24668 26414 24724
rect 30482 24668 30492 24724
rect 30548 24668 30716 24724
rect 30772 24668 30782 24724
rect 32498 24668 32508 24724
rect 32564 24668 33852 24724
rect 33908 24668 33918 24724
rect 34066 24668 34076 24724
rect 34132 24668 34524 24724
rect 34580 24668 35308 24724
rect 35364 24668 35374 24724
rect 64978 24668 64988 24724
rect 65044 24668 65436 24724
rect 65492 24668 67788 24724
rect 67844 24668 67854 24724
rect 75282 24668 75292 24724
rect 75348 24668 76412 24724
rect 76468 24668 76478 24724
rect 76636 24668 77532 24724
rect 77588 24668 77598 24724
rect 7420 24388 7476 24668
rect 11554 24556 11564 24612
rect 11620 24556 12012 24612
rect 12068 24556 12078 24612
rect 14914 24556 14924 24612
rect 14980 24556 16044 24612
rect 16100 24556 16110 24612
rect 22978 24556 22988 24612
rect 23044 24556 23212 24612
rect 23268 24556 23996 24612
rect 24052 24556 24062 24612
rect 25554 24556 25564 24612
rect 25620 24556 26572 24612
rect 26628 24556 26638 24612
rect 32834 24556 32844 24612
rect 32900 24556 33628 24612
rect 33684 24556 33694 24612
rect 34626 24556 34636 24612
rect 34692 24556 37100 24612
rect 37156 24556 37996 24612
rect 38052 24556 38062 24612
rect 44258 24556 44268 24612
rect 44324 24556 45388 24612
rect 45444 24556 60844 24612
rect 60900 24556 60910 24612
rect 66770 24556 66780 24612
rect 66836 24556 67228 24612
rect 67284 24556 67294 24612
rect 73490 24556 73500 24612
rect 73556 24556 74060 24612
rect 74116 24556 74126 24612
rect 75170 24556 75180 24612
rect 75236 24556 76300 24612
rect 76356 24556 77420 24612
rect 77476 24556 77486 24612
rect 15922 24444 15932 24500
rect 15988 24444 31052 24500
rect 31108 24444 31118 24500
rect 7410 24332 7420 24388
rect 7476 24332 7486 24388
rect 10862 24276 10872 24332
rect 10928 24276 10976 24332
rect 11032 24276 11080 24332
rect 11136 24276 11146 24332
rect 30182 24276 30192 24332
rect 30248 24276 30296 24332
rect 30352 24276 30400 24332
rect 30456 24276 30466 24332
rect 49502 24276 49512 24332
rect 49568 24276 49616 24332
rect 49672 24276 49720 24332
rect 49776 24276 49786 24332
rect 68822 24276 68832 24332
rect 68888 24276 68936 24332
rect 68992 24276 69040 24332
rect 69096 24276 69106 24332
rect 12226 24220 12236 24276
rect 12292 24220 15148 24276
rect 15204 24220 15214 24276
rect 17602 24220 17612 24276
rect 17668 24220 19852 24276
rect 19908 24220 19918 24276
rect 35746 24220 35756 24276
rect 35812 24220 42364 24276
rect 42420 24220 42430 24276
rect 7634 24108 7644 24164
rect 7700 24108 8092 24164
rect 8148 24108 10108 24164
rect 10164 24108 10174 24164
rect 10780 24108 22988 24164
rect 23044 24108 23054 24164
rect 24434 24108 24444 24164
rect 24500 24108 48748 24164
rect 48804 24108 49756 24164
rect 49812 24108 50316 24164
rect 50372 24108 50382 24164
rect 10780 23940 10836 24108
rect 11778 23996 11788 24052
rect 11844 23996 12124 24052
rect 12180 23996 12190 24052
rect 19506 23996 19516 24052
rect 19572 23996 22876 24052
rect 22932 23996 22942 24052
rect 26002 23996 26012 24052
rect 26068 23996 27244 24052
rect 27300 23996 27310 24052
rect 28242 23996 28252 24052
rect 28308 23996 37828 24052
rect 38098 23996 38108 24052
rect 38164 23996 38892 24052
rect 38948 23996 38958 24052
rect 49298 23996 49308 24052
rect 49364 23996 49868 24052
rect 49924 23996 49934 24052
rect 65538 23996 65548 24052
rect 65604 23996 67116 24052
rect 67172 23996 67340 24052
rect 67396 23996 67406 24052
rect 11788 23940 11844 23996
rect 37772 23940 37828 23996
rect 7858 23884 7868 23940
rect 7924 23884 8428 23940
rect 8484 23884 10836 23940
rect 10994 23884 11004 23940
rect 11060 23884 11228 23940
rect 11284 23884 11844 23940
rect 12898 23884 12908 23940
rect 12964 23884 14028 23940
rect 14084 23884 14094 23940
rect 18610 23884 18620 23940
rect 18676 23884 19292 23940
rect 19348 23884 19358 23940
rect 21858 23884 21868 23940
rect 21924 23884 23100 23940
rect 23156 23884 23166 23940
rect 33954 23884 33964 23940
rect 34020 23884 34636 23940
rect 34692 23884 34702 23940
rect 37772 23884 56812 23940
rect 56868 23884 57596 23940
rect 57652 23884 57662 23940
rect 58370 23884 58380 23940
rect 58436 23884 61740 23940
rect 61796 23884 61806 23940
rect 62066 23884 62076 23940
rect 62132 23884 69244 23940
rect 69300 23884 69310 23940
rect 76178 23884 76188 23940
rect 76244 23884 77308 23940
rect 77364 23884 77374 23940
rect 57596 23828 57652 23884
rect 3154 23772 3164 23828
rect 3220 23772 3612 23828
rect 3668 23772 3678 23828
rect 10546 23772 10556 23828
rect 10612 23772 11340 23828
rect 11396 23772 11406 23828
rect 11666 23772 11676 23828
rect 11732 23772 24892 23828
rect 24948 23772 25452 23828
rect 25508 23772 25518 23828
rect 25666 23772 25676 23828
rect 25732 23772 27916 23828
rect 27972 23772 28252 23828
rect 28308 23772 28318 23828
rect 29698 23772 29708 23828
rect 29764 23772 30044 23828
rect 30100 23772 30268 23828
rect 30324 23772 30334 23828
rect 41122 23772 41132 23828
rect 41188 23772 42700 23828
rect 42756 23772 42766 23828
rect 46946 23772 46956 23828
rect 47012 23772 47516 23828
rect 47572 23772 47582 23828
rect 57596 23772 59052 23828
rect 59108 23772 59118 23828
rect 59714 23772 59724 23828
rect 59780 23772 60396 23828
rect 60452 23772 60732 23828
rect 60788 23772 60798 23828
rect 66322 23772 66332 23828
rect 66388 23772 67900 23828
rect 67956 23772 67966 23828
rect 0 23716 800 23744
rect 79200 23716 80000 23744
rect 0 23660 1932 23716
rect 1988 23660 1998 23716
rect 2930 23660 2940 23716
rect 2996 23660 3836 23716
rect 3892 23660 3902 23716
rect 9202 23660 9212 23716
rect 9268 23660 9996 23716
rect 10052 23660 10062 23716
rect 21858 23660 21868 23716
rect 21924 23660 22316 23716
rect 22372 23660 22988 23716
rect 23044 23660 23054 23716
rect 23538 23660 23548 23716
rect 23604 23660 24444 23716
rect 24500 23660 25900 23716
rect 25956 23660 25966 23716
rect 26898 23660 26908 23716
rect 26964 23660 30380 23716
rect 30436 23660 30716 23716
rect 30772 23660 30782 23716
rect 32610 23660 32620 23716
rect 32676 23660 33628 23716
rect 33684 23660 34748 23716
rect 34804 23660 34814 23716
rect 34962 23660 34972 23716
rect 35028 23660 35532 23716
rect 35588 23660 35598 23716
rect 36866 23660 36876 23716
rect 36932 23660 37772 23716
rect 37828 23660 37838 23716
rect 41682 23660 41692 23716
rect 41748 23660 42140 23716
rect 42196 23660 42206 23716
rect 49970 23660 49980 23716
rect 50036 23660 52556 23716
rect 52612 23660 53788 23716
rect 53844 23660 54348 23716
rect 54404 23660 54414 23716
rect 58258 23660 58268 23716
rect 58324 23660 59276 23716
rect 59332 23660 59342 23716
rect 59826 23660 59836 23716
rect 59892 23660 60284 23716
rect 60340 23660 60844 23716
rect 60900 23660 60910 23716
rect 66434 23660 66444 23716
rect 66500 23660 67452 23716
rect 67508 23660 67518 23716
rect 75506 23660 75516 23716
rect 75572 23660 80000 23716
rect 0 23632 800 23660
rect 8754 23548 8764 23604
rect 8820 23548 9660 23604
rect 9716 23548 11116 23604
rect 11172 23548 18060 23604
rect 18116 23548 18126 23604
rect 60050 23548 60060 23604
rect 60116 23548 61852 23604
rect 61908 23548 61918 23604
rect 64082 23548 64092 23604
rect 64148 23548 64988 23604
rect 65044 23548 65324 23604
rect 65380 23548 65390 23604
rect 20522 23492 20532 23548
rect 20588 23492 20636 23548
rect 20692 23492 20740 23548
rect 20796 23492 20806 23548
rect 39842 23492 39852 23548
rect 39908 23492 39956 23548
rect 40012 23492 40060 23548
rect 40116 23492 40126 23548
rect 59162 23492 59172 23548
rect 59228 23492 59276 23548
rect 59332 23492 59380 23548
rect 59436 23492 59446 23548
rect 66444 23492 66500 23660
rect 79200 23632 80000 23660
rect 78482 23492 78492 23548
rect 78548 23492 78596 23548
rect 78652 23492 78700 23548
rect 78756 23492 78766 23548
rect 4386 23436 4396 23492
rect 4452 23436 4732 23492
rect 4788 23436 5628 23492
rect 5684 23436 5694 23492
rect 17266 23436 17276 23492
rect 17332 23436 18284 23492
rect 18340 23436 18350 23492
rect 19170 23436 19180 23492
rect 19236 23436 20188 23492
rect 20244 23436 20254 23492
rect 26562 23436 26572 23492
rect 26628 23436 27356 23492
rect 27412 23436 27422 23492
rect 50082 23436 50092 23492
rect 50148 23436 50988 23492
rect 51044 23436 56140 23492
rect 56196 23436 56700 23492
rect 56756 23436 56766 23492
rect 64866 23436 64876 23492
rect 64932 23436 66500 23492
rect 72594 23436 72604 23492
rect 72660 23436 73612 23492
rect 73668 23436 75628 23492
rect 75684 23436 75694 23492
rect 5842 23324 5852 23380
rect 5908 23324 29596 23380
rect 29652 23324 29662 23380
rect 42242 23324 42252 23380
rect 42308 23324 50428 23380
rect 52546 23324 52556 23380
rect 52612 23324 53452 23380
rect 53508 23324 53518 23380
rect 60050 23324 60060 23380
rect 60116 23324 60620 23380
rect 60676 23324 61292 23380
rect 61348 23324 61358 23380
rect 72146 23324 72156 23380
rect 72212 23324 73500 23380
rect 73556 23324 73566 23380
rect 50372 23268 50428 23324
rect 18050 23212 18060 23268
rect 18116 23212 19068 23268
rect 19124 23212 19134 23268
rect 19954 23212 19964 23268
rect 20020 23212 21196 23268
rect 21252 23212 21644 23268
rect 21700 23212 21710 23268
rect 25218 23212 25228 23268
rect 25284 23212 25900 23268
rect 25956 23212 26572 23268
rect 26628 23212 37212 23268
rect 37268 23212 37278 23268
rect 46162 23212 46172 23268
rect 46228 23212 47180 23268
rect 47236 23212 47740 23268
rect 47796 23212 47806 23268
rect 50372 23212 78316 23268
rect 78372 23212 78382 23268
rect 6962 23100 6972 23156
rect 7028 23100 8204 23156
rect 8260 23100 9940 23156
rect 10098 23100 10108 23156
rect 10164 23100 13468 23156
rect 13524 23100 13916 23156
rect 13972 23100 13982 23156
rect 9884 23044 9940 23100
rect 19068 23044 19124 23212
rect 19394 23100 19404 23156
rect 19460 23100 20636 23156
rect 20692 23100 21308 23156
rect 21364 23100 21374 23156
rect 34066 23100 34076 23156
rect 34132 23100 38668 23156
rect 38724 23100 38734 23156
rect 39554 23100 39564 23156
rect 39620 23100 40236 23156
rect 40292 23100 40302 23156
rect 40898 23100 40908 23156
rect 40964 23100 41916 23156
rect 41972 23100 41982 23156
rect 44258 23100 44268 23156
rect 44324 23100 45500 23156
rect 45556 23100 45566 23156
rect 52434 23100 52444 23156
rect 52500 23100 53676 23156
rect 53732 23100 53742 23156
rect 55570 23100 55580 23156
rect 55636 23100 56700 23156
rect 56756 23100 57484 23156
rect 57540 23100 58156 23156
rect 58212 23100 58222 23156
rect 60022 23100 60060 23156
rect 60116 23100 60126 23156
rect 60284 23100 62748 23156
rect 62804 23100 62814 23156
rect 66098 23100 66108 23156
rect 66164 23100 68572 23156
rect 68628 23100 68638 23156
rect 72146 23100 72156 23156
rect 72212 23100 73612 23156
rect 73668 23100 73678 23156
rect 60284 23044 60340 23100
rect 3378 22988 3388 23044
rect 3444 22988 5068 23044
rect 5124 22988 5134 23044
rect 6402 22988 6412 23044
rect 6468 22988 7084 23044
rect 7140 22988 7756 23044
rect 7812 22988 9828 23044
rect 9884 22988 18284 23044
rect 18340 22988 18350 23044
rect 19068 22988 23548 23044
rect 23604 22988 24108 23044
rect 24164 22988 24174 23044
rect 36194 22988 36204 23044
rect 36260 22988 36764 23044
rect 36820 22988 36830 23044
rect 44482 22988 44492 23044
rect 44548 22988 45612 23044
rect 45668 22988 45678 23044
rect 47842 22988 47852 23044
rect 47908 22988 48636 23044
rect 48692 22988 48702 23044
rect 58930 22988 58940 23044
rect 58996 22988 59500 23044
rect 59556 22988 60340 23044
rect 65986 22988 65996 23044
rect 66052 22988 70588 23044
rect 70644 22988 71260 23044
rect 71316 22988 71326 23044
rect 73266 22988 73276 23044
rect 73332 22988 75740 23044
rect 75796 22988 76860 23044
rect 76916 22988 76926 23044
rect 9772 22932 9828 22988
rect 4610 22876 4620 22932
rect 4676 22876 9324 22932
rect 9380 22876 9390 22932
rect 9772 22876 17836 22932
rect 17892 22876 17902 22932
rect 18498 22876 18508 22932
rect 18564 22876 19180 22932
rect 19236 22876 19246 22932
rect 47282 22876 47292 22932
rect 47348 22876 48076 22932
rect 48132 22876 48142 22932
rect 57586 22876 57596 22932
rect 57652 22876 58044 22932
rect 58100 22876 59948 22932
rect 60004 22876 60014 22932
rect 12674 22764 12684 22820
rect 12740 22764 21028 22820
rect 10862 22708 10872 22764
rect 10928 22708 10976 22764
rect 11032 22708 11080 22764
rect 11136 22708 11146 22764
rect 8978 22652 8988 22708
rect 9044 22652 9772 22708
rect 9828 22652 9838 22708
rect 13346 22652 13356 22708
rect 13412 22652 16212 22708
rect 2482 22540 2492 22596
rect 2548 22540 2828 22596
rect 2884 22540 4508 22596
rect 4564 22540 11676 22596
rect 11732 22540 11742 22596
rect 12114 22540 12124 22596
rect 12180 22540 12572 22596
rect 12628 22540 14812 22596
rect 14868 22540 14878 22596
rect 16156 22484 16212 22652
rect 20972 22596 21028 22764
rect 30182 22708 30192 22764
rect 30248 22708 30296 22764
rect 30352 22708 30400 22764
rect 30456 22708 30466 22764
rect 49502 22708 49512 22764
rect 49568 22708 49616 22764
rect 49672 22708 49720 22764
rect 49776 22708 49786 22764
rect 68822 22708 68832 22764
rect 68888 22708 68936 22764
rect 68992 22708 69040 22764
rect 69096 22708 69106 22764
rect 26674 22652 26684 22708
rect 26740 22652 27916 22708
rect 27972 22652 29148 22708
rect 29204 22652 29214 22708
rect 30706 22652 30716 22708
rect 30772 22652 38668 22708
rect 40562 22652 40572 22708
rect 40628 22652 41580 22708
rect 41636 22652 41646 22708
rect 50978 22652 50988 22708
rect 51044 22652 55916 22708
rect 55972 22652 56476 22708
rect 56532 22652 56542 22708
rect 71148 22652 71372 22708
rect 71428 22652 71438 22708
rect 38612 22596 38668 22652
rect 71148 22596 71204 22652
rect 20972 22540 33740 22596
rect 33796 22540 33806 22596
rect 38612 22540 47404 22596
rect 47460 22540 47470 22596
rect 49522 22540 49532 22596
rect 49588 22540 52220 22596
rect 52276 22540 53900 22596
rect 53956 22540 53966 22596
rect 63522 22540 63532 22596
rect 63588 22540 71148 22596
rect 71204 22540 71214 22596
rect 71474 22540 71484 22596
rect 71540 22540 73948 22596
rect 74004 22540 74014 22596
rect 3042 22428 3052 22484
rect 3108 22428 3388 22484
rect 3444 22428 3454 22484
rect 6178 22428 6188 22484
rect 6244 22428 6748 22484
rect 6804 22428 6814 22484
rect 8530 22428 8540 22484
rect 8596 22428 9436 22484
rect 9492 22428 9772 22484
rect 9828 22428 9838 22484
rect 13794 22428 13804 22484
rect 13860 22428 15148 22484
rect 16156 22428 51436 22484
rect 51492 22428 51502 22484
rect 58370 22428 58380 22484
rect 58436 22428 59164 22484
rect 59220 22428 59836 22484
rect 59892 22428 60620 22484
rect 60676 22428 60686 22484
rect 69234 22428 69244 22484
rect 69300 22428 72492 22484
rect 72548 22428 73388 22484
rect 73444 22428 73454 22484
rect 15092 22372 15148 22428
rect 12898 22316 12908 22372
rect 12964 22316 13692 22372
rect 13748 22316 13758 22372
rect 15092 22316 21084 22372
rect 21140 22316 21150 22372
rect 32946 22316 32956 22372
rect 33012 22316 34076 22372
rect 34132 22316 34142 22372
rect 40338 22316 40348 22372
rect 40404 22316 40908 22372
rect 40964 22316 40974 22372
rect 42466 22316 42476 22372
rect 42532 22316 45724 22372
rect 45780 22316 45790 22372
rect 48066 22316 48076 22372
rect 48132 22316 49420 22372
rect 49476 22316 49486 22372
rect 57484 22316 60396 22372
rect 60452 22316 60462 22372
rect 65090 22316 65100 22372
rect 65156 22316 66668 22372
rect 66724 22316 67116 22372
rect 67172 22316 67182 22372
rect 72930 22316 72940 22372
rect 72996 22316 75628 22372
rect 75684 22316 76748 22372
rect 76804 22316 76814 22372
rect 45724 22260 45780 22316
rect 57484 22260 57540 22316
rect 8082 22204 8092 22260
rect 8148 22204 9436 22260
rect 9492 22204 9996 22260
rect 10052 22204 10062 22260
rect 12786 22204 12796 22260
rect 12852 22204 14924 22260
rect 14980 22204 14990 22260
rect 16482 22204 16492 22260
rect 16548 22204 20076 22260
rect 20132 22204 20142 22260
rect 24770 22204 24780 22260
rect 24836 22204 25228 22260
rect 25284 22204 26348 22260
rect 26404 22204 26796 22260
rect 26852 22204 26862 22260
rect 43026 22204 43036 22260
rect 43092 22204 43820 22260
rect 43876 22204 44828 22260
rect 44884 22204 44894 22260
rect 45724 22204 48188 22260
rect 48244 22204 48254 22260
rect 51762 22204 51772 22260
rect 51828 22204 53452 22260
rect 53508 22204 53518 22260
rect 57474 22204 57484 22260
rect 57540 22204 57550 22260
rect 58594 22204 58604 22260
rect 58660 22204 59948 22260
rect 60004 22204 60014 22260
rect 63746 22204 63756 22260
rect 63812 22204 64876 22260
rect 64932 22204 65324 22260
rect 65380 22204 65390 22260
rect 65538 22204 65548 22260
rect 65604 22204 66108 22260
rect 66164 22204 68348 22260
rect 68404 22204 68414 22260
rect 74386 22204 74396 22260
rect 74452 22204 75404 22260
rect 75460 22204 77532 22260
rect 77588 22204 77598 22260
rect 13916 22148 13972 22204
rect 13906 22092 13916 22148
rect 13972 22092 13982 22148
rect 27122 22092 27132 22148
rect 27188 22092 27692 22148
rect 27748 22092 28140 22148
rect 28196 22092 30604 22148
rect 30660 22092 30670 22148
rect 36754 22092 36764 22148
rect 36820 22092 36988 22148
rect 37044 22092 37660 22148
rect 37716 22092 37996 22148
rect 38052 22092 38444 22148
rect 38500 22092 38510 22148
rect 38612 22092 45388 22148
rect 45444 22092 45948 22148
rect 46004 22092 47292 22148
rect 47348 22092 47852 22148
rect 47908 22092 47918 22148
rect 49970 22092 49980 22148
rect 50036 22092 52444 22148
rect 52500 22092 52510 22148
rect 55458 22092 55468 22148
rect 55524 22092 56476 22148
rect 56532 22092 58268 22148
rect 58324 22092 58334 22148
rect 58706 22092 58716 22148
rect 58772 22092 59388 22148
rect 59444 22092 59724 22148
rect 59780 22092 61348 22148
rect 65650 22092 65660 22148
rect 65716 22092 66444 22148
rect 66500 22092 67900 22148
rect 67956 22092 67966 22148
rect 71026 22092 71036 22148
rect 71092 22092 74732 22148
rect 74788 22092 74798 22148
rect 77074 22092 77084 22148
rect 77140 22092 77756 22148
rect 77812 22092 77822 22148
rect 38612 22036 38668 22092
rect 61292 22036 61348 22092
rect 27570 21980 27580 22036
rect 27636 21980 28588 22036
rect 28644 21980 36204 22036
rect 36260 21980 36270 22036
rect 36642 21980 36652 22036
rect 36708 21980 38668 22036
rect 52108 21980 58380 22036
rect 58436 21980 58446 22036
rect 61282 21980 61292 22036
rect 61348 21980 65660 22036
rect 65716 21980 65726 22036
rect 67218 21980 67228 22036
rect 67284 21980 73276 22036
rect 73332 21980 73342 22036
rect 20522 21924 20532 21980
rect 20588 21924 20636 21980
rect 20692 21924 20740 21980
rect 20796 21924 20806 21980
rect 39842 21924 39852 21980
rect 39908 21924 39956 21980
rect 40012 21924 40060 21980
rect 40116 21924 40126 21980
rect 9314 21868 9324 21924
rect 9380 21868 9940 21924
rect 24434 21868 24444 21924
rect 24500 21868 25676 21924
rect 25732 21868 26460 21924
rect 26516 21868 26526 21924
rect 50194 21868 50204 21924
rect 50260 21868 51884 21924
rect 51940 21868 51950 21924
rect 9884 21812 9940 21868
rect 52108 21812 52164 21980
rect 59162 21924 59172 21980
rect 59228 21924 59276 21980
rect 59332 21924 59380 21980
rect 59436 21924 59446 21980
rect 78482 21924 78492 21980
rect 78548 21924 78596 21980
rect 78652 21924 78700 21980
rect 78756 21924 78766 21980
rect 52434 21868 52444 21924
rect 52500 21868 57596 21924
rect 57652 21868 57988 21924
rect 58146 21868 58156 21924
rect 58212 21868 58996 21924
rect 65762 21868 65772 21924
rect 65828 21868 67452 21924
rect 67508 21868 67518 21924
rect 57932 21812 57988 21868
rect 58940 21812 58996 21868
rect 2034 21756 2044 21812
rect 2100 21756 2716 21812
rect 2772 21756 5292 21812
rect 5348 21756 5358 21812
rect 5506 21756 5516 21812
rect 5572 21756 7644 21812
rect 7700 21756 8876 21812
rect 8932 21756 8942 21812
rect 9874 21756 9884 21812
rect 9940 21756 9950 21812
rect 10108 21756 51884 21812
rect 51940 21756 51950 21812
rect 52098 21756 52108 21812
rect 52164 21756 52174 21812
rect 57932 21756 58884 21812
rect 58940 21756 59052 21812
rect 59108 21756 59500 21812
rect 59556 21756 59566 21812
rect 59724 21756 63756 21812
rect 63812 21756 64540 21812
rect 64596 21756 66108 21812
rect 66164 21756 66174 21812
rect 72146 21756 72156 21812
rect 72212 21756 75852 21812
rect 75908 21756 76860 21812
rect 76916 21756 76926 21812
rect 10108 21700 10164 21756
rect 58828 21700 58884 21756
rect 59724 21700 59780 21756
rect 2146 21644 2156 21700
rect 2212 21644 2604 21700
rect 2660 21644 2670 21700
rect 3938 21644 3948 21700
rect 4004 21644 4732 21700
rect 4788 21644 5404 21700
rect 5460 21644 6972 21700
rect 7028 21644 7038 21700
rect 7186 21644 7196 21700
rect 7252 21644 8204 21700
rect 8260 21644 8428 21700
rect 8530 21644 8540 21700
rect 8596 21644 10164 21700
rect 18162 21644 18172 21700
rect 18228 21644 20300 21700
rect 20356 21644 20366 21700
rect 21410 21644 21420 21700
rect 21476 21644 21868 21700
rect 21924 21644 22092 21700
rect 22148 21644 22158 21700
rect 23650 21644 23660 21700
rect 23716 21644 30716 21700
rect 30772 21644 30782 21700
rect 33954 21644 33964 21700
rect 34020 21644 35756 21700
rect 35812 21644 35822 21700
rect 37874 21644 37884 21700
rect 37940 21644 44268 21700
rect 44324 21644 44334 21700
rect 50306 21644 50316 21700
rect 50372 21644 52332 21700
rect 52388 21644 52398 21700
rect 58828 21644 59164 21700
rect 59220 21644 59780 21700
rect 60050 21644 60060 21700
rect 60116 21644 61516 21700
rect 61572 21644 61582 21700
rect 63298 21644 63308 21700
rect 63364 21644 64652 21700
rect 64708 21644 65548 21700
rect 65604 21644 65614 21700
rect 71698 21644 71708 21700
rect 71764 21644 74620 21700
rect 74676 21644 77308 21700
rect 77364 21644 77374 21700
rect 8372 21588 8428 21644
rect 6626 21532 6636 21588
rect 6692 21532 7308 21588
rect 7364 21532 7374 21588
rect 8372 21532 8764 21588
rect 8820 21532 8830 21588
rect 16146 21532 16156 21588
rect 16212 21532 16716 21588
rect 16772 21532 19516 21588
rect 19572 21532 21532 21588
rect 21588 21532 24892 21588
rect 24948 21532 26124 21588
rect 26180 21532 26190 21588
rect 26562 21532 26572 21588
rect 26628 21532 27580 21588
rect 27636 21532 27646 21588
rect 36530 21532 36540 21588
rect 36596 21532 37772 21588
rect 37828 21532 37838 21588
rect 46498 21532 46508 21588
rect 46564 21532 46956 21588
rect 47012 21532 47740 21588
rect 47796 21532 47806 21588
rect 48290 21532 48300 21588
rect 48356 21532 49868 21588
rect 49924 21532 49934 21588
rect 51874 21532 51884 21588
rect 51940 21532 55748 21588
rect 55906 21532 55916 21588
rect 55972 21532 61292 21588
rect 61348 21532 61740 21588
rect 61796 21532 61806 21588
rect 63970 21532 63980 21588
rect 64036 21532 64316 21588
rect 64372 21532 65436 21588
rect 65492 21532 65502 21588
rect 65650 21532 65660 21588
rect 65716 21532 65754 21588
rect 65874 21532 65884 21588
rect 65940 21532 66556 21588
rect 66612 21532 67116 21588
rect 67172 21532 67564 21588
rect 67620 21532 67630 21588
rect 73714 21532 73724 21588
rect 73780 21532 74396 21588
rect 74452 21532 74956 21588
rect 75012 21532 75022 21588
rect 55692 21476 55748 21532
rect 9874 21420 9884 21476
rect 9940 21420 15372 21476
rect 15428 21420 15438 21476
rect 19954 21420 19964 21476
rect 20020 21420 20748 21476
rect 20804 21420 21644 21476
rect 21700 21420 21710 21476
rect 22306 21420 22316 21476
rect 22372 21420 23100 21476
rect 23156 21420 23166 21476
rect 36306 21420 36316 21476
rect 36372 21420 37324 21476
rect 37380 21420 37390 21476
rect 39442 21420 39452 21476
rect 39508 21420 40124 21476
rect 40180 21420 40190 21476
rect 53778 21420 53788 21476
rect 53844 21420 54236 21476
rect 54292 21420 55020 21476
rect 55076 21420 55086 21476
rect 55692 21420 60508 21476
rect 60564 21420 60956 21476
rect 61012 21420 61022 21476
rect 66322 21420 66332 21476
rect 66388 21420 67452 21476
rect 67508 21420 67518 21476
rect 20178 21308 20188 21364
rect 20244 21308 20636 21364
rect 20692 21308 20702 21364
rect 0 21252 800 21280
rect 79200 21252 80000 21280
rect 0 21196 1932 21252
rect 1988 21196 1998 21252
rect 76066 21196 76076 21252
rect 76132 21196 80000 21252
rect 0 21168 800 21196
rect 10862 21140 10872 21196
rect 10928 21140 10976 21196
rect 11032 21140 11080 21196
rect 11136 21140 11146 21196
rect 30182 21140 30192 21196
rect 30248 21140 30296 21196
rect 30352 21140 30400 21196
rect 30456 21140 30466 21196
rect 49502 21140 49512 21196
rect 49568 21140 49616 21196
rect 49672 21140 49720 21196
rect 49776 21140 49786 21196
rect 68822 21140 68832 21196
rect 68888 21140 68936 21196
rect 68992 21140 69040 21196
rect 69096 21140 69106 21196
rect 79200 21168 80000 21196
rect 3154 20972 3164 21028
rect 3220 20972 10612 21028
rect 10770 20972 10780 21028
rect 10836 20972 22988 21028
rect 23044 20972 23548 21028
rect 23604 20972 24780 21028
rect 24836 20972 25788 21028
rect 25844 20972 25854 21028
rect 30594 20972 30604 21028
rect 30660 20972 31948 21028
rect 34962 20972 34972 21028
rect 35028 20972 36652 21028
rect 36708 20972 36718 21028
rect 55010 20972 55020 21028
rect 55076 20972 55804 21028
rect 55860 20972 55870 21028
rect 69906 20972 69916 21028
rect 69972 20972 70812 21028
rect 70868 20972 70878 21028
rect 74162 20972 74172 21028
rect 74228 20972 75068 21028
rect 75124 20972 75134 21028
rect 10556 20916 10612 20972
rect 3042 20860 3052 20916
rect 3108 20860 6524 20916
rect 6580 20860 6590 20916
rect 7634 20860 7644 20916
rect 7700 20860 8764 20916
rect 8820 20860 9324 20916
rect 9380 20860 9390 20916
rect 10556 20860 13356 20916
rect 13412 20860 13422 20916
rect 15092 20804 15148 20916
rect 15204 20860 19964 20916
rect 20020 20860 20030 20916
rect 20402 20860 20412 20916
rect 20468 20860 21868 20916
rect 21924 20860 21934 20916
rect 26002 20860 26012 20916
rect 26068 20860 27468 20916
rect 27524 20860 27534 20916
rect 31892 20804 31948 20972
rect 36194 20860 36204 20916
rect 36260 20860 38108 20916
rect 38164 20860 38668 20916
rect 38724 20860 38734 20916
rect 39218 20860 39228 20916
rect 39284 20860 41916 20916
rect 41972 20860 41982 20916
rect 56130 20860 56140 20916
rect 56196 20860 58716 20916
rect 58772 20860 59612 20916
rect 59668 20860 59678 20916
rect 65202 20860 65212 20916
rect 65268 20860 67788 20916
rect 67844 20860 67854 20916
rect 68002 20860 68012 20916
rect 68068 20860 69244 20916
rect 69300 20860 69580 20916
rect 69636 20860 72716 20916
rect 72772 20860 72782 20916
rect 74834 20860 74844 20916
rect 74900 20860 75516 20916
rect 75572 20860 77532 20916
rect 77588 20860 77598 20916
rect 7186 20748 7196 20804
rect 7252 20748 8204 20804
rect 8260 20748 8270 20804
rect 10658 20748 10668 20804
rect 10724 20748 11564 20804
rect 11620 20748 15148 20804
rect 17938 20748 17948 20804
rect 18004 20748 19852 20804
rect 19908 20748 19918 20804
rect 20860 20748 22092 20804
rect 22148 20748 23660 20804
rect 23716 20748 23726 20804
rect 24210 20748 24220 20804
rect 24276 20748 25116 20804
rect 25172 20748 25182 20804
rect 31892 20748 36148 20804
rect 48402 20748 48412 20804
rect 48468 20748 49644 20804
rect 49700 20748 49710 20804
rect 54338 20748 54348 20804
rect 54404 20748 55580 20804
rect 55636 20748 55646 20804
rect 58594 20748 58604 20804
rect 58660 20748 60060 20804
rect 60116 20748 60126 20804
rect 60386 20748 60396 20804
rect 60452 20748 61628 20804
rect 61684 20748 61694 20804
rect 61842 20748 61852 20804
rect 61908 20748 62972 20804
rect 63028 20748 63038 20804
rect 65538 20748 65548 20804
rect 65604 20748 66108 20804
rect 66164 20748 66668 20804
rect 66724 20748 66734 20804
rect 69794 20748 69804 20804
rect 69860 20748 70364 20804
rect 70420 20748 70430 20804
rect 73714 20748 73724 20804
rect 73780 20748 77868 20804
rect 77924 20748 77934 20804
rect 20860 20692 20916 20748
rect 36092 20692 36148 20748
rect 4946 20636 4956 20692
rect 5012 20636 6076 20692
rect 6132 20636 6142 20692
rect 9202 20636 9212 20692
rect 9268 20636 9884 20692
rect 9940 20636 9950 20692
rect 10546 20636 10556 20692
rect 10612 20636 11116 20692
rect 11172 20636 14028 20692
rect 14084 20636 14094 20692
rect 18610 20636 18620 20692
rect 18676 20636 19628 20692
rect 19684 20636 20860 20692
rect 20916 20636 20926 20692
rect 25554 20636 25564 20692
rect 25620 20636 26460 20692
rect 26516 20636 26526 20692
rect 26852 20636 29036 20692
rect 29092 20636 29708 20692
rect 29764 20636 35700 20692
rect 36082 20636 36092 20692
rect 36148 20636 36158 20692
rect 44594 20636 44604 20692
rect 44660 20636 48300 20692
rect 48356 20636 48366 20692
rect 55906 20636 55916 20692
rect 55972 20636 56364 20692
rect 56420 20636 61964 20692
rect 62020 20636 62030 20692
rect 65314 20636 65324 20692
rect 65380 20636 65772 20692
rect 65828 20636 65838 20692
rect 68226 20636 68236 20692
rect 68292 20636 71708 20692
rect 71764 20636 72268 20692
rect 72324 20636 72334 20692
rect 26852 20580 26908 20636
rect 12002 20524 12012 20580
rect 12068 20524 13020 20580
rect 13076 20524 13916 20580
rect 13972 20524 13982 20580
rect 17714 20524 17724 20580
rect 17780 20524 18732 20580
rect 18788 20524 18798 20580
rect 25106 20524 25116 20580
rect 25172 20524 26572 20580
rect 26628 20524 26908 20580
rect 27794 20524 27804 20580
rect 27860 20524 32732 20580
rect 32788 20524 32798 20580
rect 35644 20468 35700 20636
rect 35858 20524 35868 20580
rect 35924 20524 39900 20580
rect 39956 20524 39966 20580
rect 44370 20524 44380 20580
rect 44436 20524 45388 20580
rect 45444 20524 45454 20580
rect 53554 20524 53564 20580
rect 53620 20524 54348 20580
rect 54404 20524 55468 20580
rect 55524 20524 56140 20580
rect 56196 20524 56206 20580
rect 69458 20524 69468 20580
rect 69524 20524 69804 20580
rect 69860 20524 69870 20580
rect 70466 20524 70476 20580
rect 70532 20524 70924 20580
rect 70980 20524 70990 20580
rect 73938 20524 73948 20580
rect 74004 20524 75180 20580
rect 75236 20524 77308 20580
rect 77364 20524 77374 20580
rect 4834 20412 4844 20468
rect 4900 20412 5628 20468
rect 5684 20412 10780 20468
rect 10836 20412 10846 20468
rect 21634 20412 21644 20468
rect 21700 20412 24556 20468
rect 24612 20412 26124 20468
rect 26180 20412 26190 20468
rect 27458 20412 27468 20468
rect 27524 20412 31948 20468
rect 35644 20412 37772 20468
rect 37828 20412 39116 20468
rect 39172 20412 39732 20468
rect 67218 20412 67228 20468
rect 67284 20412 71148 20468
rect 71204 20412 71214 20468
rect 20522 20356 20532 20412
rect 20588 20356 20636 20412
rect 20692 20356 20740 20412
rect 20796 20356 20806 20412
rect 31892 20356 31948 20412
rect 18274 20300 18284 20356
rect 18340 20300 19460 20356
rect 26450 20300 26460 20356
rect 26516 20300 28364 20356
rect 28420 20300 28812 20356
rect 28868 20300 29596 20356
rect 29652 20300 29662 20356
rect 31892 20300 39452 20356
rect 39508 20300 39518 20356
rect 19404 20244 19460 20300
rect 39676 20244 39732 20412
rect 39842 20356 39852 20412
rect 39908 20356 39956 20412
rect 40012 20356 40060 20412
rect 40116 20356 40126 20412
rect 59162 20356 59172 20412
rect 59228 20356 59276 20412
rect 59332 20356 59380 20412
rect 59436 20356 59446 20412
rect 78482 20356 78492 20412
rect 78548 20356 78596 20412
rect 78652 20356 78700 20412
rect 78756 20356 78766 20412
rect 48514 20300 48524 20356
rect 48580 20300 50092 20356
rect 50148 20300 50158 20356
rect 69458 20300 69468 20356
rect 69524 20300 71596 20356
rect 71652 20300 71662 20356
rect 18386 20188 18396 20244
rect 18452 20188 18462 20244
rect 19394 20188 19404 20244
rect 19460 20188 20076 20244
rect 20132 20188 20860 20244
rect 20916 20188 21756 20244
rect 21812 20188 21822 20244
rect 22530 20188 22540 20244
rect 22596 20188 22606 20244
rect 25778 20188 25788 20244
rect 25844 20188 27468 20244
rect 27524 20188 27534 20244
rect 27794 20188 27804 20244
rect 27860 20188 29148 20244
rect 29204 20188 30828 20244
rect 30884 20188 30894 20244
rect 39676 20188 40908 20244
rect 40964 20188 40974 20244
rect 47618 20188 47628 20244
rect 47684 20188 48412 20244
rect 48468 20188 48478 20244
rect 18396 20132 18452 20188
rect 22540 20132 22596 20188
rect 3490 20076 3500 20132
rect 3556 20076 4620 20132
rect 4676 20076 4686 20132
rect 8306 20076 8316 20132
rect 8372 20076 10108 20132
rect 10164 20076 10174 20132
rect 13010 20076 13020 20132
rect 13076 20076 14252 20132
rect 14308 20076 14318 20132
rect 18396 20076 19516 20132
rect 19572 20076 19582 20132
rect 21522 20076 21532 20132
rect 21588 20076 22596 20132
rect 24658 20076 24668 20132
rect 24724 20076 33012 20132
rect 33170 20076 33180 20132
rect 33236 20076 35196 20132
rect 35252 20076 35262 20132
rect 38098 20076 38108 20132
rect 38164 20076 38668 20132
rect 39554 20076 39564 20132
rect 39620 20076 40348 20132
rect 40404 20076 41804 20132
rect 41860 20076 41870 20132
rect 44706 20076 44716 20132
rect 44772 20076 46508 20132
rect 46564 20076 46574 20132
rect 62402 20076 62412 20132
rect 62468 20076 63084 20132
rect 63140 20076 63868 20132
rect 63924 20076 70028 20132
rect 70084 20076 70094 20132
rect 74610 20076 74620 20132
rect 74676 20076 76972 20132
rect 77028 20076 77038 20132
rect 77522 20076 77532 20132
rect 77588 20076 78988 20132
rect 79044 20076 79054 20132
rect 32956 20020 33012 20076
rect 1810 19964 1820 20020
rect 1876 19964 2380 20020
rect 2436 19964 3388 20020
rect 3444 19964 3454 20020
rect 3714 19964 3724 20020
rect 3780 19964 5068 20020
rect 5124 19964 5134 20020
rect 14130 19964 14140 20020
rect 14196 19964 15036 20020
rect 15092 19964 15102 20020
rect 17490 19964 17500 20020
rect 17556 19964 19180 20020
rect 19236 19964 19246 20020
rect 23538 19964 23548 20020
rect 23604 19964 24332 20020
rect 24388 19964 24398 20020
rect 32956 19964 37660 20020
rect 37716 19964 37726 20020
rect 38612 19964 38668 20076
rect 38724 19964 39676 20020
rect 39732 19964 39742 20020
rect 40674 19964 40684 20020
rect 40740 19964 42140 20020
rect 42196 19964 42206 20020
rect 44146 19964 44156 20020
rect 44212 19964 46172 20020
rect 46228 19964 46238 20020
rect 48066 19964 48076 20020
rect 48132 19964 49532 20020
rect 49588 19964 50988 20020
rect 51044 19964 51054 20020
rect 53554 19964 53564 20020
rect 53620 19964 54460 20020
rect 54516 19964 55804 20020
rect 55860 19964 55870 20020
rect 59938 19964 59948 20020
rect 60004 19964 63644 20020
rect 63700 19964 64204 20020
rect 64260 19964 64270 20020
rect 69010 19964 69020 20020
rect 69076 19964 69916 20020
rect 69972 19964 70812 20020
rect 70868 19964 70878 20020
rect 71250 19964 71260 20020
rect 71316 19964 72044 20020
rect 72100 19964 72110 20020
rect 74386 19964 74396 20020
rect 74452 19964 75292 20020
rect 75348 19964 75358 20020
rect 3602 19852 3612 19908
rect 3668 19852 4844 19908
rect 4900 19852 4910 19908
rect 13906 19852 13916 19908
rect 13972 19852 15148 19908
rect 15204 19852 15214 19908
rect 26898 19852 26908 19908
rect 26964 19852 27692 19908
rect 27748 19852 29036 19908
rect 29092 19852 29596 19908
rect 29652 19852 29662 19908
rect 31154 19852 31164 19908
rect 31220 19852 32788 19908
rect 34626 19852 34636 19908
rect 34692 19852 35196 19908
rect 35252 19852 35262 19908
rect 43362 19852 43372 19908
rect 43428 19852 43932 19908
rect 43988 19852 43998 19908
rect 45490 19852 45500 19908
rect 45556 19852 48636 19908
rect 48692 19852 48702 19908
rect 64754 19852 64764 19908
rect 64820 19852 66332 19908
rect 66388 19852 66398 19908
rect 66994 19852 67004 19908
rect 67060 19852 67900 19908
rect 67956 19852 67966 19908
rect 68674 19852 68684 19908
rect 68740 19852 69356 19908
rect 69412 19852 69692 19908
rect 69748 19852 70252 19908
rect 70308 19852 70318 19908
rect 71922 19852 71932 19908
rect 71988 19852 72492 19908
rect 72548 19852 72558 19908
rect 74274 19852 74284 19908
rect 74340 19852 74732 19908
rect 74788 19852 75404 19908
rect 75460 19852 75470 19908
rect 6738 19740 6748 19796
rect 6804 19740 22204 19796
rect 22260 19740 22270 19796
rect 27906 19740 27916 19796
rect 27972 19740 28252 19796
rect 28308 19740 30604 19796
rect 30660 19740 30670 19796
rect 32732 19684 32788 19852
rect 43932 19796 43988 19852
rect 43932 19740 46284 19796
rect 46340 19740 46844 19796
rect 46900 19740 46910 19796
rect 52322 19740 52332 19796
rect 52388 19740 63980 19796
rect 64036 19740 64046 19796
rect 72034 19740 72044 19796
rect 72100 19740 73276 19796
rect 73332 19740 73836 19796
rect 73892 19740 73902 19796
rect 74050 19740 74060 19796
rect 74116 19740 75628 19796
rect 75684 19740 77084 19796
rect 77140 19740 77150 19796
rect 32732 19628 33740 19684
rect 33796 19628 35308 19684
rect 35364 19628 35374 19684
rect 35522 19628 35532 19684
rect 35588 19628 36092 19684
rect 36148 19628 36158 19684
rect 37090 19628 37100 19684
rect 37156 19628 47068 19684
rect 47124 19628 47134 19684
rect 10862 19572 10872 19628
rect 10928 19572 10976 19628
rect 11032 19572 11080 19628
rect 11136 19572 11146 19628
rect 30182 19572 30192 19628
rect 30248 19572 30296 19628
rect 30352 19572 30400 19628
rect 30456 19572 30466 19628
rect 49502 19572 49512 19628
rect 49568 19572 49616 19628
rect 49672 19572 49720 19628
rect 49776 19572 49786 19628
rect 14242 19516 14252 19572
rect 14308 19516 16156 19572
rect 16212 19516 16222 19572
rect 18620 19516 25900 19572
rect 25956 19516 26348 19572
rect 26404 19516 26414 19572
rect 33506 19516 33516 19572
rect 33572 19516 45276 19572
rect 45332 19516 45342 19572
rect 53218 19516 53228 19572
rect 53284 19516 53294 19572
rect 18620 19460 18676 19516
rect 53228 19460 53284 19516
rect 4946 19404 4956 19460
rect 5012 19404 5964 19460
rect 6020 19404 6030 19460
rect 8372 19404 8540 19460
rect 8596 19404 8606 19460
rect 9426 19404 9436 19460
rect 9492 19404 9884 19460
rect 9940 19404 9950 19460
rect 13794 19404 13804 19460
rect 13860 19404 14700 19460
rect 14756 19404 18620 19460
rect 18676 19404 18686 19460
rect 18834 19404 18844 19460
rect 18900 19404 19068 19460
rect 19124 19404 20972 19460
rect 21028 19404 21308 19460
rect 21364 19404 22316 19460
rect 22372 19404 22652 19460
rect 22708 19404 22718 19460
rect 24770 19404 24780 19460
rect 24836 19404 26236 19460
rect 26292 19404 26302 19460
rect 49634 19404 49644 19460
rect 49700 19404 53788 19460
rect 53844 19404 53854 19460
rect 8372 19348 8428 19404
rect 63980 19348 64036 19740
rect 74162 19628 74172 19684
rect 74228 19628 76636 19684
rect 76692 19628 76702 19684
rect 68822 19572 68832 19628
rect 68888 19572 68936 19628
rect 68992 19572 69040 19628
rect 69096 19572 69106 19628
rect 3938 19292 3948 19348
rect 4004 19292 4620 19348
rect 4676 19292 8428 19348
rect 15026 19292 15036 19348
rect 15092 19292 16940 19348
rect 16996 19292 17006 19348
rect 17266 19292 17276 19348
rect 17332 19292 19628 19348
rect 19684 19292 19694 19348
rect 28690 19292 28700 19348
rect 28756 19292 38724 19348
rect 39890 19292 39900 19348
rect 39956 19292 41020 19348
rect 41076 19292 41086 19348
rect 42690 19292 42700 19348
rect 42756 19292 43596 19348
rect 43652 19292 43662 19348
rect 49858 19292 49868 19348
rect 49924 19292 51100 19348
rect 51156 19292 51166 19348
rect 56578 19292 56588 19348
rect 56644 19292 57820 19348
rect 57876 19292 57886 19348
rect 63970 19292 63980 19348
rect 64036 19292 64046 19348
rect 73826 19292 73836 19348
rect 73892 19292 74396 19348
rect 74452 19292 74462 19348
rect 38668 19236 38724 19292
rect 4834 19180 4844 19236
rect 4900 19180 6076 19236
rect 6132 19180 6142 19236
rect 8866 19180 8876 19236
rect 8932 19180 9660 19236
rect 9716 19180 9726 19236
rect 16594 19180 16604 19236
rect 16660 19180 17052 19236
rect 17108 19180 17118 19236
rect 19730 19180 19740 19236
rect 19796 19180 21532 19236
rect 21588 19180 21598 19236
rect 22194 19180 22204 19236
rect 22260 19180 23436 19236
rect 23492 19180 23502 19236
rect 24994 19180 25004 19236
rect 25060 19180 26348 19236
rect 26404 19180 26414 19236
rect 30930 19180 30940 19236
rect 30996 19180 34076 19236
rect 34132 19180 34636 19236
rect 34692 19180 34702 19236
rect 38658 19180 38668 19236
rect 38724 19180 39004 19236
rect 39060 19180 40460 19236
rect 40516 19180 40526 19236
rect 58034 19180 58044 19236
rect 58100 19180 58492 19236
rect 58548 19180 59388 19236
rect 59444 19180 59454 19236
rect 60162 19180 60172 19236
rect 60228 19180 61516 19236
rect 61572 19180 61582 19236
rect 63186 19180 63196 19236
rect 63252 19180 64092 19236
rect 64148 19180 64158 19236
rect 64306 19180 64316 19236
rect 64372 19180 66780 19236
rect 66836 19180 66846 19236
rect 76178 19180 76188 19236
rect 76244 19180 77196 19236
rect 77252 19180 77262 19236
rect 3042 19068 3052 19124
rect 3108 19068 3612 19124
rect 3668 19068 3678 19124
rect 18162 19068 18172 19124
rect 18228 19068 18620 19124
rect 18676 19068 18686 19124
rect 20178 19068 20188 19124
rect 20244 19068 20860 19124
rect 20916 19068 21980 19124
rect 22036 19068 22764 19124
rect 22820 19068 22830 19124
rect 24098 19068 24108 19124
rect 24164 19068 26236 19124
rect 26292 19068 26302 19124
rect 26898 19068 26908 19124
rect 26964 19068 27468 19124
rect 27524 19068 27534 19124
rect 30482 19068 30492 19124
rect 30548 19068 31724 19124
rect 31780 19068 31790 19124
rect 34738 19068 34748 19124
rect 34804 19068 35980 19124
rect 36036 19068 36046 19124
rect 37202 19068 37212 19124
rect 37268 19068 40348 19124
rect 40404 19068 41580 19124
rect 41636 19068 62188 19124
rect 64194 19068 64204 19124
rect 64260 19068 65436 19124
rect 65492 19068 65502 19124
rect 67554 19068 67564 19124
rect 67620 19068 69356 19124
rect 69412 19068 70476 19124
rect 70532 19068 70542 19124
rect 62132 19012 62188 19068
rect 16482 18956 16492 19012
rect 16548 18956 19628 19012
rect 19684 18956 20412 19012
rect 20468 18956 21028 19012
rect 21186 18956 21196 19012
rect 21252 18956 31500 19012
rect 31556 18956 32172 19012
rect 32228 18956 33516 19012
rect 33572 18956 33582 19012
rect 39890 18956 39900 19012
rect 39956 18956 40572 19012
rect 40628 18956 42588 19012
rect 42644 18956 42654 19012
rect 50194 18956 50204 19012
rect 50260 18956 50764 19012
rect 50820 18956 50830 19012
rect 62132 18956 62748 19012
rect 62804 18956 62814 19012
rect 68674 18956 68684 19012
rect 68740 18956 69468 19012
rect 69524 18956 70364 19012
rect 70420 18956 71708 19012
rect 71764 18956 71774 19012
rect 75506 18956 75516 19012
rect 75572 18956 78932 19012
rect 18498 18844 18508 18900
rect 18564 18844 18574 18900
rect 0 18788 800 18816
rect 18508 18788 18564 18844
rect 20522 18788 20532 18844
rect 20588 18788 20636 18844
rect 20692 18788 20740 18844
rect 20796 18788 20806 18844
rect 20972 18788 21028 18956
rect 26002 18844 26012 18900
rect 26068 18844 28252 18900
rect 28308 18844 28700 18900
rect 28756 18844 28766 18900
rect 29586 18844 29596 18900
rect 29652 18844 31388 18900
rect 31444 18844 31454 18900
rect 36418 18844 36428 18900
rect 36484 18844 39116 18900
rect 39172 18844 39732 18900
rect 40226 18844 40236 18900
rect 40292 18844 50316 18900
rect 50372 18844 50382 18900
rect 0 18732 1932 18788
rect 1988 18732 1998 18788
rect 8306 18732 8316 18788
rect 0 18704 800 18732
rect 8372 18676 8428 18788
rect 15138 18732 15148 18788
rect 15204 18732 16268 18788
rect 16324 18732 16334 18788
rect 16930 18732 16940 18788
rect 16996 18732 17164 18788
rect 17220 18732 18564 18788
rect 18722 18732 18732 18788
rect 18788 18732 19740 18788
rect 19796 18732 19806 18788
rect 20972 18732 36708 18788
rect 36652 18676 36708 18732
rect 39676 18676 39732 18844
rect 39842 18788 39852 18844
rect 39908 18788 39956 18844
rect 40012 18788 40060 18844
rect 40116 18788 40126 18844
rect 59162 18788 59172 18844
rect 59228 18788 59276 18844
rect 59332 18788 59380 18844
rect 59436 18788 59446 18844
rect 78482 18788 78492 18844
rect 78548 18788 78596 18844
rect 78652 18788 78700 18844
rect 78756 18788 78766 18844
rect 78876 18788 78932 18956
rect 79200 18788 80000 18816
rect 41010 18732 41020 18788
rect 41076 18732 41692 18788
rect 41748 18732 41916 18788
rect 41972 18732 41982 18788
rect 49298 18732 49308 18788
rect 49364 18732 49868 18788
rect 49924 18732 49934 18788
rect 50866 18732 50876 18788
rect 50932 18732 51324 18788
rect 51380 18732 52444 18788
rect 52500 18732 52510 18788
rect 58146 18732 58156 18788
rect 58212 18732 58940 18788
rect 58996 18732 59006 18788
rect 78876 18732 80000 18788
rect 79200 18704 80000 18732
rect 2370 18620 2380 18676
rect 2436 18620 2716 18676
rect 2772 18620 3836 18676
rect 3892 18620 3902 18676
rect 8372 18620 8876 18676
rect 8932 18620 9884 18676
rect 9940 18620 10556 18676
rect 10612 18620 14252 18676
rect 14308 18620 14318 18676
rect 16370 18620 16380 18676
rect 16436 18620 16828 18676
rect 16884 18620 16894 18676
rect 18050 18620 18060 18676
rect 18116 18620 19516 18676
rect 19572 18620 19582 18676
rect 20178 18620 20188 18676
rect 20244 18620 21196 18676
rect 21252 18620 21262 18676
rect 23426 18620 23436 18676
rect 23492 18620 24108 18676
rect 24164 18620 24174 18676
rect 31378 18620 31388 18676
rect 31444 18620 33852 18676
rect 33908 18620 33918 18676
rect 36642 18620 36652 18676
rect 36708 18620 37100 18676
rect 37156 18620 37166 18676
rect 37650 18620 37660 18676
rect 37716 18620 38892 18676
rect 38948 18620 39228 18676
rect 39284 18620 39294 18676
rect 39676 18620 40124 18676
rect 40180 18620 40190 18676
rect 40348 18620 43372 18676
rect 43428 18620 43438 18676
rect 45826 18620 45836 18676
rect 45892 18620 48188 18676
rect 48244 18620 49756 18676
rect 49812 18620 49822 18676
rect 51650 18620 51660 18676
rect 51716 18620 52332 18676
rect 52388 18620 52398 18676
rect 55346 18620 55356 18676
rect 55412 18620 56252 18676
rect 56308 18620 56318 18676
rect 58258 18620 58268 18676
rect 58324 18620 59164 18676
rect 59220 18620 59230 18676
rect 59378 18620 59388 18676
rect 59444 18620 60172 18676
rect 60228 18620 60238 18676
rect 66098 18620 66108 18676
rect 66164 18620 67228 18676
rect 67284 18620 68012 18676
rect 68068 18620 68078 18676
rect 40348 18564 40404 18620
rect 1922 18508 1932 18564
rect 1988 18508 3164 18564
rect 3220 18508 3230 18564
rect 11442 18508 11452 18564
rect 11508 18508 13244 18564
rect 13300 18508 13310 18564
rect 15810 18508 15820 18564
rect 15876 18508 17836 18564
rect 17892 18508 18620 18564
rect 18676 18508 19292 18564
rect 19348 18508 20076 18564
rect 20132 18508 20142 18564
rect 22194 18508 22204 18564
rect 22260 18508 23548 18564
rect 23604 18508 23614 18564
rect 25666 18508 25676 18564
rect 25732 18508 25742 18564
rect 29922 18508 29932 18564
rect 29988 18508 31052 18564
rect 31108 18508 31118 18564
rect 34738 18508 34748 18564
rect 34804 18508 40404 18564
rect 40460 18508 42364 18564
rect 42420 18508 42430 18564
rect 43586 18508 43596 18564
rect 43652 18508 68124 18564
rect 68180 18508 68190 18564
rect 70130 18508 70140 18564
rect 70196 18508 71372 18564
rect 71428 18508 71438 18564
rect 73714 18508 73724 18564
rect 73780 18508 77532 18564
rect 77588 18508 77598 18564
rect 25676 18452 25732 18508
rect 40460 18452 40516 18508
rect 5394 18396 5404 18452
rect 5460 18396 6524 18452
rect 6580 18396 9548 18452
rect 9604 18396 9614 18452
rect 10210 18396 10220 18452
rect 10276 18396 11564 18452
rect 11620 18396 11630 18452
rect 16370 18396 16380 18452
rect 16436 18396 16716 18452
rect 16772 18396 16782 18452
rect 17042 18396 17052 18452
rect 17108 18396 18396 18452
rect 18452 18396 18462 18452
rect 24882 18396 24892 18452
rect 24948 18396 25732 18452
rect 25890 18396 25900 18452
rect 25956 18396 26684 18452
rect 26740 18396 27132 18452
rect 27188 18396 27580 18452
rect 27636 18396 27804 18452
rect 27860 18396 27870 18452
rect 28018 18396 28028 18452
rect 28084 18396 30156 18452
rect 30212 18396 32172 18452
rect 32228 18396 32238 18452
rect 38658 18396 38668 18452
rect 38724 18396 39452 18452
rect 39508 18396 39518 18452
rect 40450 18396 40460 18452
rect 40516 18396 40526 18452
rect 40786 18396 40796 18452
rect 40852 18396 41580 18452
rect 41636 18396 42252 18452
rect 42308 18396 43708 18452
rect 43764 18396 43774 18452
rect 44930 18396 44940 18452
rect 44996 18396 45500 18452
rect 45556 18396 45836 18452
rect 45892 18396 45902 18452
rect 47058 18396 47068 18452
rect 47124 18396 47852 18452
rect 47908 18396 50652 18452
rect 50708 18396 50718 18452
rect 51090 18396 51100 18452
rect 51156 18396 53788 18452
rect 53844 18396 54796 18452
rect 54852 18396 54862 18452
rect 59714 18396 59724 18452
rect 59780 18396 61292 18452
rect 61348 18396 61358 18452
rect 64754 18396 64764 18452
rect 64820 18396 65884 18452
rect 65940 18396 65950 18452
rect 70690 18396 70700 18452
rect 70756 18396 72156 18452
rect 72212 18396 74620 18452
rect 74676 18396 74686 18452
rect 76738 18396 76748 18452
rect 76804 18396 77756 18452
rect 77812 18396 77822 18452
rect 7858 18284 7868 18340
rect 7924 18284 8988 18340
rect 9044 18284 9054 18340
rect 10098 18284 10108 18340
rect 10164 18284 11340 18340
rect 11396 18284 11406 18340
rect 13458 18284 13468 18340
rect 13524 18284 20972 18340
rect 21028 18284 21868 18340
rect 21924 18284 23324 18340
rect 23380 18284 23390 18340
rect 22764 18228 22820 18284
rect 25676 18228 25732 18396
rect 50652 18340 50708 18396
rect 28354 18284 28364 18340
rect 28420 18284 28588 18340
rect 28644 18284 28654 18340
rect 30594 18284 30604 18340
rect 30660 18284 31276 18340
rect 31332 18284 32284 18340
rect 32340 18284 32350 18340
rect 37986 18284 37996 18340
rect 38052 18284 39004 18340
rect 39060 18284 41636 18340
rect 41794 18284 41804 18340
rect 41860 18284 42588 18340
rect 42644 18284 43484 18340
rect 43540 18284 43550 18340
rect 50652 18284 51436 18340
rect 51492 18284 51502 18340
rect 54114 18284 54124 18340
rect 54180 18284 55020 18340
rect 55076 18284 55468 18340
rect 55524 18284 55534 18340
rect 61170 18284 61180 18340
rect 61236 18284 65772 18340
rect 65828 18284 66668 18340
rect 66724 18284 66734 18340
rect 68338 18284 68348 18340
rect 68404 18284 68908 18340
rect 68964 18284 68974 18340
rect 73826 18284 73836 18340
rect 73892 18284 76076 18340
rect 76132 18284 77420 18340
rect 77476 18284 77486 18340
rect 41580 18228 41636 18284
rect 51436 18228 51492 18284
rect 9762 18172 9772 18228
rect 9828 18172 10444 18228
rect 10500 18172 12348 18228
rect 12404 18172 12414 18228
rect 15362 18172 15372 18228
rect 15428 18172 21420 18228
rect 21476 18172 21486 18228
rect 22754 18172 22764 18228
rect 22820 18172 22830 18228
rect 25676 18172 33628 18228
rect 33684 18172 33694 18228
rect 35634 18172 35644 18228
rect 35700 18172 39788 18228
rect 39844 18172 39854 18228
rect 41580 18172 51212 18228
rect 51268 18172 51278 18228
rect 51436 18172 60732 18228
rect 60788 18172 60798 18228
rect 63410 18172 63420 18228
rect 63476 18172 69580 18228
rect 69636 18172 69646 18228
rect 74050 18172 74060 18228
rect 74116 18172 75180 18228
rect 75236 18172 75246 18228
rect 14578 18060 14588 18116
rect 14644 18060 15148 18116
rect 15250 18060 15260 18116
rect 15316 18060 16940 18116
rect 16996 18060 17006 18116
rect 34178 18060 34188 18116
rect 34244 18060 35308 18116
rect 35364 18060 38668 18116
rect 39330 18060 39340 18116
rect 39396 18060 39406 18116
rect 42578 18060 42588 18116
rect 42644 18060 44492 18116
rect 44548 18060 44558 18116
rect 10862 18004 10872 18060
rect 10928 18004 10976 18060
rect 11032 18004 11080 18060
rect 11136 18004 11146 18060
rect 15092 18004 15148 18060
rect 30182 18004 30192 18060
rect 30248 18004 30296 18060
rect 30352 18004 30400 18060
rect 30456 18004 30466 18060
rect 38612 18004 38668 18060
rect 39340 18004 39396 18060
rect 49502 18004 49512 18060
rect 49568 18004 49616 18060
rect 49672 18004 49720 18060
rect 49776 18004 49786 18060
rect 68822 18004 68832 18060
rect 68888 18004 68936 18060
rect 68992 18004 69040 18060
rect 69096 18004 69106 18060
rect 15092 17948 19740 18004
rect 19796 17948 19806 18004
rect 38612 17948 43876 18004
rect 43820 17892 43876 17948
rect 3938 17836 3948 17892
rect 4004 17836 4956 17892
rect 5012 17836 5740 17892
rect 5796 17836 5806 17892
rect 8754 17836 8764 17892
rect 8820 17836 9660 17892
rect 9716 17836 11676 17892
rect 11732 17836 12460 17892
rect 12516 17836 12526 17892
rect 18162 17836 18172 17892
rect 18228 17836 18508 17892
rect 18564 17836 19180 17892
rect 19236 17836 19246 17892
rect 20402 17836 20412 17892
rect 20468 17836 43596 17892
rect 43652 17836 43662 17892
rect 43820 17836 49980 17892
rect 50036 17836 50046 17892
rect 20412 17780 20468 17836
rect 7970 17724 7980 17780
rect 8036 17724 8428 17780
rect 8484 17724 8494 17780
rect 8652 17724 15932 17780
rect 15988 17724 15998 17780
rect 18722 17724 18732 17780
rect 18788 17724 19068 17780
rect 19124 17724 19964 17780
rect 20020 17724 20468 17780
rect 33618 17724 33628 17780
rect 33684 17724 34524 17780
rect 34580 17724 35196 17780
rect 35252 17724 36540 17780
rect 36596 17724 36606 17780
rect 39666 17724 39676 17780
rect 39732 17724 41692 17780
rect 41748 17724 45724 17780
rect 45780 17724 45790 17780
rect 51202 17724 51212 17780
rect 51268 17724 53340 17780
rect 53396 17724 53406 17780
rect 63186 17724 63196 17780
rect 63252 17724 67228 17780
rect 67284 17724 68348 17780
rect 68404 17724 68414 17780
rect 75170 17724 75180 17780
rect 75236 17724 77308 17780
rect 77364 17724 77374 17780
rect 8652 17668 8708 17724
rect 6962 17612 6972 17668
rect 7028 17612 8708 17668
rect 8866 17612 8876 17668
rect 8932 17612 10220 17668
rect 10276 17612 10286 17668
rect 14354 17612 14364 17668
rect 14420 17612 17724 17668
rect 17780 17612 25228 17668
rect 25284 17612 28812 17668
rect 28868 17612 29148 17668
rect 29204 17612 29214 17668
rect 36754 17612 36764 17668
rect 36820 17612 37548 17668
rect 37604 17612 37884 17668
rect 37940 17612 37950 17668
rect 38882 17612 38892 17668
rect 38948 17612 39340 17668
rect 39396 17612 39406 17668
rect 46946 17612 46956 17668
rect 47012 17612 47516 17668
rect 47572 17612 47582 17668
rect 50306 17612 50316 17668
rect 50372 17612 56308 17668
rect 62066 17612 62076 17668
rect 62132 17612 69356 17668
rect 69412 17612 69422 17668
rect 69794 17612 69804 17668
rect 69860 17612 71260 17668
rect 71316 17612 71326 17668
rect 74610 17612 74620 17668
rect 74676 17612 76076 17668
rect 76132 17612 76748 17668
rect 76804 17612 76814 17668
rect 8530 17500 8540 17556
rect 8596 17500 11788 17556
rect 11844 17500 12572 17556
rect 12628 17500 15148 17556
rect 26338 17500 26348 17556
rect 26404 17500 32844 17556
rect 32900 17500 32910 17556
rect 38612 17500 50764 17556
rect 50820 17500 51436 17556
rect 51492 17500 53676 17556
rect 53732 17500 53742 17556
rect 2146 17388 2156 17444
rect 2212 17388 2604 17444
rect 2660 17388 4060 17444
rect 4116 17388 4956 17444
rect 5012 17388 5022 17444
rect 12450 17388 12460 17444
rect 12516 17388 12796 17444
rect 12852 17388 13804 17444
rect 13860 17388 14476 17444
rect 14532 17388 14812 17444
rect 14868 17388 14878 17444
rect 15092 17332 15148 17500
rect 38612 17444 38668 17500
rect 56252 17444 56308 17612
rect 58034 17500 58044 17556
rect 58100 17500 59500 17556
rect 59556 17500 59566 17556
rect 60386 17500 60396 17556
rect 60452 17500 61740 17556
rect 61796 17500 61806 17556
rect 69682 17500 69692 17556
rect 69748 17500 70140 17556
rect 70196 17500 70364 17556
rect 70420 17500 71036 17556
rect 71092 17500 71102 17556
rect 73938 17500 73948 17556
rect 74004 17500 74508 17556
rect 74564 17500 75628 17556
rect 75684 17500 75694 17556
rect 25890 17388 25900 17444
rect 25956 17388 26460 17444
rect 26516 17388 26526 17444
rect 27458 17388 27468 17444
rect 27524 17388 29596 17444
rect 29652 17388 30156 17444
rect 30212 17388 30222 17444
rect 31892 17388 38668 17444
rect 39218 17388 39228 17444
rect 39284 17388 40348 17444
rect 40404 17388 40414 17444
rect 40562 17388 40572 17444
rect 40628 17388 42028 17444
rect 42084 17388 42094 17444
rect 47170 17388 47180 17444
rect 47236 17388 47740 17444
rect 47796 17388 47806 17444
rect 50530 17388 50540 17444
rect 50596 17388 52220 17444
rect 52276 17388 52286 17444
rect 56252 17388 64652 17444
rect 64708 17388 65324 17444
rect 65380 17388 65390 17444
rect 70242 17388 70252 17444
rect 70308 17388 71484 17444
rect 71540 17388 71550 17444
rect 75170 17388 75180 17444
rect 75236 17388 75516 17444
rect 75572 17388 78876 17444
rect 78932 17388 78942 17444
rect 31892 17332 31948 17388
rect 51324 17332 51380 17388
rect 15092 17276 15372 17332
rect 15428 17276 19628 17332
rect 19684 17276 20188 17332
rect 20244 17276 20254 17332
rect 26562 17276 26572 17332
rect 26628 17276 31948 17332
rect 32834 17276 32844 17332
rect 32900 17276 33516 17332
rect 33572 17276 37268 17332
rect 40226 17276 40236 17332
rect 40292 17276 40908 17332
rect 40964 17276 40974 17332
rect 51314 17276 51324 17332
rect 51380 17276 51390 17332
rect 58034 17276 58044 17332
rect 58100 17276 58604 17332
rect 58660 17276 58670 17332
rect 77410 17276 77420 17332
rect 77476 17276 77756 17332
rect 77812 17276 77822 17332
rect 20522 17220 20532 17276
rect 20588 17220 20636 17276
rect 20692 17220 20740 17276
rect 20796 17220 20806 17276
rect 32722 17164 32732 17220
rect 32788 17164 33292 17220
rect 33348 17164 35196 17220
rect 35252 17164 35262 17220
rect 13458 17052 13468 17108
rect 13524 17052 14588 17108
rect 14644 17052 14654 17108
rect 17042 17052 17052 17108
rect 17108 17052 17612 17108
rect 17668 17052 17678 17108
rect 19282 17052 19292 17108
rect 19348 17052 20188 17108
rect 20244 17052 20254 17108
rect 29138 17052 29148 17108
rect 29204 17052 30268 17108
rect 30324 17052 30334 17108
rect 31938 17052 31948 17108
rect 32004 17052 34972 17108
rect 35028 17052 35038 17108
rect 37212 16996 37268 17276
rect 39842 17220 39852 17276
rect 39908 17220 39956 17276
rect 40012 17220 40060 17276
rect 40116 17220 40126 17276
rect 40236 17108 40292 17276
rect 40908 17220 40964 17276
rect 59162 17220 59172 17276
rect 59228 17220 59276 17276
rect 59332 17220 59380 17276
rect 59436 17220 59446 17276
rect 78482 17220 78492 17276
rect 78548 17220 78596 17276
rect 78652 17220 78700 17276
rect 78756 17220 78766 17276
rect 40908 17164 54460 17220
rect 54516 17164 55020 17220
rect 55076 17164 55086 17220
rect 60284 17164 61292 17220
rect 61348 17164 61358 17220
rect 63858 17164 63868 17220
rect 63924 17164 64652 17220
rect 64708 17164 64718 17220
rect 60284 17108 60340 17164
rect 39442 17052 39452 17108
rect 39508 17052 40292 17108
rect 40898 17052 40908 17108
rect 40964 17052 41804 17108
rect 41860 17052 41870 17108
rect 45266 17052 45276 17108
rect 45332 17052 47628 17108
rect 47684 17052 48636 17108
rect 48692 17052 48702 17108
rect 51650 17052 51660 17108
rect 51716 17052 52892 17108
rect 52948 17052 52958 17108
rect 54796 17052 60284 17108
rect 60340 17052 60350 17108
rect 60722 17052 60732 17108
rect 60788 17052 61404 17108
rect 61460 17052 61470 17108
rect 61852 17052 63084 17108
rect 63140 17052 63150 17108
rect 64418 17052 64428 17108
rect 64484 17052 64494 17108
rect 54796 16996 54852 17052
rect 61852 16996 61908 17052
rect 64428 16996 64484 17052
rect 12338 16940 12348 16996
rect 12404 16940 13580 16996
rect 13636 16940 14812 16996
rect 14868 16940 14878 16996
rect 16930 16940 16940 16996
rect 16996 16940 19068 16996
rect 19124 16940 19134 16996
rect 19842 16940 19852 16996
rect 19908 16940 21868 16996
rect 21924 16940 22204 16996
rect 22260 16940 22270 16996
rect 28018 16940 28028 16996
rect 28084 16940 28644 16996
rect 31826 16940 31836 16996
rect 31892 16940 32508 16996
rect 32564 16940 36988 16996
rect 37044 16940 37054 16996
rect 37212 16940 38668 16996
rect 42018 16940 42028 16996
rect 42084 16940 42476 16996
rect 42532 16940 46396 16996
rect 46452 16940 46462 16996
rect 47394 16940 47404 16996
rect 47460 16940 48188 16996
rect 48244 16940 49420 16996
rect 49476 16940 51884 16996
rect 51940 16940 54852 16996
rect 55010 16940 55020 16996
rect 55076 16940 61852 16996
rect 61908 16940 61918 16996
rect 62132 16940 63868 16996
rect 63924 16940 63934 16996
rect 64082 16940 64092 16996
rect 64148 16940 65772 16996
rect 65828 16940 65838 16996
rect 66434 16940 66444 16996
rect 66500 16940 67564 16996
rect 67620 16940 67630 16996
rect 28588 16884 28644 16940
rect 38612 16884 38668 16940
rect 62132 16884 62188 16940
rect 3042 16828 3052 16884
rect 3108 16828 3612 16884
rect 3668 16828 3678 16884
rect 4386 16828 4396 16884
rect 4452 16828 5292 16884
rect 5348 16828 5358 16884
rect 16146 16828 16156 16884
rect 16212 16828 16380 16884
rect 16436 16828 16828 16884
rect 16884 16828 16894 16884
rect 18274 16828 18284 16884
rect 18340 16828 21532 16884
rect 21588 16828 21980 16884
rect 22036 16828 22046 16884
rect 24770 16828 24780 16884
rect 24836 16828 25788 16884
rect 25844 16828 26124 16884
rect 26180 16828 26190 16884
rect 28588 16828 30828 16884
rect 30884 16828 32844 16884
rect 32900 16828 32910 16884
rect 35858 16828 35868 16884
rect 35924 16828 37772 16884
rect 37828 16828 37838 16884
rect 38612 16828 41804 16884
rect 41860 16828 41870 16884
rect 43810 16828 43820 16884
rect 43876 16828 50988 16884
rect 51044 16828 51054 16884
rect 53666 16828 53676 16884
rect 53732 16828 54236 16884
rect 54292 16828 54302 16884
rect 55122 16828 55132 16884
rect 55188 16828 55916 16884
rect 55972 16828 57484 16884
rect 57540 16828 57550 16884
rect 61394 16828 61404 16884
rect 61460 16828 61740 16884
rect 61796 16828 62188 16884
rect 63410 16828 63420 16884
rect 63476 16828 64428 16884
rect 64484 16828 64494 16884
rect 64754 16828 64764 16884
rect 64820 16828 66892 16884
rect 66948 16828 66958 16884
rect 67442 16828 67452 16884
rect 67508 16828 69468 16884
rect 69524 16828 69804 16884
rect 69860 16828 69870 16884
rect 76066 16828 76076 16884
rect 76132 16828 76142 16884
rect 47068 16772 47124 16828
rect 76076 16772 76132 16828
rect 3826 16716 3836 16772
rect 3892 16716 4508 16772
rect 4564 16716 4574 16772
rect 4834 16716 4844 16772
rect 4900 16716 6972 16772
rect 7028 16716 7038 16772
rect 15250 16716 15260 16772
rect 15316 16716 15708 16772
rect 15764 16716 16716 16772
rect 16772 16716 16782 16772
rect 18498 16716 18508 16772
rect 18564 16716 19404 16772
rect 19460 16716 20412 16772
rect 20468 16716 20636 16772
rect 20692 16716 20702 16772
rect 28018 16716 28028 16772
rect 28084 16716 29260 16772
rect 29316 16716 29326 16772
rect 29586 16716 29596 16772
rect 29652 16716 30156 16772
rect 30212 16716 30222 16772
rect 37874 16716 37884 16772
rect 37940 16716 42028 16772
rect 42084 16716 42094 16772
rect 44258 16716 44268 16772
rect 44324 16716 45388 16772
rect 45444 16716 45454 16772
rect 47058 16716 47068 16772
rect 47124 16716 47134 16772
rect 48962 16716 48972 16772
rect 49028 16716 49756 16772
rect 49812 16716 49822 16772
rect 50082 16716 50092 16772
rect 50148 16716 50652 16772
rect 50708 16716 50876 16772
rect 50932 16716 50942 16772
rect 51874 16716 51884 16772
rect 51940 16716 52668 16772
rect 52724 16716 52734 16772
rect 56354 16716 56364 16772
rect 56420 16716 56700 16772
rect 56756 16716 57708 16772
rect 57764 16716 57774 16772
rect 76076 16716 78260 16772
rect 29596 16660 29652 16716
rect 18610 16604 18620 16660
rect 18676 16604 19292 16660
rect 19348 16604 19358 16660
rect 28578 16604 28588 16660
rect 28644 16604 29652 16660
rect 29708 16604 32732 16660
rect 32788 16604 32798 16660
rect 40562 16604 40572 16660
rect 40628 16604 69468 16660
rect 69524 16604 69534 16660
rect 76066 16604 76076 16660
rect 76132 16604 76636 16660
rect 76692 16604 77420 16660
rect 77476 16604 77980 16660
rect 78036 16604 78046 16660
rect 29708 16548 29764 16604
rect 29698 16492 29708 16548
rect 29764 16492 29774 16548
rect 42018 16492 42028 16548
rect 42084 16492 45612 16548
rect 45668 16492 46284 16548
rect 46340 16492 46350 16548
rect 75282 16492 75292 16548
rect 75348 16492 75964 16548
rect 76020 16492 76030 16548
rect 10862 16436 10872 16492
rect 10928 16436 10976 16492
rect 11032 16436 11080 16492
rect 11136 16436 11146 16492
rect 30182 16436 30192 16492
rect 30248 16436 30296 16492
rect 30352 16436 30400 16492
rect 30456 16436 30466 16492
rect 49502 16436 49512 16492
rect 49568 16436 49616 16492
rect 49672 16436 49720 16492
rect 49776 16436 49786 16492
rect 68822 16436 68832 16492
rect 68888 16436 68936 16492
rect 68992 16436 69040 16492
rect 69096 16436 69106 16492
rect 40450 16380 40460 16436
rect 40516 16380 43932 16436
rect 43988 16380 43998 16436
rect 50372 16380 61628 16436
rect 61684 16380 62076 16436
rect 62132 16380 62636 16436
rect 62692 16380 62702 16436
rect 0 16324 800 16352
rect 50372 16324 50428 16380
rect 78204 16324 78260 16716
rect 79200 16324 80000 16352
rect 0 16268 2492 16324
rect 2548 16268 2558 16324
rect 15138 16268 15148 16324
rect 15204 16268 16268 16324
rect 16324 16268 18172 16324
rect 18228 16268 18732 16324
rect 18788 16268 18798 16324
rect 31714 16268 31724 16324
rect 31780 16268 34972 16324
rect 35028 16268 35038 16324
rect 41906 16268 41916 16324
rect 41972 16268 47628 16324
rect 47684 16268 49868 16324
rect 49924 16268 50428 16324
rect 52322 16268 52332 16324
rect 52388 16268 54236 16324
rect 54292 16268 54302 16324
rect 62290 16268 62300 16324
rect 62356 16268 62916 16324
rect 64978 16268 64988 16324
rect 65044 16268 65548 16324
rect 65604 16268 65614 16324
rect 78204 16268 80000 16324
rect 0 16240 800 16268
rect 62860 16212 62916 16268
rect 79200 16240 80000 16268
rect 4050 16156 4060 16212
rect 4116 16156 6188 16212
rect 6244 16156 7420 16212
rect 7476 16156 7486 16212
rect 13906 16156 13916 16212
rect 13972 16156 14364 16212
rect 14420 16156 16492 16212
rect 16548 16156 16558 16212
rect 17154 16156 17164 16212
rect 17220 16156 17388 16212
rect 17444 16156 18508 16212
rect 18564 16156 18574 16212
rect 18732 16156 23436 16212
rect 23492 16156 23502 16212
rect 30258 16156 30268 16212
rect 30324 16156 30828 16212
rect 30884 16156 30894 16212
rect 35410 16156 35420 16212
rect 35476 16156 35868 16212
rect 35924 16156 37212 16212
rect 37268 16156 37278 16212
rect 38444 16156 40124 16212
rect 40180 16156 40190 16212
rect 61954 16156 61964 16212
rect 62020 16156 62636 16212
rect 62692 16156 62702 16212
rect 62850 16156 62860 16212
rect 62916 16156 63644 16212
rect 63700 16156 75404 16212
rect 75460 16156 75470 16212
rect 18732 16100 18788 16156
rect 38444 16100 38500 16156
rect 6626 16044 6636 16100
rect 6692 16044 7756 16100
rect 7812 16044 11340 16100
rect 11396 16044 11406 16100
rect 11900 16044 15708 16100
rect 15764 16044 18788 16100
rect 19628 16044 21644 16100
rect 21700 16044 22316 16100
rect 22372 16044 22652 16100
rect 22708 16044 22718 16100
rect 23314 16044 23324 16100
rect 23380 16044 23772 16100
rect 23828 16044 24220 16100
rect 24276 16044 24668 16100
rect 24724 16044 24734 16100
rect 26450 16044 26460 16100
rect 26516 16044 27244 16100
rect 27300 16044 27310 16100
rect 11900 15988 11956 16044
rect 19628 15988 19684 16044
rect 9202 15932 9212 15988
rect 9268 15932 9996 15988
rect 10052 15932 11956 15988
rect 12114 15932 12124 15988
rect 12180 15932 12572 15988
rect 12628 15932 14588 15988
rect 14644 15932 14654 15988
rect 16706 15932 16716 15988
rect 16772 15932 17948 15988
rect 18004 15932 18956 15988
rect 19012 15932 19628 15988
rect 19684 15932 19694 15988
rect 20290 15932 20300 15988
rect 20356 15932 23156 15988
rect 26114 15932 26124 15988
rect 26180 15932 27132 15988
rect 27188 15932 27198 15988
rect 8978 15820 8988 15876
rect 9044 15820 9884 15876
rect 9940 15820 10444 15876
rect 10500 15820 10510 15876
rect 11218 15820 11228 15876
rect 11284 15820 11900 15876
rect 11956 15820 12348 15876
rect 12404 15820 12414 15876
rect 12898 15820 12908 15876
rect 12964 15820 13580 15876
rect 13636 15820 13646 15876
rect 15922 15820 15932 15876
rect 15988 15820 17836 15876
rect 17892 15820 17902 15876
rect 20626 15820 20636 15876
rect 20692 15820 21700 15876
rect 13580 15708 15148 15764
rect 15204 15708 15214 15764
rect 13580 15652 13636 15708
rect 20522 15652 20532 15708
rect 20588 15652 20636 15708
rect 20692 15652 20740 15708
rect 20796 15652 20806 15708
rect 12674 15596 12684 15652
rect 12740 15596 13580 15652
rect 13636 15596 13646 15652
rect 21644 15540 21700 15820
rect 23100 15540 23156 15932
rect 28914 15820 28924 15876
rect 28980 15820 29708 15876
rect 29764 15820 29774 15876
rect 31154 15820 31164 15876
rect 31220 15820 31724 15876
rect 31780 15820 31790 15876
rect 31892 15764 31948 16100
rect 32004 16044 32014 16100
rect 32162 16044 32172 16100
rect 32228 16044 32266 16100
rect 37650 16044 37660 16100
rect 37716 16044 38444 16100
rect 38500 16044 38510 16100
rect 39106 16044 39116 16100
rect 39172 16044 39900 16100
rect 39956 16044 39966 16100
rect 48514 16044 48524 16100
rect 48580 16044 49420 16100
rect 49476 16044 49486 16100
rect 53106 16044 53116 16100
rect 53172 16044 54572 16100
rect 54628 16044 55580 16100
rect 55636 16044 56644 16100
rect 56914 16044 56924 16100
rect 56980 16044 57484 16100
rect 57540 16044 57550 16100
rect 59938 16044 59948 16100
rect 60004 16044 60396 16100
rect 60452 16044 60462 16100
rect 64194 16044 64204 16100
rect 64260 16044 66220 16100
rect 66276 16044 67340 16100
rect 67396 16044 67406 16100
rect 73266 16044 73276 16100
rect 73332 16044 73948 16100
rect 74004 16044 74014 16100
rect 74834 16044 74844 16100
rect 74900 16044 75964 16100
rect 76020 16044 77084 16100
rect 77140 16044 77150 16100
rect 38444 15988 38500 16044
rect 56588 15988 56644 16044
rect 32050 15932 32060 15988
rect 32116 15932 32396 15988
rect 32452 15932 32462 15988
rect 32610 15932 32620 15988
rect 32676 15932 33516 15988
rect 33572 15932 34412 15988
rect 34468 15932 34478 15988
rect 38444 15932 39564 15988
rect 39620 15932 39630 15988
rect 54786 15932 54796 15988
rect 54852 15932 56364 15988
rect 56420 15932 56430 15988
rect 56588 15932 57372 15988
rect 57428 15932 57820 15988
rect 57876 15932 62972 15988
rect 63028 15932 64316 15988
rect 64372 15932 64382 15988
rect 76738 15932 76748 15988
rect 76804 15932 77308 15988
rect 77364 15932 77374 15988
rect 32498 15820 32508 15876
rect 32564 15820 33740 15876
rect 33796 15820 34524 15876
rect 34580 15820 34590 15876
rect 38658 15820 38668 15876
rect 38724 15820 39004 15876
rect 39060 15820 40236 15876
rect 40292 15820 40302 15876
rect 41682 15820 41692 15876
rect 41748 15820 42700 15876
rect 42756 15820 50428 15876
rect 50484 15820 50494 15876
rect 50866 15820 50876 15876
rect 50932 15820 52780 15876
rect 52836 15820 55692 15876
rect 55748 15820 57596 15876
rect 57652 15820 57662 15876
rect 61618 15820 61628 15876
rect 61684 15820 62076 15876
rect 62132 15820 64652 15876
rect 64708 15820 65884 15876
rect 65940 15820 69244 15876
rect 69300 15820 69310 15876
rect 31892 15708 32396 15764
rect 32452 15708 32462 15764
rect 34290 15708 34300 15764
rect 34356 15708 38892 15764
rect 38948 15708 38958 15764
rect 46498 15708 46508 15764
rect 46564 15708 47292 15764
rect 47348 15708 47358 15764
rect 39842 15652 39852 15708
rect 39908 15652 39956 15708
rect 40012 15652 40060 15708
rect 40116 15652 40126 15708
rect 59162 15652 59172 15708
rect 59228 15652 59276 15708
rect 59332 15652 59380 15708
rect 59436 15652 59446 15708
rect 78482 15652 78492 15708
rect 78548 15652 78596 15708
rect 78652 15652 78700 15708
rect 78756 15652 78766 15708
rect 23426 15596 23436 15652
rect 23492 15596 37772 15652
rect 37828 15596 37838 15652
rect 62290 15596 62300 15652
rect 62356 15596 63980 15652
rect 64036 15596 68908 15652
rect 68964 15596 70924 15652
rect 70980 15596 70990 15652
rect 14466 15484 14476 15540
rect 14532 15484 15148 15540
rect 15362 15484 15372 15540
rect 15428 15484 16716 15540
rect 16772 15484 16782 15540
rect 18050 15484 18060 15540
rect 18116 15484 18844 15540
rect 18900 15484 19404 15540
rect 19460 15484 21084 15540
rect 21140 15484 21150 15540
rect 21634 15484 21644 15540
rect 21700 15484 21868 15540
rect 21924 15484 22876 15540
rect 22932 15484 22942 15540
rect 23100 15484 37604 15540
rect 15092 15428 15148 15484
rect 37548 15428 37604 15484
rect 37996 15484 71036 15540
rect 71092 15484 71102 15540
rect 75394 15484 75404 15540
rect 75460 15484 76188 15540
rect 76244 15484 77420 15540
rect 77476 15484 78092 15540
rect 78148 15484 78158 15540
rect 37996 15428 38052 15484
rect 9650 15372 9660 15428
rect 9716 15372 11004 15428
rect 11060 15372 12684 15428
rect 12740 15372 12750 15428
rect 15092 15372 23324 15428
rect 23380 15372 23390 15428
rect 29922 15372 29932 15428
rect 29988 15372 31948 15428
rect 32004 15372 32014 15428
rect 37548 15372 38052 15428
rect 43362 15372 43372 15428
rect 43428 15372 44156 15428
rect 44212 15372 44222 15428
rect 50372 15372 50652 15428
rect 50708 15372 51212 15428
rect 51268 15372 51278 15428
rect 56578 15372 56588 15428
rect 56644 15372 62972 15428
rect 63028 15372 63868 15428
rect 63924 15372 63934 15428
rect 65762 15372 65772 15428
rect 65828 15372 66332 15428
rect 66388 15372 66398 15428
rect 69458 15372 69468 15428
rect 69524 15372 69916 15428
rect 69972 15372 71596 15428
rect 71652 15372 71662 15428
rect 72258 15372 72268 15428
rect 72324 15372 73500 15428
rect 73556 15372 74060 15428
rect 74116 15372 74508 15428
rect 74564 15372 74574 15428
rect 76850 15372 76860 15428
rect 76916 15372 77532 15428
rect 77588 15372 77598 15428
rect 50372 15316 50428 15372
rect 2370 15260 2380 15316
rect 2436 15260 3052 15316
rect 3108 15260 3118 15316
rect 3938 15260 3948 15316
rect 4004 15260 4844 15316
rect 4900 15260 5404 15316
rect 5460 15260 5470 15316
rect 9660 15260 14252 15316
rect 14308 15260 14318 15316
rect 17826 15260 17836 15316
rect 17892 15260 18732 15316
rect 18788 15260 19516 15316
rect 19572 15260 19582 15316
rect 21074 15260 21084 15316
rect 21140 15260 21150 15316
rect 21298 15260 21308 15316
rect 21364 15260 22876 15316
rect 22932 15260 22942 15316
rect 31826 15260 31836 15316
rect 31892 15260 37548 15316
rect 37604 15260 37614 15316
rect 38612 15260 42308 15316
rect 42466 15260 42476 15316
rect 42532 15260 43036 15316
rect 43092 15260 44044 15316
rect 44100 15260 44604 15316
rect 44660 15260 44670 15316
rect 46834 15260 46844 15316
rect 46900 15260 48412 15316
rect 48468 15260 49980 15316
rect 50036 15260 50428 15316
rect 50530 15260 50540 15316
rect 50596 15260 51660 15316
rect 51716 15260 51726 15316
rect 52434 15260 52444 15316
rect 52500 15260 53116 15316
rect 53172 15260 53182 15316
rect 54114 15260 54124 15316
rect 54180 15260 54796 15316
rect 54852 15260 54862 15316
rect 60386 15260 60396 15316
rect 60452 15260 61516 15316
rect 61572 15260 61582 15316
rect 67890 15260 67900 15316
rect 67956 15260 70028 15316
rect 70084 15260 70094 15316
rect 75170 15260 75180 15316
rect 75236 15260 76748 15316
rect 76804 15260 76814 15316
rect 9660 15204 9716 15260
rect 21084 15204 21140 15260
rect 38612 15204 38668 15260
rect 42252 15204 42308 15260
rect 46844 15204 46900 15260
rect 4498 15148 4508 15204
rect 4564 15148 7980 15204
rect 8036 15148 8046 15204
rect 8530 15148 8540 15204
rect 8596 15148 9660 15204
rect 9716 15148 9726 15204
rect 11218 15148 11228 15204
rect 11284 15148 12348 15204
rect 12404 15148 13804 15204
rect 13860 15148 13870 15204
rect 16258 15148 16268 15204
rect 16324 15148 18060 15204
rect 18116 15148 18126 15204
rect 18274 15148 18284 15204
rect 18340 15148 19740 15204
rect 19796 15148 20300 15204
rect 20356 15148 20366 15204
rect 21084 15148 22204 15204
rect 22260 15148 22428 15204
rect 22484 15148 22494 15204
rect 29586 15148 29596 15204
rect 29652 15148 30044 15204
rect 30100 15148 30716 15204
rect 30772 15148 30782 15204
rect 32134 15148 32172 15204
rect 32228 15148 32238 15204
rect 37762 15148 37772 15204
rect 37828 15148 38668 15204
rect 38882 15148 38892 15204
rect 38948 15148 40572 15204
rect 40628 15148 40638 15204
rect 42252 15148 46900 15204
rect 50754 15148 50764 15204
rect 50820 15148 55356 15204
rect 55412 15148 55422 15204
rect 63308 15148 64092 15204
rect 64148 15148 65324 15204
rect 65380 15148 65390 15204
rect 5628 15092 5684 15148
rect 63308 15092 63364 15148
rect 3602 15036 3612 15092
rect 3668 15036 4956 15092
rect 5012 15036 5022 15092
rect 5618 15036 5628 15092
rect 5684 15036 5694 15092
rect 16034 15036 16044 15092
rect 16100 15036 33852 15092
rect 33908 15036 33918 15092
rect 42018 15036 42028 15092
rect 42084 15036 55468 15092
rect 63298 15036 63308 15092
rect 63364 15036 63374 15092
rect 70354 15036 70364 15092
rect 70420 15036 76188 15092
rect 76244 15036 76254 15092
rect 55412 14980 55468 15036
rect 39778 14924 39788 14980
rect 39844 14924 44716 14980
rect 44772 14924 44782 14980
rect 55412 14924 64652 14980
rect 64708 14924 64718 14980
rect 10862 14868 10872 14924
rect 10928 14868 10976 14924
rect 11032 14868 11080 14924
rect 11136 14868 11146 14924
rect 30182 14868 30192 14924
rect 30248 14868 30296 14924
rect 30352 14868 30400 14924
rect 30456 14868 30466 14924
rect 49502 14868 49512 14924
rect 49568 14868 49616 14924
rect 49672 14868 49720 14924
rect 49776 14868 49786 14924
rect 68822 14868 68832 14924
rect 68888 14868 68936 14924
rect 68992 14868 69040 14924
rect 69096 14868 69106 14924
rect 14802 14812 14812 14868
rect 14868 14812 24668 14868
rect 24724 14812 25452 14868
rect 25508 14812 25518 14868
rect 34850 14812 34860 14868
rect 34916 14812 35756 14868
rect 35812 14812 35822 14868
rect 38612 14812 43596 14868
rect 43652 14812 43662 14868
rect 9426 14700 9436 14756
rect 9492 14700 12460 14756
rect 12516 14700 12526 14756
rect 32386 14700 32396 14756
rect 32452 14700 34412 14756
rect 34468 14700 35644 14756
rect 35700 14700 36204 14756
rect 36260 14700 36270 14756
rect 38612 14644 38668 14812
rect 41906 14700 41916 14756
rect 41972 14700 63980 14756
rect 64036 14700 64046 14756
rect 70018 14700 70028 14756
rect 70084 14700 71260 14756
rect 71316 14700 71820 14756
rect 71876 14700 71886 14756
rect 77410 14700 77420 14756
rect 77476 14700 77756 14756
rect 77812 14700 77822 14756
rect 2706 14588 2716 14644
rect 2772 14588 38668 14644
rect 40226 14588 40236 14644
rect 40292 14588 42476 14644
rect 42532 14588 43372 14644
rect 43428 14588 43438 14644
rect 48066 14588 48076 14644
rect 48132 14588 51996 14644
rect 52052 14588 52444 14644
rect 52500 14588 52510 14644
rect 57026 14588 57036 14644
rect 57092 14588 58156 14644
rect 58212 14588 58222 14644
rect 66322 14588 66332 14644
rect 66388 14588 67004 14644
rect 67060 14588 67676 14644
rect 67732 14588 67742 14644
rect 72370 14588 72380 14644
rect 72436 14588 73052 14644
rect 73108 14588 73118 14644
rect 3602 14476 3612 14532
rect 3668 14476 4620 14532
rect 4676 14476 5516 14532
rect 5572 14476 5582 14532
rect 8754 14476 8764 14532
rect 8820 14476 20692 14532
rect 20962 14476 20972 14532
rect 21028 14476 33628 14532
rect 33684 14476 33694 14532
rect 33954 14476 33964 14532
rect 34020 14476 34972 14532
rect 35028 14476 35980 14532
rect 36036 14476 36046 14532
rect 39106 14476 39116 14532
rect 39172 14476 40684 14532
rect 40740 14476 40750 14532
rect 46050 14476 46060 14532
rect 46116 14476 53116 14532
rect 53172 14476 54908 14532
rect 54964 14476 54974 14532
rect 66882 14476 66892 14532
rect 66948 14476 68012 14532
rect 68068 14476 68078 14532
rect 70466 14476 70476 14532
rect 70532 14476 71484 14532
rect 71540 14476 72044 14532
rect 72100 14476 72110 14532
rect 3938 14364 3948 14420
rect 4004 14364 7084 14420
rect 7140 14364 8092 14420
rect 8148 14364 8158 14420
rect 8642 14364 8652 14420
rect 8708 14364 9324 14420
rect 9380 14364 9390 14420
rect 12226 14364 12236 14420
rect 12292 14364 13468 14420
rect 13524 14364 14364 14420
rect 14420 14364 14430 14420
rect 14578 14364 14588 14420
rect 14644 14364 15596 14420
rect 15652 14364 15662 14420
rect 20636 14308 20692 14476
rect 26786 14364 26796 14420
rect 26852 14364 27692 14420
rect 27748 14364 28812 14420
rect 28868 14364 28878 14420
rect 39890 14364 39900 14420
rect 39956 14364 40348 14420
rect 40404 14364 40414 14420
rect 50306 14364 50316 14420
rect 50372 14364 50764 14420
rect 50820 14364 50830 14420
rect 60498 14364 60508 14420
rect 60564 14364 61292 14420
rect 61348 14364 66108 14420
rect 66164 14364 66174 14420
rect 68226 14364 68236 14420
rect 68292 14364 74620 14420
rect 74676 14364 74686 14420
rect 3378 14252 3388 14308
rect 3444 14252 3724 14308
rect 3780 14252 6076 14308
rect 6132 14252 6142 14308
rect 7186 14252 7196 14308
rect 7252 14252 9548 14308
rect 9604 14252 9614 14308
rect 9874 14252 9884 14308
rect 9940 14252 12348 14308
rect 12404 14252 12414 14308
rect 14690 14252 14700 14308
rect 14756 14252 15148 14308
rect 15204 14252 15214 14308
rect 20636 14252 27468 14308
rect 27524 14252 27534 14308
rect 28018 14252 28028 14308
rect 28084 14252 28700 14308
rect 28756 14252 28766 14308
rect 34738 14252 34748 14308
rect 34804 14252 35308 14308
rect 35364 14252 35374 14308
rect 37762 14252 37772 14308
rect 37828 14252 39788 14308
rect 39844 14252 39854 14308
rect 41570 14252 41580 14308
rect 41636 14252 42252 14308
rect 42308 14252 42318 14308
rect 48402 14252 48412 14308
rect 48468 14252 50876 14308
rect 50932 14252 50942 14308
rect 60274 14252 60284 14308
rect 60340 14252 61404 14308
rect 61460 14252 62524 14308
rect 62580 14252 62590 14308
rect 3826 14140 3836 14196
rect 3892 14140 4900 14196
rect 40674 14140 40684 14196
rect 40740 14140 45948 14196
rect 46004 14140 46284 14196
rect 46340 14140 46350 14196
rect 67106 14140 67116 14196
rect 67172 14140 67228 14196
rect 67284 14140 68236 14196
rect 68292 14140 68302 14196
rect 3154 13916 3164 13972
rect 3220 13916 3836 13972
rect 3892 13916 4508 13972
rect 4564 13916 4574 13972
rect 0 13860 800 13888
rect 0 13804 1932 13860
rect 1988 13804 1998 13860
rect 0 13776 800 13804
rect 4844 13748 4900 14140
rect 20522 14084 20532 14140
rect 20588 14084 20636 14140
rect 20692 14084 20740 14140
rect 20796 14084 20806 14140
rect 39842 14084 39852 14140
rect 39908 14084 39956 14140
rect 40012 14084 40060 14140
rect 40116 14084 40126 14140
rect 59162 14084 59172 14140
rect 59228 14084 59276 14140
rect 59332 14084 59380 14140
rect 59436 14084 59446 14140
rect 78482 14084 78492 14140
rect 78548 14084 78596 14140
rect 78652 14084 78700 14140
rect 78756 14084 78766 14140
rect 43250 14028 43260 14084
rect 43316 14028 48748 14084
rect 48804 14028 50092 14084
rect 50148 14028 50158 14084
rect 67442 14028 67452 14084
rect 67508 14028 69692 14084
rect 69748 14028 69758 14084
rect 16146 13916 16156 13972
rect 16212 13916 16828 13972
rect 16884 13916 16894 13972
rect 18946 13916 18956 13972
rect 19012 13916 23996 13972
rect 24052 13916 24062 13972
rect 24220 13916 67228 13972
rect 67284 13916 67788 13972
rect 67844 13916 67854 13972
rect 10434 13804 10444 13860
rect 10500 13804 12124 13860
rect 12180 13804 12190 13860
rect 15250 13804 15260 13860
rect 15316 13804 15708 13860
rect 15764 13804 21252 13860
rect 23090 13804 23100 13860
rect 23156 13804 23884 13860
rect 23940 13804 23950 13860
rect 17836 13748 17892 13804
rect 21196 13748 21252 13804
rect 24220 13748 24276 13916
rect 79200 13860 80000 13888
rect 25442 13804 25452 13860
rect 25508 13804 26012 13860
rect 26068 13804 26684 13860
rect 26740 13804 26750 13860
rect 30146 13804 30156 13860
rect 30212 13804 33404 13860
rect 33460 13804 33470 13860
rect 37314 13804 37324 13860
rect 37380 13804 37548 13860
rect 37604 13804 37884 13860
rect 37940 13804 38444 13860
rect 38500 13804 38510 13860
rect 45378 13804 45388 13860
rect 45444 13804 46172 13860
rect 46228 13804 46238 13860
rect 50418 13804 50428 13860
rect 50484 13804 55468 13860
rect 58146 13804 58156 13860
rect 58212 13804 59276 13860
rect 59332 13804 59342 13860
rect 60050 13804 60060 13860
rect 60116 13804 61068 13860
rect 61124 13804 61516 13860
rect 61572 13804 61582 13860
rect 64642 13804 64652 13860
rect 64708 13804 65436 13860
rect 65492 13804 65502 13860
rect 68226 13804 68236 13860
rect 68292 13804 70140 13860
rect 70196 13804 70206 13860
rect 71698 13804 71708 13860
rect 71764 13804 73500 13860
rect 73556 13804 73566 13860
rect 76066 13804 76076 13860
rect 76132 13804 80000 13860
rect 55412 13748 55468 13804
rect 79200 13776 80000 13804
rect 2594 13692 2604 13748
rect 2660 13692 3388 13748
rect 3444 13692 3454 13748
rect 4834 13692 4844 13748
rect 4900 13692 5516 13748
rect 5572 13692 6636 13748
rect 6692 13692 6702 13748
rect 8194 13692 8204 13748
rect 8260 13692 9884 13748
rect 9940 13692 9950 13748
rect 11442 13692 11452 13748
rect 11508 13692 11900 13748
rect 11956 13692 12908 13748
rect 12964 13692 12974 13748
rect 17826 13692 17836 13748
rect 17892 13692 17902 13748
rect 19058 13692 19068 13748
rect 19124 13692 20972 13748
rect 21028 13692 21038 13748
rect 21196 13692 24276 13748
rect 24994 13692 25004 13748
rect 25060 13692 25564 13748
rect 25620 13692 25630 13748
rect 27458 13692 27468 13748
rect 27524 13692 28140 13748
rect 28196 13692 28206 13748
rect 28802 13692 28812 13748
rect 28868 13692 29484 13748
rect 29540 13692 29550 13748
rect 32610 13692 32620 13748
rect 32676 13692 34860 13748
rect 34916 13692 34926 13748
rect 35298 13692 35308 13748
rect 35364 13692 36316 13748
rect 36372 13692 36382 13748
rect 39666 13692 39676 13748
rect 39732 13692 40348 13748
rect 40404 13692 40572 13748
rect 40628 13692 40638 13748
rect 55412 13692 64988 13748
rect 65044 13692 66556 13748
rect 66612 13692 69356 13748
rect 69412 13692 69422 13748
rect 71474 13692 71484 13748
rect 71540 13692 72268 13748
rect 72324 13692 72334 13748
rect 3490 13580 3500 13636
rect 3556 13580 4732 13636
rect 4788 13580 5292 13636
rect 5348 13580 5358 13636
rect 6066 13580 6076 13636
rect 6132 13580 7756 13636
rect 7812 13580 9772 13636
rect 9828 13580 9838 13636
rect 10210 13580 10220 13636
rect 10276 13580 15708 13636
rect 15764 13580 16716 13636
rect 16772 13580 16782 13636
rect 17714 13580 17724 13636
rect 17780 13580 20972 13636
rect 21028 13580 21038 13636
rect 26114 13580 26124 13636
rect 26180 13580 28028 13636
rect 28084 13580 28094 13636
rect 34066 13580 34076 13636
rect 34132 13580 34636 13636
rect 34692 13580 35756 13636
rect 35812 13580 35822 13636
rect 39890 13580 39900 13636
rect 39956 13580 40796 13636
rect 40852 13580 40862 13636
rect 45938 13580 45948 13636
rect 46004 13580 48636 13636
rect 48692 13580 49980 13636
rect 50036 13580 50046 13636
rect 66098 13580 66108 13636
rect 66164 13580 66174 13636
rect 68002 13580 68012 13636
rect 68068 13580 70364 13636
rect 70420 13580 70812 13636
rect 70868 13580 71372 13636
rect 71428 13580 71438 13636
rect 76402 13580 76412 13636
rect 76468 13580 76972 13636
rect 77028 13580 77038 13636
rect 4946 13468 4956 13524
rect 5012 13468 5628 13524
rect 5684 13468 5694 13524
rect 11666 13468 11676 13524
rect 11732 13468 13804 13524
rect 13860 13468 14140 13524
rect 14196 13468 14206 13524
rect 18162 13468 18172 13524
rect 18228 13468 19740 13524
rect 19796 13468 19806 13524
rect 32722 13468 32732 13524
rect 32788 13468 41580 13524
rect 41636 13468 41646 13524
rect 53106 13468 53116 13524
rect 53172 13468 54012 13524
rect 54068 13468 54078 13524
rect 54338 13468 54348 13524
rect 54404 13468 59836 13524
rect 59892 13468 61628 13524
rect 61684 13468 61694 13524
rect 66108 13412 66164 13580
rect 75394 13468 75404 13524
rect 75460 13468 77420 13524
rect 77476 13468 77486 13524
rect 2594 13356 2604 13412
rect 2660 13356 4620 13412
rect 4676 13356 4686 13412
rect 15092 13356 25452 13412
rect 25508 13356 25518 13412
rect 46834 13356 46844 13412
rect 46900 13356 48300 13412
rect 48356 13356 48366 13412
rect 55346 13356 55356 13412
rect 55412 13356 56924 13412
rect 56980 13356 56990 13412
rect 65538 13356 65548 13412
rect 65604 13356 66164 13412
rect 75282 13356 75292 13412
rect 75348 13356 76300 13412
rect 76356 13356 76366 13412
rect 10862 13300 10872 13356
rect 10928 13300 10976 13356
rect 11032 13300 11080 13356
rect 11136 13300 11146 13356
rect 2370 13244 2380 13300
rect 2436 13244 2828 13300
rect 2884 13244 6636 13300
rect 6692 13244 6702 13300
rect 15092 13188 15148 13356
rect 30182 13300 30192 13356
rect 30248 13300 30296 13356
rect 30352 13300 30400 13356
rect 30456 13300 30466 13356
rect 49502 13300 49512 13356
rect 49568 13300 49616 13356
rect 49672 13300 49720 13356
rect 49776 13300 49786 13356
rect 68822 13300 68832 13356
rect 68888 13300 68936 13356
rect 68992 13300 69040 13356
rect 69096 13300 69106 13356
rect 24546 13244 24556 13300
rect 24612 13244 28924 13300
rect 28980 13244 28990 13300
rect 35634 13244 35644 13300
rect 35700 13244 44100 13300
rect 54450 13244 54460 13300
rect 54516 13244 55356 13300
rect 55412 13244 55422 13300
rect 44044 13188 44100 13244
rect 7858 13132 7868 13188
rect 7924 13132 15148 13188
rect 16706 13132 16716 13188
rect 16772 13132 28476 13188
rect 28532 13132 28542 13188
rect 30706 13132 30716 13188
rect 30772 13132 43988 13188
rect 44044 13132 55916 13188
rect 55972 13132 55982 13188
rect 65538 13132 65548 13188
rect 65604 13132 65614 13188
rect 66994 13132 67004 13188
rect 67060 13132 69804 13188
rect 69860 13132 70252 13188
rect 70308 13132 70318 13188
rect 75506 13132 75516 13188
rect 75572 13132 77308 13188
rect 77364 13132 77374 13188
rect 43932 13076 43988 13132
rect 65548 13076 65604 13132
rect 12338 13020 12348 13076
rect 12404 13020 13356 13076
rect 13412 13020 13422 13076
rect 13682 13020 13692 13076
rect 13748 13020 14364 13076
rect 14420 13020 14430 13076
rect 18134 13020 18172 13076
rect 18228 13020 18238 13076
rect 18834 13020 18844 13076
rect 18900 13020 19292 13076
rect 19348 13020 19358 13076
rect 26852 13020 42028 13076
rect 42084 13020 42094 13076
rect 43932 13020 44100 13076
rect 50978 13020 50988 13076
rect 51044 13020 57148 13076
rect 57204 13020 58044 13076
rect 58100 13020 58110 13076
rect 59164 13020 60620 13076
rect 60676 13020 64428 13076
rect 64484 13020 65604 13076
rect 67218 13020 67228 13076
rect 67284 13020 68124 13076
rect 68180 13020 68190 13076
rect 13692 12852 13748 13020
rect 26852 12964 26908 13020
rect 15922 12908 15932 12964
rect 15988 12908 18396 12964
rect 18452 12908 19404 12964
rect 19460 12908 21700 12964
rect 22978 12908 22988 12964
rect 23044 12908 26908 12964
rect 40786 12908 40796 12964
rect 40852 12908 42476 12964
rect 42532 12908 43596 12964
rect 43652 12908 43662 12964
rect 21644 12852 21700 12908
rect 4162 12796 4172 12852
rect 4228 12796 4844 12852
rect 4900 12796 4910 12852
rect 12338 12796 12348 12852
rect 12404 12796 13020 12852
rect 13076 12796 13748 12852
rect 17938 12796 17948 12852
rect 18004 12796 18508 12852
rect 18564 12796 18574 12852
rect 18722 12796 18732 12852
rect 18788 12796 19180 12852
rect 19236 12796 20300 12852
rect 20356 12796 20366 12852
rect 21634 12796 21644 12852
rect 21700 12796 22092 12852
rect 22148 12796 29260 12852
rect 29316 12796 29326 12852
rect 35970 12796 35980 12852
rect 36036 12796 36540 12852
rect 36596 12796 37884 12852
rect 37940 12796 37950 12852
rect 7186 12684 7196 12740
rect 7252 12684 7756 12740
rect 7812 12684 8540 12740
rect 8596 12684 8606 12740
rect 19282 12684 19292 12740
rect 19348 12684 19964 12740
rect 20020 12684 20030 12740
rect 20178 12684 20188 12740
rect 20244 12684 25004 12740
rect 25060 12684 25070 12740
rect 27346 12684 27356 12740
rect 27412 12684 28028 12740
rect 28084 12684 29596 12740
rect 29652 12684 30044 12740
rect 30100 12684 30268 12740
rect 30324 12684 30334 12740
rect 31490 12684 31500 12740
rect 31556 12684 32172 12740
rect 32228 12684 34076 12740
rect 34132 12684 34142 12740
rect 35522 12684 35532 12740
rect 35588 12684 36652 12740
rect 36708 12684 37212 12740
rect 37268 12684 37772 12740
rect 37828 12684 37838 12740
rect 44044 12628 44100 13020
rect 44930 12908 44940 12964
rect 44996 12908 45836 12964
rect 45892 12908 45902 12964
rect 49634 12908 49644 12964
rect 49700 12908 50876 12964
rect 50932 12908 50942 12964
rect 53778 12908 53788 12964
rect 53844 12908 55132 12964
rect 55188 12908 56140 12964
rect 56196 12908 56206 12964
rect 59164 12852 59220 13020
rect 60162 12908 60172 12964
rect 60228 12908 61292 12964
rect 61348 12908 61358 12964
rect 66770 12908 66780 12964
rect 66836 12908 67900 12964
rect 67956 12908 67966 12964
rect 76066 12908 76076 12964
rect 76132 12908 77420 12964
rect 77476 12908 77486 12964
rect 44482 12796 44492 12852
rect 44548 12796 46060 12852
rect 46116 12796 46126 12852
rect 50082 12796 50092 12852
rect 50148 12796 51100 12852
rect 51156 12796 51166 12852
rect 51314 12796 51324 12852
rect 51380 12796 59220 12852
rect 59378 12796 59388 12852
rect 59444 12796 59948 12852
rect 60004 12796 61740 12852
rect 61796 12796 61806 12852
rect 70130 12796 70140 12852
rect 70196 12796 72380 12852
rect 72436 12796 72446 12852
rect 44258 12684 44268 12740
rect 44324 12684 45612 12740
rect 45668 12684 45678 12740
rect 48850 12684 48860 12740
rect 48916 12684 50652 12740
rect 50708 12684 50718 12740
rect 53666 12684 53676 12740
rect 53732 12684 61964 12740
rect 62020 12684 62412 12740
rect 62468 12684 62972 12740
rect 63028 12684 63038 12740
rect 65314 12684 65324 12740
rect 65380 12684 66220 12740
rect 66276 12684 66668 12740
rect 66724 12684 66734 12740
rect 70466 12684 70476 12740
rect 70532 12684 71148 12740
rect 71204 12684 71214 12740
rect 32834 12572 32844 12628
rect 32900 12572 37100 12628
rect 37156 12572 37166 12628
rect 44044 12572 57372 12628
rect 57428 12572 58044 12628
rect 58100 12572 58492 12628
rect 58548 12572 58558 12628
rect 63074 12572 63084 12628
rect 63140 12572 65996 12628
rect 66052 12572 66556 12628
rect 66612 12572 66622 12628
rect 20522 12516 20532 12572
rect 20588 12516 20636 12572
rect 20692 12516 20740 12572
rect 20796 12516 20806 12572
rect 39842 12516 39852 12572
rect 39908 12516 39956 12572
rect 40012 12516 40060 12572
rect 40116 12516 40126 12572
rect 59162 12516 59172 12572
rect 59228 12516 59276 12572
rect 59332 12516 59380 12572
rect 59436 12516 59446 12572
rect 78482 12516 78492 12572
rect 78548 12516 78596 12572
rect 78652 12516 78700 12572
rect 78756 12516 78766 12572
rect 8866 12460 8876 12516
rect 8932 12460 17724 12516
rect 17780 12460 17790 12516
rect 40338 12460 40348 12516
rect 40404 12460 52668 12516
rect 52724 12460 53788 12516
rect 53844 12460 53854 12516
rect 62402 12460 62412 12516
rect 62468 12460 66780 12516
rect 66836 12460 66846 12516
rect 16146 12348 16156 12404
rect 16212 12348 17052 12404
rect 17108 12348 18284 12404
rect 18340 12348 19068 12404
rect 19124 12348 19134 12404
rect 19282 12348 19292 12404
rect 19348 12348 20860 12404
rect 20916 12348 20926 12404
rect 21074 12348 21084 12404
rect 21140 12348 21980 12404
rect 22036 12348 22204 12404
rect 22260 12348 23324 12404
rect 23380 12348 55468 12404
rect 55906 12348 55916 12404
rect 55972 12348 56588 12404
rect 56644 12348 67004 12404
rect 67060 12348 67070 12404
rect 68226 12348 68236 12404
rect 68292 12348 73500 12404
rect 73556 12348 74060 12404
rect 74116 12348 74126 12404
rect 4946 12236 4956 12292
rect 5012 12236 5852 12292
rect 5908 12236 8092 12292
rect 8148 12236 8158 12292
rect 11778 12236 11788 12292
rect 11844 12236 12460 12292
rect 12516 12236 12796 12292
rect 12852 12236 14476 12292
rect 14532 12236 14542 12292
rect 15092 12236 30660 12292
rect 30818 12236 30828 12292
rect 30884 12236 33180 12292
rect 33236 12236 33246 12292
rect 34738 12236 34748 12292
rect 34804 12236 40460 12292
rect 40516 12236 40526 12292
rect 45378 12236 45388 12292
rect 45444 12236 48636 12292
rect 48692 12236 49756 12292
rect 49812 12236 49822 12292
rect 50866 12236 50876 12292
rect 50932 12236 53564 12292
rect 53620 12236 53630 12292
rect 54450 12236 54460 12292
rect 54516 12236 55244 12292
rect 55300 12236 55310 12292
rect 8978 12124 8988 12180
rect 9044 12124 10108 12180
rect 10164 12124 10174 12180
rect 12674 12124 12684 12180
rect 12740 12124 13804 12180
rect 13860 12124 13870 12180
rect 15092 12068 15148 12236
rect 30604 12180 30660 12236
rect 55412 12180 55468 12348
rect 66780 12292 66836 12348
rect 57474 12236 57484 12292
rect 57540 12236 62076 12292
rect 62132 12236 62524 12292
rect 62580 12236 62590 12292
rect 63410 12236 63420 12292
rect 63476 12236 63868 12292
rect 63924 12236 63934 12292
rect 66770 12236 66780 12292
rect 66836 12236 66846 12292
rect 68114 12236 68124 12292
rect 68180 12236 68796 12292
rect 68852 12236 69244 12292
rect 69300 12236 76748 12292
rect 76804 12236 76814 12292
rect 16146 12124 16156 12180
rect 16212 12124 16492 12180
rect 16548 12124 18172 12180
rect 18228 12124 18238 12180
rect 18722 12124 18732 12180
rect 18788 12124 19964 12180
rect 20020 12124 20524 12180
rect 20580 12124 20590 12180
rect 20850 12124 20860 12180
rect 20916 12124 24668 12180
rect 24724 12124 25228 12180
rect 25284 12124 25294 12180
rect 26786 12124 26796 12180
rect 26852 12124 27916 12180
rect 27972 12124 28588 12180
rect 28644 12124 29708 12180
rect 29764 12124 29774 12180
rect 30604 12124 31500 12180
rect 31556 12124 31566 12180
rect 31724 12124 38668 12180
rect 43586 12124 43596 12180
rect 43652 12124 43932 12180
rect 43988 12124 51324 12180
rect 51380 12124 51390 12180
rect 55412 12124 61964 12180
rect 62020 12124 62860 12180
rect 62916 12124 65436 12180
rect 65492 12124 65502 12180
rect 76178 12124 76188 12180
rect 76244 12124 77868 12180
rect 77924 12124 77934 12180
rect 9874 12012 9884 12068
rect 9940 12012 15148 12068
rect 20524 12068 20580 12124
rect 31724 12068 31780 12124
rect 20524 12012 21308 12068
rect 21364 12012 21532 12068
rect 21588 12012 21598 12068
rect 28354 12012 28364 12068
rect 28420 12012 31780 12068
rect 33394 12012 33404 12068
rect 33460 12012 35980 12068
rect 36036 12012 36046 12068
rect 6178 11900 6188 11956
rect 6244 11900 7532 11956
rect 7588 11900 7598 11956
rect 10770 11900 10780 11956
rect 10836 11900 12908 11956
rect 12964 11900 12974 11956
rect 18946 11900 18956 11956
rect 19012 11900 20076 11956
rect 20132 11900 20524 11956
rect 20580 11900 20590 11956
rect 20738 11900 20748 11956
rect 20804 11900 21084 11956
rect 21140 11900 21150 11956
rect 29698 11900 29708 11956
rect 29764 11900 35532 11956
rect 35588 11900 35598 11956
rect 38612 11844 38668 12124
rect 40114 12012 40124 12068
rect 40180 12012 42588 12068
rect 42644 12012 43596 12068
rect 43652 12012 43662 12068
rect 48402 12012 48412 12068
rect 48468 12012 49868 12068
rect 49924 12012 49934 12068
rect 56466 12012 56476 12068
rect 56532 12012 56924 12068
rect 56980 12012 65548 12068
rect 65604 12012 65614 12068
rect 69570 12012 69580 12068
rect 69636 12012 70028 12068
rect 70084 12012 70364 12068
rect 70420 12012 70430 12068
rect 59714 11900 59724 11956
rect 59780 11900 60956 11956
rect 61012 11900 61022 11956
rect 63532 11900 63756 11956
rect 63812 11900 63822 11956
rect 66770 11900 66780 11956
rect 66836 11900 67004 11956
rect 67060 11900 67452 11956
rect 67508 11900 67518 11956
rect 72370 11900 72380 11956
rect 72436 11900 76188 11956
rect 76244 11900 76254 11956
rect 63532 11844 63588 11900
rect 15362 11788 15372 11844
rect 15428 11788 24892 11844
rect 24948 11788 26012 11844
rect 26068 11788 26684 11844
rect 26740 11788 26750 11844
rect 38612 11788 48188 11844
rect 48244 11788 48254 11844
rect 63522 11788 63532 11844
rect 63588 11788 63598 11844
rect 10862 11732 10872 11788
rect 10928 11732 10976 11788
rect 11032 11732 11080 11788
rect 11136 11732 11146 11788
rect 30182 11732 30192 11788
rect 30248 11732 30296 11788
rect 30352 11732 30400 11788
rect 30456 11732 30466 11788
rect 49502 11732 49512 11788
rect 49568 11732 49616 11788
rect 49672 11732 49720 11788
rect 49776 11732 49786 11788
rect 68822 11732 68832 11788
rect 68888 11732 68936 11788
rect 68992 11732 69040 11788
rect 69096 11732 69106 11788
rect 2034 11676 2044 11732
rect 2100 11676 3164 11732
rect 3220 11676 4396 11732
rect 4452 11676 4462 11732
rect 8866 11676 8876 11732
rect 8932 11676 9996 11732
rect 10052 11676 10062 11732
rect 21970 11676 21980 11732
rect 22036 11676 22876 11732
rect 22932 11676 22942 11732
rect 35410 11676 35420 11732
rect 35476 11676 43596 11732
rect 43652 11676 43662 11732
rect 19282 11564 19292 11620
rect 19348 11564 27580 11620
rect 27636 11564 27646 11620
rect 35522 11564 35532 11620
rect 35588 11564 36204 11620
rect 36260 11564 43932 11620
rect 43988 11564 43998 11620
rect 2818 11452 2828 11508
rect 2884 11452 3276 11508
rect 3332 11452 5852 11508
rect 5908 11452 5918 11508
rect 18610 11452 18620 11508
rect 18676 11452 21644 11508
rect 21700 11452 21710 11508
rect 24322 11452 24332 11508
rect 24388 11452 25004 11508
rect 25060 11452 25676 11508
rect 25732 11452 25742 11508
rect 34290 11452 34300 11508
rect 34356 11452 41916 11508
rect 41972 11452 41982 11508
rect 54226 11452 54236 11508
rect 54292 11452 56364 11508
rect 56420 11452 56430 11508
rect 57250 11452 57260 11508
rect 57316 11452 57932 11508
rect 57988 11452 57998 11508
rect 62290 11452 62300 11508
rect 62356 11452 63308 11508
rect 63364 11452 63374 11508
rect 63746 11452 63756 11508
rect 63812 11452 66668 11508
rect 66724 11452 66734 11508
rect 75506 11452 75516 11508
rect 75572 11452 76356 11508
rect 76514 11452 76524 11508
rect 76580 11452 77532 11508
rect 77588 11452 77598 11508
rect 0 11396 800 11424
rect 76300 11396 76356 11452
rect 79200 11396 80000 11424
rect 0 11340 1932 11396
rect 1988 11340 1998 11396
rect 4162 11340 4172 11396
rect 4228 11340 5740 11396
rect 5796 11340 5806 11396
rect 8754 11340 8764 11396
rect 8820 11340 14252 11396
rect 14308 11340 14318 11396
rect 15250 11340 15260 11396
rect 15316 11340 15484 11396
rect 15540 11340 16156 11396
rect 16212 11340 16222 11396
rect 22194 11340 22204 11396
rect 22260 11340 24892 11396
rect 24948 11340 24958 11396
rect 25778 11340 25788 11396
rect 25844 11340 26908 11396
rect 26964 11340 26974 11396
rect 27906 11340 27916 11396
rect 27972 11340 29596 11396
rect 29652 11340 29662 11396
rect 46946 11340 46956 11396
rect 47012 11340 48860 11396
rect 48916 11340 51548 11396
rect 51604 11340 51614 11396
rect 57026 11340 57036 11396
rect 57092 11340 58268 11396
rect 58324 11340 58334 11396
rect 70130 11340 70140 11396
rect 70196 11340 70812 11396
rect 70868 11340 73388 11396
rect 73444 11340 73836 11396
rect 73892 11340 73902 11396
rect 74946 11340 74956 11396
rect 75012 11340 75628 11396
rect 75684 11340 75694 11396
rect 76300 11340 80000 11396
rect 0 11312 800 11340
rect 15586 11228 15596 11284
rect 15652 11228 16716 11284
rect 16772 11228 17724 11284
rect 17780 11228 19068 11284
rect 19124 11228 19134 11284
rect 24892 11172 24948 11340
rect 79200 11312 80000 11340
rect 48738 11228 48748 11284
rect 48804 11228 58940 11284
rect 58996 11228 59500 11284
rect 59556 11228 60508 11284
rect 60564 11228 60574 11284
rect 76962 11228 76972 11284
rect 77028 11228 77196 11284
rect 77252 11228 77644 11284
rect 77700 11228 77710 11284
rect 4610 11116 4620 11172
rect 4676 11116 8876 11172
rect 8932 11116 8942 11172
rect 15138 11116 15148 11172
rect 15204 11116 15708 11172
rect 15764 11116 15774 11172
rect 17266 11116 17276 11172
rect 17332 11116 17836 11172
rect 17892 11116 17902 11172
rect 24892 11116 25788 11172
rect 25844 11116 25854 11172
rect 34962 11116 34972 11172
rect 35028 11116 35644 11172
rect 35700 11116 35710 11172
rect 38546 11116 38556 11172
rect 38612 11116 39116 11172
rect 39172 11116 39788 11172
rect 39844 11116 39854 11172
rect 43586 11116 43596 11172
rect 43652 11116 44268 11172
rect 44324 11116 44334 11172
rect 50978 11116 50988 11172
rect 51044 11116 51996 11172
rect 52052 11116 52220 11172
rect 52276 11116 52286 11172
rect 55412 11116 63868 11172
rect 63924 11116 64764 11172
rect 64820 11116 64830 11172
rect 66546 11116 66556 11172
rect 66612 11116 67452 11172
rect 67508 11116 67518 11172
rect 74722 11116 74732 11172
rect 74788 11116 75852 11172
rect 75908 11116 75918 11172
rect 29922 11004 29932 11060
rect 29988 11004 36092 11060
rect 36148 11004 36158 11060
rect 20522 10948 20532 11004
rect 20588 10948 20636 11004
rect 20692 10948 20740 11004
rect 20796 10948 20806 11004
rect 39842 10948 39852 11004
rect 39908 10948 39956 11004
rect 40012 10948 40060 11004
rect 40116 10948 40126 11004
rect 55412 10948 55468 11116
rect 69346 11004 69356 11060
rect 69412 11004 70140 11060
rect 70196 11004 71036 11060
rect 71092 11004 72268 11060
rect 72324 11004 72334 11060
rect 59162 10948 59172 11004
rect 59228 10948 59276 11004
rect 59332 10948 59380 11004
rect 59436 10948 59446 11004
rect 78482 10948 78492 11004
rect 78548 10948 78596 11004
rect 78652 10948 78700 11004
rect 78756 10948 78766 11004
rect 12898 10892 12908 10948
rect 12964 10892 20356 10948
rect 52770 10892 52780 10948
rect 52836 10892 55468 10948
rect 63298 10892 63308 10948
rect 63364 10892 63532 10948
rect 63588 10892 63598 10948
rect 20300 10836 20356 10892
rect 12786 10780 12796 10836
rect 12852 10780 13244 10836
rect 13300 10780 14364 10836
rect 14420 10780 14430 10836
rect 14914 10780 14924 10836
rect 14980 10780 15932 10836
rect 15988 10780 15998 10836
rect 20300 10780 28140 10836
rect 28196 10780 28812 10836
rect 28868 10780 29820 10836
rect 29876 10780 29886 10836
rect 30818 10780 30828 10836
rect 30884 10780 31052 10836
rect 31108 10780 31836 10836
rect 31892 10780 55804 10836
rect 55860 10780 56476 10836
rect 56532 10780 56542 10836
rect 57698 10780 57708 10836
rect 57764 10780 62188 10836
rect 62244 10780 63196 10836
rect 63252 10780 63262 10836
rect 69346 10780 69356 10836
rect 69412 10780 74732 10836
rect 74788 10780 74798 10836
rect 14924 10724 14980 10780
rect 2594 10668 2604 10724
rect 2660 10668 7700 10724
rect 7858 10668 7868 10724
rect 7924 10668 8652 10724
rect 8708 10668 8718 10724
rect 12450 10668 12460 10724
rect 12516 10668 12684 10724
rect 12740 10668 14980 10724
rect 18162 10668 18172 10724
rect 18228 10668 19628 10724
rect 19684 10668 19694 10724
rect 21522 10668 21532 10724
rect 21588 10668 22316 10724
rect 22372 10668 22382 10724
rect 28466 10668 28476 10724
rect 28532 10668 32284 10724
rect 32340 10668 34972 10724
rect 35028 10668 35038 10724
rect 42242 10668 42252 10724
rect 42308 10668 47124 10724
rect 47282 10668 47292 10724
rect 47348 10668 47516 10724
rect 47572 10668 48636 10724
rect 48692 10668 49644 10724
rect 49700 10668 49710 10724
rect 52434 10668 52444 10724
rect 52500 10668 53228 10724
rect 53284 10668 53294 10724
rect 75730 10668 75740 10724
rect 75796 10668 76412 10724
rect 76468 10668 76478 10724
rect 77522 10668 77532 10724
rect 77588 10668 77980 10724
rect 78036 10668 78046 10724
rect 7644 10612 7700 10668
rect 47068 10612 47124 10668
rect 4386 10556 4396 10612
rect 4452 10556 6076 10612
rect 6132 10556 6142 10612
rect 7644 10556 7980 10612
rect 8036 10556 8046 10612
rect 11218 10556 11228 10612
rect 11284 10556 31276 10612
rect 31332 10556 31342 10612
rect 32386 10556 32396 10612
rect 32452 10556 35420 10612
rect 35476 10556 35486 10612
rect 35644 10556 40124 10612
rect 40180 10556 40572 10612
rect 40628 10556 40638 10612
rect 40786 10556 40796 10612
rect 40852 10556 43820 10612
rect 43876 10556 45276 10612
rect 45332 10556 45342 10612
rect 47068 10556 54236 10612
rect 54292 10556 54796 10612
rect 54852 10556 54862 10612
rect 56578 10556 56588 10612
rect 56644 10556 57484 10612
rect 57540 10556 57550 10612
rect 61506 10556 61516 10612
rect 61572 10556 62188 10612
rect 62244 10556 62254 10612
rect 67330 10556 67340 10612
rect 67396 10556 68572 10612
rect 68628 10556 68638 10612
rect 73714 10556 73724 10612
rect 73780 10556 74844 10612
rect 74900 10556 74910 10612
rect 76514 10556 76524 10612
rect 76580 10556 78092 10612
rect 78148 10556 78158 10612
rect 35644 10500 35700 10556
rect 40572 10500 40628 10556
rect 12002 10444 12012 10500
rect 12068 10444 12572 10500
rect 12628 10444 12908 10500
rect 12964 10444 13468 10500
rect 13524 10444 13534 10500
rect 14354 10444 14364 10500
rect 14420 10444 15148 10500
rect 15204 10444 15214 10500
rect 19058 10444 19068 10500
rect 19124 10444 27020 10500
rect 27076 10444 27086 10500
rect 29810 10444 29820 10500
rect 29876 10444 32844 10500
rect 32900 10444 32910 10500
rect 33170 10444 33180 10500
rect 33236 10444 33964 10500
rect 34020 10444 34030 10500
rect 34178 10444 34188 10500
rect 34244 10444 35700 10500
rect 36306 10444 36316 10500
rect 36372 10444 38668 10500
rect 38724 10444 38734 10500
rect 39218 10444 39228 10500
rect 39284 10444 40012 10500
rect 40068 10444 40078 10500
rect 40572 10444 41468 10500
rect 41524 10444 41534 10500
rect 44034 10444 44044 10500
rect 44100 10444 45500 10500
rect 45556 10444 45566 10500
rect 50306 10444 50316 10500
rect 50372 10444 50764 10500
rect 50820 10444 50830 10500
rect 56690 10444 56700 10500
rect 56756 10444 58380 10500
rect 58436 10444 67004 10500
rect 67060 10444 68348 10500
rect 68404 10444 68414 10500
rect 72482 10444 72492 10500
rect 72548 10444 73388 10500
rect 73444 10444 74956 10500
rect 75012 10444 75022 10500
rect 75618 10444 75628 10500
rect 75684 10444 76300 10500
rect 76356 10444 76366 10500
rect 14924 10388 14980 10444
rect 1922 10332 1932 10388
rect 1988 10332 3500 10388
rect 3556 10332 5740 10388
rect 5796 10332 5806 10388
rect 14914 10332 14924 10388
rect 14980 10332 14990 10388
rect 15092 10332 15484 10388
rect 15540 10332 15550 10388
rect 16594 10332 16604 10388
rect 16660 10332 18732 10388
rect 18788 10332 19404 10388
rect 19460 10332 19470 10388
rect 26786 10332 26796 10388
rect 26852 10332 33404 10388
rect 33460 10332 33470 10388
rect 35746 10332 35756 10388
rect 35812 10332 42476 10388
rect 42532 10332 42542 10388
rect 42802 10332 42812 10388
rect 42868 10332 50988 10388
rect 51044 10332 51054 10388
rect 67554 10332 67564 10388
rect 67620 10332 68236 10388
rect 68292 10332 68302 10388
rect 68562 10332 68572 10388
rect 68628 10332 69244 10388
rect 69300 10332 69310 10388
rect 74498 10332 74508 10388
rect 74564 10332 77980 10388
rect 78036 10332 78046 10388
rect 13234 10220 13244 10276
rect 13300 10220 14252 10276
rect 14308 10220 14318 10276
rect 10862 10164 10872 10220
rect 10928 10164 10976 10220
rect 11032 10164 11080 10220
rect 11136 10164 11146 10220
rect 15092 10164 15148 10332
rect 17154 10220 17164 10276
rect 17220 10220 19516 10276
rect 19572 10220 20300 10276
rect 20356 10220 20366 10276
rect 32946 10220 32956 10276
rect 33012 10220 39116 10276
rect 39172 10220 39182 10276
rect 50754 10220 50764 10276
rect 50820 10220 64652 10276
rect 64708 10220 65996 10276
rect 66052 10220 67340 10276
rect 67396 10220 67406 10276
rect 30182 10164 30192 10220
rect 30248 10164 30296 10220
rect 30352 10164 30400 10220
rect 30456 10164 30466 10220
rect 49502 10164 49512 10220
rect 49568 10164 49616 10220
rect 49672 10164 49720 10220
rect 49776 10164 49786 10220
rect 68822 10164 68832 10220
rect 68888 10164 68936 10220
rect 68992 10164 69040 10220
rect 69096 10164 69106 10220
rect 4722 10108 4732 10164
rect 4788 10108 7420 10164
rect 7476 10108 8652 10164
rect 8708 10108 8718 10164
rect 8978 10108 8988 10164
rect 9044 10108 10220 10164
rect 10276 10108 10286 10164
rect 13682 10108 13692 10164
rect 13748 10108 14700 10164
rect 14756 10108 15148 10164
rect 15362 10108 15372 10164
rect 15428 10108 15438 10164
rect 17938 10108 17948 10164
rect 18004 10108 25116 10164
rect 25172 10108 25182 10164
rect 39890 10108 39900 10164
rect 39956 10108 40460 10164
rect 40516 10108 40526 10164
rect 15372 10052 15428 10108
rect 6402 9996 6412 10052
rect 6468 9996 7644 10052
rect 7700 9996 7710 10052
rect 15092 9996 15428 10052
rect 17042 9996 17052 10052
rect 17108 9996 18172 10052
rect 18228 9996 18238 10052
rect 18386 9996 18396 10052
rect 18452 9996 19516 10052
rect 19572 9996 20188 10052
rect 20244 9996 20254 10052
rect 21186 9996 21196 10052
rect 21252 9996 21644 10052
rect 21700 9996 24220 10052
rect 24276 9996 24286 10052
rect 35634 9996 35644 10052
rect 35700 9996 61628 10052
rect 61684 9996 61694 10052
rect 61954 9996 61964 10052
rect 62020 9996 63420 10052
rect 63476 9996 63486 10052
rect 64530 9996 64540 10052
rect 64596 9996 66668 10052
rect 66724 9996 66734 10052
rect 4946 9884 4956 9940
rect 5012 9884 7868 9940
rect 7924 9884 7934 9940
rect 8194 9884 8204 9940
rect 8260 9884 10444 9940
rect 10500 9884 11004 9940
rect 11060 9884 11070 9940
rect 12562 9884 12572 9940
rect 12628 9884 13356 9940
rect 13412 9884 15036 9940
rect 15092 9884 15148 9996
rect 17378 9884 17388 9940
rect 17444 9884 18844 9940
rect 18900 9884 22092 9940
rect 22148 9884 22158 9940
rect 22306 9884 22316 9940
rect 22372 9884 22988 9940
rect 23044 9884 23054 9940
rect 27010 9884 27020 9940
rect 27076 9884 27804 9940
rect 27860 9884 28812 9940
rect 28868 9884 30268 9940
rect 30324 9884 30334 9940
rect 30930 9884 30940 9940
rect 30996 9884 32844 9940
rect 32900 9884 32910 9940
rect 38612 9884 61516 9940
rect 61572 9884 61582 9940
rect 61842 9884 61852 9940
rect 61908 9884 65548 9940
rect 65604 9884 66444 9940
rect 66500 9884 66510 9940
rect 74946 9884 74956 9940
rect 75012 9884 78316 9940
rect 78372 9884 78382 9940
rect 38612 9828 38668 9884
rect 2482 9772 2492 9828
rect 2548 9772 5516 9828
rect 5572 9772 7084 9828
rect 7140 9772 7150 9828
rect 7970 9772 7980 9828
rect 8036 9772 8876 9828
rect 8932 9772 8942 9828
rect 11666 9772 11676 9828
rect 11732 9772 25004 9828
rect 25060 9772 25452 9828
rect 25508 9772 26124 9828
rect 26180 9772 26190 9828
rect 28242 9772 28252 9828
rect 28308 9772 28476 9828
rect 28532 9772 38668 9828
rect 40562 9772 40572 9828
rect 40628 9772 41356 9828
rect 41412 9772 41422 9828
rect 44706 9772 44716 9828
rect 44772 9772 45724 9828
rect 45780 9772 45790 9828
rect 50978 9772 50988 9828
rect 51044 9772 51548 9828
rect 51604 9772 52108 9828
rect 52164 9772 52174 9828
rect 69682 9772 69692 9828
rect 69748 9772 70588 9828
rect 70644 9772 72156 9828
rect 72212 9772 72222 9828
rect 8876 9716 8932 9772
rect 8876 9660 15260 9716
rect 15316 9660 15326 9716
rect 15484 9660 34748 9716
rect 34804 9660 34972 9716
rect 35028 9660 35756 9716
rect 35812 9660 36540 9716
rect 36596 9660 36606 9716
rect 44594 9660 44604 9716
rect 44660 9660 45948 9716
rect 46004 9660 46014 9716
rect 50530 9660 50540 9716
rect 50596 9660 52780 9716
rect 52836 9660 52846 9716
rect 55412 9660 59948 9716
rect 60004 9660 60014 9716
rect 62402 9660 62412 9716
rect 62468 9660 63420 9716
rect 63476 9660 63486 9716
rect 69010 9660 69020 9716
rect 69076 9660 70028 9716
rect 70084 9660 71148 9716
rect 71204 9660 73724 9716
rect 73780 9660 73790 9716
rect 1922 9548 1932 9604
rect 1988 9548 4508 9604
rect 4564 9548 4574 9604
rect 5842 9548 5852 9604
rect 5908 9548 6412 9604
rect 6468 9548 6860 9604
rect 6916 9548 6926 9604
rect 13794 9548 13804 9604
rect 13860 9548 14476 9604
rect 14532 9548 15260 9604
rect 15316 9548 15326 9604
rect 10546 9436 10556 9492
rect 10612 9436 14588 9492
rect 14644 9436 15148 9492
rect 15204 9436 15214 9492
rect 15484 9380 15540 9660
rect 55412 9604 55468 9660
rect 15922 9548 15932 9604
rect 15988 9548 16268 9604
rect 16324 9548 17276 9604
rect 17332 9548 21028 9604
rect 22642 9548 22652 9604
rect 22708 9548 22988 9604
rect 23044 9548 24444 9604
rect 24500 9548 24510 9604
rect 37202 9548 37212 9604
rect 37268 9548 37436 9604
rect 37492 9548 37502 9604
rect 38210 9548 38220 9604
rect 38276 9548 38668 9604
rect 38724 9548 38734 9604
rect 40002 9548 40012 9604
rect 40068 9548 40348 9604
rect 40404 9548 40414 9604
rect 42130 9548 42140 9604
rect 42196 9548 42364 9604
rect 42420 9548 42430 9604
rect 42690 9548 42700 9604
rect 42756 9548 43260 9604
rect 43316 9548 43326 9604
rect 45378 9548 45388 9604
rect 45444 9548 50988 9604
rect 51044 9548 51054 9604
rect 54450 9548 54460 9604
rect 54516 9548 55468 9604
rect 57362 9548 57372 9604
rect 57428 9548 58492 9604
rect 58548 9548 67228 9604
rect 20972 9492 21028 9548
rect 67172 9492 67228 9548
rect 16706 9436 16716 9492
rect 16772 9436 17388 9492
rect 17444 9436 18396 9492
rect 18452 9436 18462 9492
rect 20972 9436 24052 9492
rect 24210 9436 24220 9492
rect 24276 9436 36428 9492
rect 36484 9436 37884 9492
rect 37940 9436 37950 9492
rect 43474 9436 43484 9492
rect 43540 9436 43932 9492
rect 43988 9436 56700 9492
rect 56756 9436 58044 9492
rect 58100 9436 58110 9492
rect 60162 9436 60172 9492
rect 60228 9436 62748 9492
rect 62804 9436 63084 9492
rect 63140 9436 63532 9492
rect 63588 9436 63598 9492
rect 67172 9436 68908 9492
rect 68964 9436 69468 9492
rect 69524 9436 70028 9492
rect 70084 9436 70094 9492
rect 20522 9380 20532 9436
rect 20588 9380 20636 9436
rect 20692 9380 20740 9436
rect 20796 9380 20806 9436
rect 23996 9380 24052 9436
rect 39842 9380 39852 9436
rect 39908 9380 39956 9436
rect 40012 9380 40060 9436
rect 40116 9380 40126 9436
rect 57372 9380 57428 9436
rect 59162 9380 59172 9436
rect 59228 9380 59276 9436
rect 59332 9380 59380 9436
rect 59436 9380 59446 9436
rect 78482 9380 78492 9436
rect 78548 9380 78596 9436
rect 78652 9380 78700 9436
rect 78756 9380 78766 9436
rect 12898 9324 12908 9380
rect 12964 9324 14476 9380
rect 14532 9324 14542 9380
rect 15092 9324 15540 9380
rect 17910 9324 17948 9380
rect 18004 9324 18014 9380
rect 23538 9324 23548 9380
rect 23604 9324 23772 9380
rect 23828 9324 23838 9380
rect 23996 9324 34300 9380
rect 34356 9324 34860 9380
rect 34916 9324 34926 9380
rect 42914 9324 42924 9380
rect 42980 9324 43708 9380
rect 48290 9324 48300 9380
rect 48356 9324 49868 9380
rect 49924 9324 54348 9380
rect 54404 9324 54414 9380
rect 57362 9324 57372 9380
rect 57428 9324 57438 9380
rect 62850 9324 62860 9380
rect 62916 9324 75852 9380
rect 75908 9324 76748 9380
rect 76804 9324 77532 9380
rect 77588 9324 77598 9380
rect 15092 9268 15148 9324
rect 43652 9268 43708 9324
rect 7186 9212 7196 9268
rect 7252 9212 8876 9268
rect 8932 9212 9772 9268
rect 9828 9212 15148 9268
rect 15250 9212 15260 9268
rect 15316 9212 18172 9268
rect 18228 9212 18238 9268
rect 19506 9212 19516 9268
rect 19572 9212 20524 9268
rect 20580 9212 20590 9268
rect 21634 9212 21644 9268
rect 21700 9212 22652 9268
rect 22708 9212 22718 9268
rect 23986 9212 23996 9268
rect 24052 9212 25900 9268
rect 25956 9212 25966 9268
rect 26226 9212 26236 9268
rect 26292 9212 29708 9268
rect 29764 9212 29774 9268
rect 32274 9212 32284 9268
rect 32340 9212 32732 9268
rect 32788 9212 32798 9268
rect 34066 9212 34076 9268
rect 34132 9212 34972 9268
rect 35028 9212 35308 9268
rect 35364 9212 36540 9268
rect 36596 9212 37212 9268
rect 37268 9212 37278 9268
rect 39554 9212 39564 9268
rect 39620 9212 40684 9268
rect 40740 9212 43036 9268
rect 43092 9212 43102 9268
rect 43652 9212 44044 9268
rect 44100 9212 45276 9268
rect 45332 9212 45342 9268
rect 49186 9212 49196 9268
rect 49252 9212 49980 9268
rect 50036 9212 52108 9268
rect 52164 9212 62748 9268
rect 62804 9212 63532 9268
rect 63588 9212 63598 9268
rect 67554 9212 67564 9268
rect 67620 9212 69580 9268
rect 69636 9212 70252 9268
rect 70308 9212 72268 9268
rect 72324 9212 72334 9268
rect 75170 9212 75180 9268
rect 75236 9212 75964 9268
rect 76020 9212 77420 9268
rect 77476 9212 77486 9268
rect 4498 9100 4508 9156
rect 4564 9100 5740 9156
rect 5796 9100 6524 9156
rect 6580 9100 6590 9156
rect 10882 9100 10892 9156
rect 10948 9100 12012 9156
rect 12068 9100 13580 9156
rect 13636 9100 13646 9156
rect 18274 9100 18284 9156
rect 18340 9100 19292 9156
rect 19348 9100 19358 9156
rect 24322 9100 24332 9156
rect 24388 9100 26012 9156
rect 26068 9100 26348 9156
rect 26404 9100 26414 9156
rect 29474 9100 29484 9156
rect 29540 9100 30044 9156
rect 30100 9100 30604 9156
rect 30660 9100 30670 9156
rect 34850 9100 34860 9156
rect 34916 9100 40012 9156
rect 40068 9100 40572 9156
rect 40628 9100 40638 9156
rect 42354 9100 42364 9156
rect 42420 9100 48748 9156
rect 48804 9100 49420 9156
rect 49476 9100 49756 9156
rect 49812 9100 50876 9156
rect 50932 9100 50942 9156
rect 54786 9100 54796 9156
rect 54852 9100 56140 9156
rect 56196 9100 56206 9156
rect 61506 9100 61516 9156
rect 61572 9100 66780 9156
rect 66836 9100 67452 9156
rect 67508 9100 69020 9156
rect 69076 9100 69086 9156
rect 75618 9100 75628 9156
rect 75684 9100 76860 9156
rect 76916 9100 76926 9156
rect 4274 8988 4284 9044
rect 4340 8988 5516 9044
rect 5572 8988 5582 9044
rect 6738 8988 6748 9044
rect 6804 8988 7084 9044
rect 7140 8988 8540 9044
rect 8596 8988 8606 9044
rect 10434 8988 10444 9044
rect 10500 8988 11900 9044
rect 11956 8988 11966 9044
rect 17042 8988 17052 9044
rect 17108 8988 18060 9044
rect 18116 8988 22316 9044
rect 22372 8988 22382 9044
rect 28130 8988 28140 9044
rect 28196 8988 28700 9044
rect 28756 8988 29932 9044
rect 29988 8988 30492 9044
rect 30548 8988 30558 9044
rect 31490 8988 31500 9044
rect 31556 8988 34188 9044
rect 34244 8988 34254 9044
rect 40898 8988 40908 9044
rect 40964 8988 41580 9044
rect 41636 8988 41646 9044
rect 43652 8988 50764 9044
rect 50820 8988 50830 9044
rect 54674 8988 54684 9044
rect 54740 8988 55916 9044
rect 55972 8988 55982 9044
rect 64082 8988 64092 9044
rect 64148 8988 65436 9044
rect 65492 8988 65502 9044
rect 68338 8988 68348 9044
rect 68404 8988 69132 9044
rect 69188 8988 69198 9044
rect 70354 8988 70364 9044
rect 70420 8988 71596 9044
rect 71652 8988 71662 9044
rect 71922 8988 71932 9044
rect 71988 8988 73948 9044
rect 74004 8988 74014 9044
rect 74946 8988 74956 9044
rect 75012 8988 76748 9044
rect 76804 8988 76814 9044
rect 0 8932 800 8960
rect 0 8876 1932 8932
rect 1988 8876 1998 8932
rect 18610 8876 18620 8932
rect 18676 8876 20972 8932
rect 21028 8876 21038 8932
rect 37538 8876 37548 8932
rect 37604 8876 42252 8932
rect 42308 8876 42318 8932
rect 0 8848 800 8876
rect 43652 8820 43708 8988
rect 68348 8932 68404 8988
rect 79200 8932 80000 8960
rect 52770 8876 52780 8932
rect 52836 8876 54796 8932
rect 54852 8876 54862 8932
rect 56018 8876 56028 8932
rect 56084 8876 60844 8932
rect 60900 8876 62412 8932
rect 62468 8876 62478 8932
rect 65202 8876 65212 8932
rect 65268 8876 65772 8932
rect 65828 8876 65838 8932
rect 68002 8876 68012 8932
rect 68068 8876 68404 8932
rect 69794 8876 69804 8932
rect 69860 8876 70476 8932
rect 70532 8876 70542 8932
rect 70914 8876 70924 8932
rect 70980 8876 73052 8932
rect 73108 8876 73118 8932
rect 75506 8876 75516 8932
rect 75572 8876 80000 8932
rect 79200 8848 80000 8876
rect 28802 8764 28812 8820
rect 28868 8764 29708 8820
rect 29764 8764 31444 8820
rect 36530 8764 36540 8820
rect 36596 8764 40460 8820
rect 40516 8764 40526 8820
rect 41682 8764 41692 8820
rect 41748 8764 43708 8820
rect 45266 8764 45276 8820
rect 45332 8764 65100 8820
rect 65156 8764 65324 8820
rect 65380 8764 65390 8820
rect 31388 8708 31444 8764
rect 5394 8652 5404 8708
rect 5460 8652 9884 8708
rect 9940 8652 9950 8708
rect 31388 8652 42700 8708
rect 42756 8652 42766 8708
rect 43250 8652 43260 8708
rect 43316 8652 49196 8708
rect 49252 8652 49262 8708
rect 10862 8596 10872 8652
rect 10928 8596 10976 8652
rect 11032 8596 11080 8652
rect 11136 8596 11146 8652
rect 30182 8596 30192 8652
rect 30248 8596 30296 8652
rect 30352 8596 30400 8652
rect 30456 8596 30466 8652
rect 49502 8596 49512 8652
rect 49568 8596 49616 8652
rect 49672 8596 49720 8652
rect 49776 8596 49786 8652
rect 68822 8596 68832 8652
rect 68888 8596 68936 8652
rect 68992 8596 69040 8652
rect 69096 8596 69106 8652
rect 4946 8540 4956 8596
rect 5012 8540 10444 8596
rect 10500 8540 10510 8596
rect 20514 8540 20524 8596
rect 20580 8540 21420 8596
rect 21476 8540 26908 8596
rect 32834 8540 32844 8596
rect 32900 8540 33068 8596
rect 33124 8540 33134 8596
rect 40562 8540 40572 8596
rect 40628 8540 41692 8596
rect 41748 8540 41758 8596
rect 65772 8540 66332 8596
rect 66388 8540 66780 8596
rect 66836 8540 66846 8596
rect 77858 8540 77868 8596
rect 77924 8540 77934 8596
rect 26852 8484 26908 8540
rect 65772 8484 65828 8540
rect 8194 8428 8204 8484
rect 8260 8428 8932 8484
rect 16146 8428 16156 8484
rect 16212 8428 21196 8484
rect 21252 8428 21262 8484
rect 22652 8428 23548 8484
rect 23604 8428 23614 8484
rect 26852 8428 35756 8484
rect 35812 8428 35822 8484
rect 37314 8428 37324 8484
rect 37380 8428 37884 8484
rect 37940 8428 42924 8484
rect 42980 8428 42990 8484
rect 65314 8428 65324 8484
rect 65380 8428 65772 8484
rect 65828 8428 65838 8484
rect 66658 8428 66668 8484
rect 66724 8428 66734 8484
rect 8876 8372 8932 8428
rect 22652 8372 22708 8428
rect 66668 8372 66724 8428
rect 77868 8372 77924 8540
rect 2146 8316 2156 8372
rect 2212 8316 3836 8372
rect 3892 8316 3902 8372
rect 7186 8316 7196 8372
rect 7252 8316 7756 8372
rect 7812 8316 8652 8372
rect 8708 8316 8718 8372
rect 8866 8316 8876 8372
rect 8932 8316 9660 8372
rect 9716 8316 19908 8372
rect 20066 8316 20076 8372
rect 20132 8316 22708 8372
rect 24210 8316 24220 8372
rect 24276 8316 29596 8372
rect 29652 8316 29662 8372
rect 38220 8316 40796 8372
rect 40852 8316 41580 8372
rect 41636 8316 41646 8372
rect 55570 8316 55580 8372
rect 55636 8316 56700 8372
rect 56756 8316 56766 8372
rect 60386 8316 60396 8372
rect 60452 8316 61628 8372
rect 61684 8316 62412 8372
rect 62468 8316 62478 8372
rect 62962 8316 62972 8372
rect 63028 8316 63756 8372
rect 63812 8316 63822 8372
rect 66668 8316 67564 8372
rect 67620 8316 67630 8372
rect 75394 8316 75404 8372
rect 75460 8316 76636 8372
rect 76692 8316 76702 8372
rect 77298 8316 77308 8372
rect 77364 8316 77924 8372
rect 19852 8260 19908 8316
rect 4610 8204 4620 8260
rect 4676 8204 7868 8260
rect 7924 8204 7934 8260
rect 8306 8204 8316 8260
rect 8372 8204 9772 8260
rect 9828 8204 9838 8260
rect 14578 8204 14588 8260
rect 14644 8204 15260 8260
rect 15316 8204 15326 8260
rect 16594 8204 16604 8260
rect 16660 8204 17164 8260
rect 17220 8204 18620 8260
rect 18676 8204 18686 8260
rect 19852 8204 22484 8260
rect 22642 8204 22652 8260
rect 22708 8204 23436 8260
rect 23492 8204 23502 8260
rect 22428 8148 22484 8204
rect 26852 8148 26908 8260
rect 26964 8204 28476 8260
rect 28532 8204 28542 8260
rect 28802 8204 28812 8260
rect 28868 8204 31388 8260
rect 31444 8204 31724 8260
rect 31780 8204 31790 8260
rect 36754 8204 36764 8260
rect 36820 8204 37772 8260
rect 37828 8204 37838 8260
rect 38220 8148 38276 8316
rect 43474 8204 43484 8260
rect 43540 8204 46284 8260
rect 46340 8204 46350 8260
rect 46722 8204 46732 8260
rect 46788 8204 47404 8260
rect 47460 8204 47470 8260
rect 50306 8204 50316 8260
rect 50372 8204 50764 8260
rect 50820 8204 50830 8260
rect 57474 8204 57484 8260
rect 57540 8204 58380 8260
rect 58436 8204 58446 8260
rect 58818 8204 58828 8260
rect 58884 8204 59612 8260
rect 59668 8204 59678 8260
rect 60274 8204 60284 8260
rect 60340 8204 61068 8260
rect 61124 8204 64988 8260
rect 65044 8204 69692 8260
rect 69748 8204 69758 8260
rect 72034 8204 72044 8260
rect 72100 8204 72716 8260
rect 72772 8204 73388 8260
rect 73444 8204 73454 8260
rect 73602 8204 73612 8260
rect 73668 8204 74620 8260
rect 74676 8204 75516 8260
rect 75572 8204 75582 8260
rect 76850 8204 76860 8260
rect 76916 8204 77532 8260
rect 77588 8204 77598 8260
rect 46284 8148 46340 8204
rect 5842 8092 5852 8148
rect 5908 8092 9324 8148
rect 9380 8092 9390 8148
rect 19058 8092 19068 8148
rect 19124 8092 20188 8148
rect 20244 8092 20254 8148
rect 22428 8092 26348 8148
rect 26404 8092 26908 8148
rect 27234 8092 27244 8148
rect 27300 8092 28028 8148
rect 28084 8092 31612 8148
rect 31668 8092 31678 8148
rect 36866 8092 36876 8148
rect 36932 8092 38220 8148
rect 38276 8092 38286 8148
rect 38612 8092 45388 8148
rect 45444 8092 45454 8148
rect 46284 8092 47628 8148
rect 47684 8092 47694 8148
rect 54226 8092 54236 8148
rect 54292 8092 55132 8148
rect 55188 8092 59052 8148
rect 59108 8092 59118 8148
rect 68460 8092 69804 8148
rect 69860 8092 69870 8148
rect 70354 8092 70364 8148
rect 70420 8092 71148 8148
rect 71204 8092 71214 8148
rect 74508 8092 75292 8148
rect 75348 8092 76300 8148
rect 76356 8092 77308 8148
rect 77364 8092 77374 8148
rect 38612 8036 38668 8092
rect 3154 7980 3164 8036
rect 3220 7980 3724 8036
rect 3780 7980 3790 8036
rect 8194 7980 8204 8036
rect 8260 7980 9996 8036
rect 10052 7980 10668 8036
rect 10724 7980 10734 8036
rect 15810 7980 15820 8036
rect 15876 7980 18508 8036
rect 18564 7980 19964 8036
rect 20020 7980 20030 8036
rect 21634 7980 21644 8036
rect 21700 7980 22428 8036
rect 22484 7980 23548 8036
rect 23604 7980 24668 8036
rect 24724 7980 24734 8036
rect 27682 7980 27692 8036
rect 27748 7980 38668 8036
rect 48514 7980 48524 8036
rect 48580 7980 49196 8036
rect 49252 7980 49262 8036
rect 57362 7980 57372 8036
rect 57428 7980 57932 8036
rect 57988 7980 57998 8036
rect 58370 7980 58380 8036
rect 58436 7980 64260 8036
rect 64204 7924 64260 7980
rect 68460 7924 68516 8092
rect 74508 8036 74564 8092
rect 69244 7980 74564 8036
rect 74722 7980 74732 8036
rect 74788 7980 75964 8036
rect 76020 7980 76030 8036
rect 1810 7868 1820 7924
rect 1876 7868 2492 7924
rect 2548 7868 3276 7924
rect 3332 7868 5964 7924
rect 6020 7868 6188 7924
rect 6244 7868 10108 7924
rect 10164 7868 10892 7924
rect 10948 7868 10958 7924
rect 22530 7868 22540 7924
rect 22596 7868 33404 7924
rect 33460 7868 33470 7924
rect 40674 7868 40684 7924
rect 40740 7868 43260 7924
rect 43316 7868 50652 7924
rect 50708 7868 52332 7924
rect 52388 7868 52398 7924
rect 64204 7868 65548 7924
rect 65604 7868 66556 7924
rect 66612 7868 66622 7924
rect 66780 7868 67900 7924
rect 67956 7868 68460 7924
rect 68516 7868 68526 7924
rect 4722 7644 4732 7700
rect 4788 7644 4798 7700
rect 4732 7588 4788 7644
rect 9772 7588 9828 7868
rect 20522 7812 20532 7868
rect 20588 7812 20636 7868
rect 20692 7812 20740 7868
rect 20796 7812 20806 7868
rect 39842 7812 39852 7868
rect 39908 7812 39956 7868
rect 40012 7812 40060 7868
rect 40116 7812 40126 7868
rect 59162 7812 59172 7868
rect 59228 7812 59276 7868
rect 59332 7812 59380 7868
rect 59436 7812 59446 7868
rect 66780 7812 66836 7868
rect 69244 7812 69300 7980
rect 78482 7812 78492 7868
rect 78548 7812 78596 7868
rect 78652 7812 78700 7868
rect 78756 7812 78766 7868
rect 10658 7756 10668 7812
rect 10724 7756 20356 7812
rect 20300 7700 20356 7756
rect 21980 7756 26684 7812
rect 26740 7756 26750 7812
rect 36418 7756 36428 7812
rect 36484 7756 37772 7812
rect 37828 7756 37838 7812
rect 46834 7756 46844 7812
rect 46900 7756 51772 7812
rect 51828 7756 52444 7812
rect 52500 7756 53340 7812
rect 53396 7756 53406 7812
rect 61282 7756 61292 7812
rect 61348 7756 66836 7812
rect 67228 7756 69300 7812
rect 69682 7756 69692 7812
rect 69748 7756 73276 7812
rect 73332 7756 73342 7812
rect 21980 7700 22036 7756
rect 37772 7700 37828 7756
rect 67228 7700 67284 7756
rect 13458 7644 13468 7700
rect 13524 7644 14252 7700
rect 14308 7644 14588 7700
rect 14644 7644 14654 7700
rect 14914 7644 14924 7700
rect 14980 7644 15372 7700
rect 15428 7644 15438 7700
rect 15922 7644 15932 7700
rect 15988 7644 16604 7700
rect 16660 7644 16670 7700
rect 20300 7644 22036 7700
rect 22194 7644 22204 7700
rect 22260 7644 23660 7700
rect 23716 7644 23726 7700
rect 37772 7644 42028 7700
rect 42084 7644 42094 7700
rect 48178 7644 48188 7700
rect 48244 7644 48636 7700
rect 48692 7644 49644 7700
rect 49700 7644 60732 7700
rect 60788 7644 60798 7700
rect 63074 7644 63084 7700
rect 63140 7644 63532 7700
rect 63588 7644 63598 7700
rect 67172 7644 67284 7700
rect 67442 7644 67452 7700
rect 67508 7644 68460 7700
rect 68516 7644 68526 7700
rect 69906 7644 69916 7700
rect 69972 7644 71372 7700
rect 71428 7644 71438 7700
rect 1362 7532 1372 7588
rect 1428 7532 2492 7588
rect 2548 7532 2716 7588
rect 2772 7532 2782 7588
rect 4162 7532 4172 7588
rect 4228 7532 6412 7588
rect 6468 7532 6478 7588
rect 9762 7532 9772 7588
rect 9828 7532 9838 7588
rect 15092 7532 21644 7588
rect 21700 7532 21710 7588
rect 22082 7532 22092 7588
rect 22148 7532 22764 7588
rect 22820 7532 23884 7588
rect 23940 7532 23950 7588
rect 26338 7532 26348 7588
rect 26404 7532 29484 7588
rect 29540 7532 29820 7588
rect 29876 7532 43708 7588
rect 48850 7532 48860 7588
rect 48916 7532 49308 7588
rect 49364 7532 50428 7588
rect 50484 7532 58828 7588
rect 58884 7532 58894 7588
rect 15092 7476 15148 7532
rect 43652 7476 43708 7532
rect 3602 7420 3612 7476
rect 3668 7420 4508 7476
rect 4564 7420 5740 7476
rect 5796 7420 5806 7476
rect 9884 7420 15148 7476
rect 31154 7420 31164 7476
rect 31220 7420 32620 7476
rect 32676 7420 32686 7476
rect 32844 7420 42924 7476
rect 42980 7420 42990 7476
rect 43652 7420 43932 7476
rect 43988 7420 43998 7476
rect 51538 7420 51548 7476
rect 51604 7420 54572 7476
rect 54628 7420 54638 7476
rect 58034 7420 58044 7476
rect 58100 7420 61292 7476
rect 61348 7420 61358 7476
rect 64978 7420 64988 7476
rect 65044 7420 65436 7476
rect 65492 7420 66108 7476
rect 66164 7420 66174 7476
rect 9884 7364 9940 7420
rect 32844 7364 32900 7420
rect 67172 7364 67228 7644
rect 67340 7532 67564 7588
rect 67620 7532 68124 7588
rect 68180 7532 70588 7588
rect 70644 7532 70654 7588
rect 67340 7476 67396 7532
rect 67330 7420 67340 7476
rect 67396 7420 67406 7476
rect 67666 7420 67676 7476
rect 67732 7420 69356 7476
rect 69412 7420 71708 7476
rect 71764 7420 71774 7476
rect 4610 7308 4620 7364
rect 4676 7308 9940 7364
rect 14914 7308 14924 7364
rect 14980 7308 15820 7364
rect 15876 7308 15886 7364
rect 20402 7308 20412 7364
rect 20468 7308 22316 7364
rect 22372 7308 23996 7364
rect 24052 7308 24062 7364
rect 24210 7308 24220 7364
rect 24276 7308 25340 7364
rect 25396 7308 25406 7364
rect 30930 7308 30940 7364
rect 30996 7308 32900 7364
rect 35186 7308 35196 7364
rect 35252 7308 36316 7364
rect 36372 7308 37548 7364
rect 37604 7308 37614 7364
rect 38434 7308 38444 7364
rect 38500 7308 43036 7364
rect 43092 7308 44492 7364
rect 44548 7308 44558 7364
rect 51874 7308 51884 7364
rect 51940 7308 52332 7364
rect 52388 7308 52668 7364
rect 52724 7308 53788 7364
rect 53844 7308 55692 7364
rect 55748 7308 57372 7364
rect 57428 7308 57438 7364
rect 58370 7308 58380 7364
rect 58436 7308 60620 7364
rect 60676 7308 60686 7364
rect 63186 7308 63196 7364
rect 63252 7308 67228 7364
rect 69570 7308 69580 7364
rect 69636 7308 71820 7364
rect 71876 7308 71886 7364
rect 37202 7196 37212 7252
rect 37268 7196 37660 7252
rect 37716 7196 38332 7252
rect 38388 7196 39844 7252
rect 42802 7196 42812 7252
rect 42868 7196 45388 7252
rect 45444 7196 45454 7252
rect 47282 7196 47292 7252
rect 47348 7196 48412 7252
rect 48468 7196 51324 7252
rect 51380 7196 51390 7252
rect 58034 7196 58044 7252
rect 58100 7196 59388 7252
rect 59444 7196 60060 7252
rect 60116 7196 60126 7252
rect 39788 7140 39844 7196
rect 38612 7084 39564 7140
rect 39620 7084 39630 7140
rect 39788 7084 48524 7140
rect 48580 7084 48590 7140
rect 58930 7084 58940 7140
rect 58996 7084 60284 7140
rect 60340 7084 61404 7140
rect 61460 7084 64876 7140
rect 64932 7084 64942 7140
rect 65650 7084 65660 7140
rect 65716 7084 67676 7140
rect 67732 7084 67742 7140
rect 10862 7028 10872 7084
rect 10928 7028 10976 7084
rect 11032 7028 11080 7084
rect 11136 7028 11146 7084
rect 30182 7028 30192 7084
rect 30248 7028 30296 7084
rect 30352 7028 30400 7084
rect 30456 7028 30466 7084
rect 28242 6972 28252 7028
rect 28308 6972 28588 7028
rect 28644 6972 28654 7028
rect 38612 6916 38668 7084
rect 49502 7028 49512 7084
rect 49568 7028 49616 7084
rect 49672 7028 49720 7084
rect 49776 7028 49786 7084
rect 68822 7028 68832 7084
rect 68888 7028 68936 7084
rect 68992 7028 69040 7084
rect 69096 7028 69106 7084
rect 38882 6972 38892 7028
rect 38948 6972 49196 7028
rect 49252 6972 49262 7028
rect 49868 6972 53004 7028
rect 53060 6972 53676 7028
rect 53732 6972 53742 7028
rect 54674 6972 54684 7028
rect 54740 6972 55356 7028
rect 55412 6972 55422 7028
rect 55906 6972 55916 7028
rect 55972 6972 62076 7028
rect 62132 6972 62860 7028
rect 62916 6972 62926 7028
rect 49868 6916 49924 6972
rect 9314 6860 9324 6916
rect 9380 6860 38668 6916
rect 47394 6860 47404 6916
rect 47460 6860 49924 6916
rect 50082 6860 50092 6916
rect 50148 6860 50876 6916
rect 50932 6860 50942 6916
rect 52882 6860 52892 6916
rect 52948 6860 54348 6916
rect 54404 6860 56868 6916
rect 63830 6860 63868 6916
rect 63924 6860 63934 6916
rect 66434 6860 66444 6916
rect 66500 6860 69580 6916
rect 69636 6860 69646 6916
rect 9650 6748 9660 6804
rect 9716 6748 9996 6804
rect 10052 6748 10062 6804
rect 12898 6748 12908 6804
rect 12964 6748 13132 6804
rect 13188 6748 13692 6804
rect 13748 6748 13758 6804
rect 28130 6748 28140 6804
rect 28196 6748 28206 6804
rect 28914 6748 28924 6804
rect 28980 6748 29484 6804
rect 29540 6748 29550 6804
rect 31490 6748 31500 6804
rect 31556 6748 32060 6804
rect 32116 6748 32126 6804
rect 43474 6748 43484 6804
rect 43540 6748 44156 6804
rect 44212 6748 44222 6804
rect 45938 6748 45948 6804
rect 46004 6748 46620 6804
rect 46676 6748 46686 6804
rect 47842 6748 47852 6804
rect 47908 6748 52332 6804
rect 52388 6748 52398 6804
rect 28140 6692 28196 6748
rect 56812 6692 56868 6860
rect 59042 6748 59052 6804
rect 59108 6748 74284 6804
rect 74340 6748 74350 6804
rect 76066 6748 76076 6804
rect 76132 6748 77532 6804
rect 77588 6748 77598 6804
rect 8642 6636 8652 6692
rect 8708 6636 9324 6692
rect 9380 6636 10220 6692
rect 10276 6636 10286 6692
rect 10434 6636 10444 6692
rect 10500 6636 10892 6692
rect 10948 6636 12572 6692
rect 12628 6636 12638 6692
rect 15586 6636 15596 6692
rect 15652 6636 16044 6692
rect 16100 6636 16268 6692
rect 16324 6636 16334 6692
rect 22642 6636 22652 6692
rect 22708 6636 23548 6692
rect 23604 6636 23614 6692
rect 24322 6636 24332 6692
rect 24388 6636 25116 6692
rect 25172 6636 26012 6692
rect 26068 6636 26078 6692
rect 28140 6636 28812 6692
rect 28868 6636 28878 6692
rect 31602 6636 31612 6692
rect 31668 6636 32396 6692
rect 32452 6636 34972 6692
rect 35028 6636 35038 6692
rect 39666 6636 39676 6692
rect 39732 6636 41356 6692
rect 41412 6636 42588 6692
rect 42644 6636 42654 6692
rect 51202 6636 51212 6692
rect 51268 6636 51996 6692
rect 52052 6636 52556 6692
rect 52612 6636 52622 6692
rect 52770 6636 52780 6692
rect 52836 6636 55580 6692
rect 55636 6636 55646 6692
rect 55794 6636 55804 6692
rect 55860 6636 55898 6692
rect 56018 6636 56028 6692
rect 56084 6636 56476 6692
rect 56532 6636 56542 6692
rect 56802 6636 56812 6692
rect 56868 6636 56878 6692
rect 57810 6636 57820 6692
rect 57876 6636 59724 6692
rect 59780 6636 59790 6692
rect 59938 6636 59948 6692
rect 60004 6636 61068 6692
rect 61124 6636 61134 6692
rect 63746 6636 63756 6692
rect 63812 6636 64764 6692
rect 64820 6636 65660 6692
rect 65716 6636 65726 6692
rect 68338 6636 68348 6692
rect 68404 6636 68572 6692
rect 68628 6636 70028 6692
rect 70084 6636 70094 6692
rect 70914 6636 70924 6692
rect 70980 6636 73164 6692
rect 73220 6636 73230 6692
rect 75282 6636 75292 6692
rect 75348 6636 77420 6692
rect 77476 6636 77486 6692
rect 9426 6524 9436 6580
rect 9492 6524 9884 6580
rect 9940 6524 15148 6580
rect 24098 6524 24108 6580
rect 24164 6524 24780 6580
rect 24836 6524 25228 6580
rect 25284 6524 25564 6580
rect 25620 6524 25630 6580
rect 28130 6524 28140 6580
rect 28196 6524 31052 6580
rect 31108 6524 32060 6580
rect 32116 6524 32126 6580
rect 34850 6524 34860 6580
rect 34916 6524 36428 6580
rect 36484 6524 36494 6580
rect 39330 6524 39340 6580
rect 39396 6524 40124 6580
rect 40180 6524 40190 6580
rect 48850 6524 48860 6580
rect 48916 6524 49980 6580
rect 50036 6524 50046 6580
rect 51426 6524 51436 6580
rect 51492 6524 55468 6580
rect 55524 6524 56588 6580
rect 56644 6524 56654 6580
rect 58146 6524 58156 6580
rect 58212 6524 59164 6580
rect 59220 6524 60508 6580
rect 60564 6524 60574 6580
rect 67218 6524 67228 6580
rect 67284 6524 70252 6580
rect 70308 6524 70318 6580
rect 72258 6524 72268 6580
rect 72324 6524 77308 6580
rect 77364 6524 77374 6580
rect 0 6468 800 6496
rect 15092 6468 15148 6524
rect 79200 6468 80000 6496
rect 0 6412 1932 6468
rect 1988 6412 1998 6468
rect 3714 6412 3724 6468
rect 3780 6412 5068 6468
rect 5124 6412 5134 6468
rect 8642 6412 8652 6468
rect 8708 6412 10108 6468
rect 10164 6412 10174 6468
rect 10322 6412 10332 6468
rect 10388 6412 11340 6468
rect 11396 6412 11406 6468
rect 12002 6412 12012 6468
rect 12068 6412 12684 6468
rect 12740 6412 14812 6468
rect 14868 6412 14878 6468
rect 15092 6412 25788 6468
rect 25844 6412 28028 6468
rect 28084 6412 28094 6468
rect 34178 6412 34188 6468
rect 34244 6412 35084 6468
rect 35140 6412 35150 6468
rect 35970 6412 35980 6468
rect 36036 6412 37436 6468
rect 37492 6412 37660 6468
rect 37716 6412 37726 6468
rect 40338 6412 40348 6468
rect 40404 6412 41244 6468
rect 41300 6412 41310 6468
rect 46498 6412 46508 6468
rect 46564 6412 47068 6468
rect 47124 6412 47134 6468
rect 51090 6412 51100 6468
rect 51156 6412 53564 6468
rect 53620 6412 53630 6468
rect 56028 6412 57372 6468
rect 57428 6412 60172 6468
rect 60228 6412 60238 6468
rect 64530 6412 64540 6468
rect 64596 6412 65212 6468
rect 65268 6412 65278 6468
rect 65762 6412 65772 6468
rect 65828 6412 67900 6468
rect 67956 6412 67966 6468
rect 68898 6412 68908 6468
rect 68964 6412 69468 6468
rect 69524 6412 71036 6468
rect 71092 6412 71102 6468
rect 71474 6412 71484 6468
rect 71540 6412 72380 6468
rect 72436 6412 72716 6468
rect 72772 6412 72782 6468
rect 74050 6412 74060 6468
rect 74116 6412 74620 6468
rect 74676 6412 74686 6468
rect 75058 6412 75068 6468
rect 75124 6412 80000 6468
rect 0 6384 800 6412
rect 3490 6300 3500 6356
rect 3556 6300 4508 6356
rect 4564 6300 4732 6356
rect 4788 6300 6076 6356
rect 6132 6300 14252 6356
rect 14308 6300 14318 6356
rect 20962 6300 20972 6356
rect 21028 6300 23772 6356
rect 23828 6300 24444 6356
rect 24500 6300 24510 6356
rect 30594 6300 30604 6356
rect 30660 6300 39676 6356
rect 39732 6300 39742 6356
rect 44594 6300 44604 6356
rect 44660 6300 45948 6356
rect 46004 6300 47852 6356
rect 47908 6300 47918 6356
rect 48738 6300 48748 6356
rect 48804 6300 54460 6356
rect 54516 6300 54526 6356
rect 20522 6244 20532 6300
rect 20588 6244 20636 6300
rect 20692 6244 20740 6300
rect 20796 6244 20806 6300
rect 39842 6244 39852 6300
rect 39908 6244 39956 6300
rect 40012 6244 40060 6300
rect 40116 6244 40126 6300
rect 56028 6244 56084 6412
rect 71036 6356 71092 6412
rect 79200 6384 80000 6412
rect 56690 6300 56700 6356
rect 56756 6300 57932 6356
rect 57988 6300 57998 6356
rect 60050 6300 60060 6356
rect 60116 6300 63420 6356
rect 63476 6300 63486 6356
rect 66658 6300 66668 6356
rect 66724 6300 67340 6356
rect 67396 6300 67406 6356
rect 67666 6300 67676 6356
rect 67732 6300 70700 6356
rect 70756 6300 70766 6356
rect 71036 6300 73612 6356
rect 73668 6300 73678 6356
rect 59162 6244 59172 6300
rect 59228 6244 59276 6300
rect 59332 6244 59380 6300
rect 59436 6244 59446 6300
rect 78482 6244 78492 6300
rect 78548 6244 78596 6300
rect 78652 6244 78700 6300
rect 78756 6244 78766 6300
rect 9986 6188 9996 6244
rect 10052 6188 11116 6244
rect 11172 6188 11182 6244
rect 23202 6188 23212 6244
rect 23268 6188 23660 6244
rect 23716 6188 23726 6244
rect 27010 6188 27020 6244
rect 27076 6188 38668 6244
rect 42914 6188 42924 6244
rect 42980 6188 49756 6244
rect 49812 6188 52444 6244
rect 52500 6188 52510 6244
rect 56018 6188 56028 6244
rect 56084 6188 56094 6244
rect 61842 6188 61852 6244
rect 61908 6188 63756 6244
rect 63812 6188 64316 6244
rect 64372 6188 64988 6244
rect 65044 6188 65054 6244
rect 66546 6188 66556 6244
rect 66612 6188 67228 6244
rect 67284 6188 67294 6244
rect 38612 6132 38668 6188
rect 8530 6076 8540 6132
rect 8596 6076 8876 6132
rect 8932 6076 9548 6132
rect 9604 6076 9716 6132
rect 9874 6076 9884 6132
rect 9940 6076 10444 6132
rect 10500 6076 24276 6132
rect 36978 6076 36988 6132
rect 37044 6076 38276 6132
rect 38612 6076 46172 6132
rect 46228 6076 47516 6132
rect 47572 6076 48300 6132
rect 48356 6076 48366 6132
rect 48626 6076 48636 6132
rect 48692 6076 49868 6132
rect 49924 6076 49934 6132
rect 51324 6076 52108 6132
rect 52164 6076 53340 6132
rect 53396 6076 55916 6132
rect 55972 6076 55982 6132
rect 56130 6076 56140 6132
rect 56196 6076 57036 6132
rect 57092 6076 58940 6132
rect 58996 6076 59006 6132
rect 59164 6076 67228 6132
rect 67284 6076 67294 6132
rect 67442 6076 67452 6132
rect 67508 6076 69804 6132
rect 69860 6076 70588 6132
rect 70644 6076 70654 6132
rect 74498 6076 74508 6132
rect 74564 6076 77756 6132
rect 77812 6076 77822 6132
rect 9660 6020 9716 6076
rect 5618 5964 5628 6020
rect 5684 5964 6748 6020
rect 6804 5964 7420 6020
rect 7476 5964 8428 6020
rect 8484 5964 9436 6020
rect 9492 5964 9502 6020
rect 9660 5964 10332 6020
rect 10388 5964 10398 6020
rect 18498 5964 18508 6020
rect 18564 5964 19516 6020
rect 19572 5964 19582 6020
rect 5394 5852 5404 5908
rect 5460 5852 8652 5908
rect 8708 5852 8718 5908
rect 16482 5852 16492 5908
rect 16548 5852 17612 5908
rect 17668 5852 17678 5908
rect 18274 5852 18284 5908
rect 18340 5852 22876 5908
rect 22932 5852 22942 5908
rect 24220 5796 24276 6076
rect 38220 6020 38276 6076
rect 48300 6020 48356 6076
rect 51324 6020 51380 6076
rect 59164 6020 59220 6076
rect 25106 5964 25116 6020
rect 25172 5964 25676 6020
rect 25732 5964 25742 6020
rect 35074 5964 35084 6020
rect 35140 5964 36540 6020
rect 36596 5964 37996 6020
rect 38052 5964 38062 6020
rect 38220 5964 40852 6020
rect 40796 5908 40852 5964
rect 45724 5964 46732 6020
rect 46788 5964 46798 6020
rect 48300 5964 49644 6020
rect 49700 5964 49710 6020
rect 49970 5964 49980 6020
rect 50036 5964 51380 6020
rect 51538 5964 51548 6020
rect 51604 5964 53900 6020
rect 53956 5964 53966 6020
rect 54674 5964 54684 6020
rect 54740 5964 55356 6020
rect 55412 5964 56028 6020
rect 56084 5964 56094 6020
rect 56242 5964 56252 6020
rect 56308 5964 57708 6020
rect 57764 5964 58156 6020
rect 58212 5964 58222 6020
rect 58370 5964 58380 6020
rect 58436 5964 59220 6020
rect 62178 5964 62188 6020
rect 62244 5964 62972 6020
rect 63028 5964 63038 6020
rect 64418 5964 64428 6020
rect 64484 5964 66556 6020
rect 66612 5964 66622 6020
rect 67106 5964 67116 6020
rect 67172 5964 67452 6020
rect 67508 5964 70924 6020
rect 70980 5964 70990 6020
rect 45724 5908 45780 5964
rect 24434 5852 24444 5908
rect 24500 5852 29540 5908
rect 29698 5852 29708 5908
rect 29764 5852 30044 5908
rect 30100 5852 30940 5908
rect 30996 5852 31006 5908
rect 32722 5852 32732 5908
rect 32788 5852 38668 5908
rect 38724 5852 39340 5908
rect 39396 5852 39564 5908
rect 39620 5852 39630 5908
rect 40786 5852 40796 5908
rect 40852 5852 42140 5908
rect 42196 5852 45780 5908
rect 45836 5852 50092 5908
rect 50148 5852 51996 5908
rect 52052 5852 54908 5908
rect 54964 5852 55468 5908
rect 55524 5852 55534 5908
rect 55906 5852 55916 5908
rect 55972 5852 58828 5908
rect 58884 5852 58894 5908
rect 62514 5852 62524 5908
rect 62580 5852 63644 5908
rect 63700 5852 63710 5908
rect 65426 5852 65436 5908
rect 65492 5852 65884 5908
rect 65940 5852 65950 5908
rect 66882 5852 66892 5908
rect 66948 5852 68124 5908
rect 68180 5852 69692 5908
rect 69748 5852 69758 5908
rect 72034 5852 72044 5908
rect 72100 5852 72492 5908
rect 72548 5852 72558 5908
rect 76962 5852 76972 5908
rect 77028 5852 77532 5908
rect 77588 5852 77598 5908
rect 29484 5796 29540 5852
rect 45836 5796 45892 5852
rect 65884 5796 65940 5852
rect 8978 5740 8988 5796
rect 9044 5740 9996 5796
rect 10052 5740 10062 5796
rect 14690 5740 14700 5796
rect 14756 5740 21980 5796
rect 22036 5740 22046 5796
rect 22530 5740 22540 5796
rect 22596 5740 23436 5796
rect 23492 5740 23502 5796
rect 24220 5740 27468 5796
rect 27524 5740 27534 5796
rect 29484 5740 30380 5796
rect 30436 5740 30446 5796
rect 35522 5740 35532 5796
rect 35588 5740 36316 5796
rect 36372 5740 36876 5796
rect 36932 5740 45892 5796
rect 46050 5740 46060 5796
rect 46116 5740 48188 5796
rect 48244 5740 48254 5796
rect 49522 5740 49532 5796
rect 49588 5740 50652 5796
rect 50708 5740 50718 5796
rect 51202 5740 51212 5796
rect 51268 5740 54796 5796
rect 54852 5740 57596 5796
rect 57652 5740 57662 5796
rect 58034 5740 58044 5796
rect 58100 5740 58492 5796
rect 58548 5740 59948 5796
rect 60004 5740 60014 5796
rect 61058 5740 61068 5796
rect 61124 5740 64652 5796
rect 64708 5740 64718 5796
rect 65884 5740 69356 5796
rect 69412 5740 69422 5796
rect 72594 5740 72604 5796
rect 72660 5740 75068 5796
rect 75124 5740 75134 5796
rect 30380 5684 30436 5740
rect 50652 5684 50708 5740
rect 30380 5628 35980 5684
rect 36036 5628 36046 5684
rect 36194 5628 36204 5684
rect 36260 5628 37324 5684
rect 37380 5628 37390 5684
rect 42466 5628 42476 5684
rect 42532 5628 50596 5684
rect 50652 5628 51436 5684
rect 51492 5628 52220 5684
rect 52276 5628 52892 5684
rect 52948 5628 53340 5684
rect 53396 5628 53406 5684
rect 56130 5628 56140 5684
rect 56196 5628 56588 5684
rect 56644 5628 56654 5684
rect 62066 5628 62076 5684
rect 62132 5628 63644 5684
rect 63700 5628 65884 5684
rect 65940 5628 65950 5684
rect 67218 5628 67228 5684
rect 67284 5628 68796 5684
rect 68852 5628 73500 5684
rect 73556 5628 73566 5684
rect 50540 5572 50596 5628
rect 13010 5516 13020 5572
rect 13076 5516 13916 5572
rect 13972 5516 14364 5572
rect 14420 5516 14924 5572
rect 14980 5516 16940 5572
rect 16996 5516 18844 5572
rect 18900 5516 18910 5572
rect 46498 5516 46508 5572
rect 46564 5516 47180 5572
rect 47236 5516 48636 5572
rect 48692 5516 48702 5572
rect 50540 5516 51324 5572
rect 51380 5516 51390 5572
rect 54002 5516 54012 5572
rect 54068 5516 54460 5572
rect 54516 5516 55580 5572
rect 55636 5516 55646 5572
rect 72034 5516 72044 5572
rect 72100 5516 73836 5572
rect 73892 5516 73902 5572
rect 10862 5460 10872 5516
rect 10928 5460 10976 5516
rect 11032 5460 11080 5516
rect 11136 5460 11146 5516
rect 30182 5460 30192 5516
rect 30248 5460 30296 5516
rect 30352 5460 30400 5516
rect 30456 5460 30466 5516
rect 49502 5460 49512 5516
rect 49568 5460 49616 5516
rect 49672 5460 49720 5516
rect 49776 5460 49786 5516
rect 68822 5460 68832 5516
rect 68888 5460 68936 5516
rect 68992 5460 69040 5516
rect 69096 5460 69106 5516
rect 12114 5404 12124 5460
rect 12180 5404 26684 5460
rect 26740 5404 26750 5460
rect 27906 5404 27916 5460
rect 27972 5404 29708 5460
rect 29764 5404 29774 5460
rect 38612 5404 42140 5460
rect 42196 5404 42924 5460
rect 42980 5404 42990 5460
rect 46162 5404 46172 5460
rect 46228 5404 46844 5460
rect 46900 5404 47404 5460
rect 47460 5404 47470 5460
rect 55458 5404 55468 5460
rect 55524 5404 56364 5460
rect 56420 5404 56430 5460
rect 6626 5292 6636 5348
rect 6692 5292 8652 5348
rect 8708 5292 9772 5348
rect 9828 5292 9838 5348
rect 18834 5292 18844 5348
rect 18900 5292 34188 5348
rect 34244 5292 34254 5348
rect 35186 5292 35196 5348
rect 35252 5292 37660 5348
rect 37716 5292 37726 5348
rect 38612 5236 38668 5404
rect 40450 5292 40460 5348
rect 40516 5292 46396 5348
rect 46452 5292 47628 5348
rect 47684 5292 47694 5348
rect 47954 5292 47964 5348
rect 48020 5292 48524 5348
rect 48580 5292 51772 5348
rect 51828 5292 51838 5348
rect 56578 5292 56588 5348
rect 56644 5292 60060 5348
rect 60116 5292 60126 5348
rect 66322 5292 66332 5348
rect 66388 5292 67004 5348
rect 67060 5292 67228 5348
rect 74274 5292 74284 5348
rect 74340 5292 75516 5348
rect 75572 5292 75582 5348
rect 76290 5292 76300 5348
rect 76356 5292 76972 5348
rect 77028 5292 77038 5348
rect 67172 5236 67228 5292
rect 7634 5180 7644 5236
rect 7700 5180 8764 5236
rect 8820 5180 8830 5236
rect 12786 5180 12796 5236
rect 12852 5180 13468 5236
rect 13524 5180 14252 5236
rect 14308 5180 16268 5236
rect 16324 5180 16334 5236
rect 16706 5180 16716 5236
rect 16772 5180 19964 5236
rect 20020 5180 20030 5236
rect 21970 5180 21980 5236
rect 22036 5180 25452 5236
rect 25508 5180 25518 5236
rect 28364 5180 29820 5236
rect 29876 5180 29886 5236
rect 30034 5180 30044 5236
rect 30100 5180 32284 5236
rect 32340 5180 32350 5236
rect 34066 5180 34076 5236
rect 34132 5180 35532 5236
rect 35588 5180 35598 5236
rect 37100 5180 38668 5236
rect 39106 5180 39116 5236
rect 39172 5180 40348 5236
rect 40404 5180 40414 5236
rect 44818 5180 44828 5236
rect 44884 5180 45724 5236
rect 45780 5180 50428 5236
rect 50484 5180 50494 5236
rect 53890 5180 53900 5236
rect 53956 5180 57596 5236
rect 57652 5180 57662 5236
rect 60498 5180 60508 5236
rect 60564 5180 61964 5236
rect 62020 5180 62030 5236
rect 65538 5180 65548 5236
rect 65604 5180 66108 5236
rect 66164 5180 66668 5236
rect 66724 5180 66734 5236
rect 67172 5180 69692 5236
rect 69748 5180 69758 5236
rect 73378 5180 73388 5236
rect 73444 5180 77196 5236
rect 77252 5180 77262 5236
rect 28364 5124 28420 5180
rect 32284 5124 32340 5180
rect 37100 5124 37156 5180
rect 1474 5068 1484 5124
rect 1540 5068 3836 5124
rect 3892 5068 4844 5124
rect 4900 5068 4910 5124
rect 9986 5068 9996 5124
rect 10052 5068 10332 5124
rect 10388 5068 10668 5124
rect 10724 5068 10734 5124
rect 14018 5068 14028 5124
rect 14084 5068 15036 5124
rect 15092 5068 15820 5124
rect 15876 5068 15886 5124
rect 16370 5068 16380 5124
rect 16436 5068 17052 5124
rect 17108 5068 17500 5124
rect 17556 5068 17566 5124
rect 17714 5068 17724 5124
rect 17780 5068 18732 5124
rect 18788 5068 19180 5124
rect 19236 5068 28364 5124
rect 28420 5068 28430 5124
rect 29138 5068 29148 5124
rect 29204 5068 30492 5124
rect 30548 5068 30558 5124
rect 32284 5068 34412 5124
rect 34468 5068 34860 5124
rect 34916 5068 34926 5124
rect 36540 5068 37156 5124
rect 38098 5068 38108 5124
rect 38164 5068 38892 5124
rect 38948 5068 38958 5124
rect 39778 5068 39788 5124
rect 39844 5068 41020 5124
rect 41076 5068 41086 5124
rect 48402 5068 48412 5124
rect 48468 5068 49308 5124
rect 49364 5068 50540 5124
rect 50596 5068 50606 5124
rect 53554 5068 53564 5124
rect 53620 5068 55804 5124
rect 55860 5068 55870 5124
rect 56578 5068 56588 5124
rect 56644 5068 58268 5124
rect 58324 5068 58334 5124
rect 59154 5068 59164 5124
rect 59220 5068 59612 5124
rect 59668 5068 65660 5124
rect 65716 5068 65726 5124
rect 66546 5068 66556 5124
rect 66612 5068 67228 5124
rect 36540 5012 36596 5068
rect 67172 5012 67228 5068
rect 70476 5068 73948 5124
rect 74004 5068 74014 5124
rect 75506 5068 75516 5124
rect 75572 5068 78092 5124
rect 78148 5068 78158 5124
rect 16594 4956 16604 5012
rect 16660 4956 17164 5012
rect 17220 4956 17230 5012
rect 18498 4956 18508 5012
rect 18564 4956 19068 5012
rect 19124 4956 19134 5012
rect 19730 4956 19740 5012
rect 19796 4956 23436 5012
rect 23492 4956 24668 5012
rect 24724 4956 24734 5012
rect 24882 4956 24892 5012
rect 24948 4956 25452 5012
rect 25508 4956 27916 5012
rect 27972 4956 27982 5012
rect 28914 4956 28924 5012
rect 28980 4956 30828 5012
rect 30884 4956 36596 5012
rect 36754 4956 36764 5012
rect 36820 4956 39004 5012
rect 39060 4956 39070 5012
rect 40114 4956 40124 5012
rect 40180 4956 41804 5012
rect 41860 4956 41870 5012
rect 44930 4956 44940 5012
rect 44996 4956 45612 5012
rect 45668 4956 45678 5012
rect 50978 4956 50988 5012
rect 51044 4956 53788 5012
rect 53844 4956 53854 5012
rect 54012 4956 54796 5012
rect 54852 4956 54862 5012
rect 55010 4956 55020 5012
rect 55076 4956 55412 5012
rect 55468 4956 55478 5012
rect 55570 4956 55580 5012
rect 55636 4956 57148 5012
rect 57204 4956 60396 5012
rect 60452 4956 64204 5012
rect 64260 4956 64270 5012
rect 67172 4956 67676 5012
rect 67732 4956 69132 5012
rect 69188 4956 69198 5012
rect 54012 4900 54068 4956
rect 70476 4900 70532 5068
rect 74162 4956 74172 5012
rect 74228 4956 74732 5012
rect 74788 4956 75628 5012
rect 75684 4956 77644 5012
rect 77700 4956 77710 5012
rect 3042 4844 3052 4900
rect 3108 4844 3612 4900
rect 3668 4844 3678 4900
rect 19954 4844 19964 4900
rect 20020 4844 31164 4900
rect 31220 4844 31230 4900
rect 31938 4844 31948 4900
rect 32004 4844 32172 4900
rect 32228 4844 33068 4900
rect 33124 4844 33134 4900
rect 37874 4844 37884 4900
rect 37940 4844 39452 4900
rect 39508 4844 40348 4900
rect 40404 4844 40414 4900
rect 41906 4844 41916 4900
rect 41972 4844 42252 4900
rect 42308 4844 42318 4900
rect 43586 4844 43596 4900
rect 43652 4844 44268 4900
rect 44324 4844 45836 4900
rect 45892 4844 45902 4900
rect 46722 4844 46732 4900
rect 46788 4844 54068 4900
rect 54674 4844 54684 4900
rect 54740 4844 55916 4900
rect 55972 4844 57708 4900
rect 57764 4844 58716 4900
rect 58772 4844 58782 4900
rect 58930 4844 58940 4900
rect 58996 4844 61516 4900
rect 61572 4844 61582 4900
rect 61954 4844 61964 4900
rect 62020 4844 63196 4900
rect 63252 4844 63756 4900
rect 63812 4844 63822 4900
rect 64530 4844 64540 4900
rect 64596 4844 65100 4900
rect 65156 4844 66332 4900
rect 66388 4844 66398 4900
rect 66546 4844 66556 4900
rect 66612 4844 70532 4900
rect 72370 4844 72380 4900
rect 72436 4844 74396 4900
rect 74452 4844 74462 4900
rect 5058 4732 5068 4788
rect 5124 4732 18956 4788
rect 19012 4732 19022 4788
rect 23986 4732 23996 4788
rect 24052 4732 24780 4788
rect 24836 4732 24846 4788
rect 26226 4732 26236 4788
rect 26292 4732 26852 4788
rect 26908 4732 26918 4788
rect 27020 4732 27692 4788
rect 27748 4732 28140 4788
rect 28196 4732 30716 4788
rect 30772 4732 31388 4788
rect 31444 4732 31454 4788
rect 31602 4732 31612 4788
rect 31668 4732 39676 4788
rect 39732 4732 39742 4788
rect 40226 4732 40236 4788
rect 40292 4732 41468 4788
rect 41524 4732 41534 4788
rect 42354 4732 42364 4788
rect 42420 4732 43372 4788
rect 43428 4732 43438 4788
rect 43698 4732 43708 4788
rect 43764 4732 44156 4788
rect 44212 4732 44222 4788
rect 44706 4732 44716 4788
rect 44772 4732 46844 4788
rect 46900 4732 46910 4788
rect 51314 4732 51324 4788
rect 51380 4732 53676 4788
rect 53732 4732 53742 4788
rect 54786 4732 54796 4788
rect 54852 4732 58380 4788
rect 58436 4732 58446 4788
rect 63858 4732 63868 4788
rect 63924 4732 64092 4788
rect 64148 4732 66220 4788
rect 66276 4732 66286 4788
rect 66994 4732 67004 4788
rect 67060 4732 68124 4788
rect 68180 4732 68190 4788
rect 68338 4732 68348 4788
rect 68404 4732 73052 4788
rect 73108 4732 73118 4788
rect 20522 4676 20532 4732
rect 20588 4676 20636 4732
rect 20692 4676 20740 4732
rect 20796 4676 20806 4732
rect 27020 4676 27076 4732
rect 39842 4676 39852 4732
rect 39908 4676 39956 4732
rect 40012 4676 40060 4732
rect 40116 4676 40126 4732
rect 43372 4676 43428 4732
rect 44716 4676 44772 4732
rect 59162 4676 59172 4732
rect 59228 4676 59276 4732
rect 59332 4676 59380 4732
rect 59436 4676 59446 4732
rect 78482 4676 78492 4732
rect 78548 4676 78596 4732
rect 78652 4676 78700 4732
rect 78756 4676 78766 4732
rect 25666 4620 25676 4676
rect 25732 4620 27076 4676
rect 27234 4620 27244 4676
rect 27300 4620 27804 4676
rect 27860 4620 39732 4676
rect 39676 4564 39732 4620
rect 40236 4620 41356 4676
rect 41412 4620 41422 4676
rect 41570 4620 41580 4676
rect 41636 4620 42028 4676
rect 42084 4620 42094 4676
rect 43372 4620 44772 4676
rect 46498 4620 46508 4676
rect 46564 4620 48748 4676
rect 48804 4620 48814 4676
rect 51650 4620 51660 4676
rect 51716 4620 52444 4676
rect 52500 4620 53004 4676
rect 53060 4620 53900 4676
rect 53956 4620 55020 4676
rect 55076 4620 55086 4676
rect 55458 4620 55468 4676
rect 55524 4620 56700 4676
rect 56756 4620 56766 4676
rect 61282 4620 61292 4676
rect 61348 4620 63868 4676
rect 63924 4620 67116 4676
rect 67172 4620 69580 4676
rect 69636 4620 69646 4676
rect 40236 4564 40292 4620
rect 46956 4564 47012 4620
rect 2930 4508 2940 4564
rect 2996 4508 3612 4564
rect 3668 4508 3678 4564
rect 11442 4508 11452 4564
rect 11508 4508 14028 4564
rect 14084 4508 14094 4564
rect 16370 4508 16380 4564
rect 16436 4508 19740 4564
rect 19796 4508 20076 4564
rect 20132 4508 20142 4564
rect 24658 4508 24668 4564
rect 24724 4508 26124 4564
rect 26180 4508 26190 4564
rect 31266 4508 31276 4564
rect 31332 4508 31948 4564
rect 32004 4508 34076 4564
rect 34132 4508 34142 4564
rect 37762 4508 37772 4564
rect 37828 4508 39116 4564
rect 39172 4508 39182 4564
rect 39676 4508 40292 4564
rect 40450 4508 40460 4564
rect 40516 4508 41692 4564
rect 41748 4508 42700 4564
rect 42756 4508 42766 4564
rect 44146 4508 44156 4564
rect 44212 4508 46172 4564
rect 46228 4508 46238 4564
rect 46946 4508 46956 4564
rect 47012 4508 47022 4564
rect 47394 4508 47404 4564
rect 47460 4508 50204 4564
rect 50260 4508 55916 4564
rect 55972 4508 55982 4564
rect 56130 4508 56140 4564
rect 56196 4508 56206 4564
rect 56802 4508 56812 4564
rect 56868 4508 58604 4564
rect 58660 4508 58670 4564
rect 59938 4508 59948 4564
rect 60004 4508 61068 4564
rect 61124 4508 61134 4564
rect 61292 4508 63084 4564
rect 63140 4508 64428 4564
rect 64484 4508 66892 4564
rect 66948 4508 66958 4564
rect 68114 4508 68124 4564
rect 68180 4508 70252 4564
rect 70308 4508 72604 4564
rect 72660 4508 72670 4564
rect 73266 4508 73276 4564
rect 73332 4508 74620 4564
rect 74676 4508 74686 4564
rect 56140 4452 56196 4508
rect 1586 4396 1596 4452
rect 1652 4396 3948 4452
rect 4004 4396 4508 4452
rect 4564 4396 4574 4452
rect 6850 4396 6860 4452
rect 6916 4396 18284 4452
rect 18340 4396 18350 4452
rect 23090 4396 23100 4452
rect 23156 4396 24108 4452
rect 24164 4396 24174 4452
rect 26898 4396 26908 4452
rect 26964 4396 29932 4452
rect 29988 4396 30156 4452
rect 30212 4396 31612 4452
rect 31668 4396 31678 4452
rect 33842 4396 33852 4452
rect 33908 4396 35644 4452
rect 35700 4396 36988 4452
rect 37044 4396 37054 4452
rect 38612 4396 39508 4452
rect 40338 4396 40348 4452
rect 40404 4396 42252 4452
rect 42308 4396 42644 4452
rect 38612 4340 38668 4396
rect 8642 4284 8652 4340
rect 8708 4284 11228 4340
rect 11284 4284 12236 4340
rect 12292 4284 12302 4340
rect 20290 4284 20300 4340
rect 20356 4284 21420 4340
rect 21476 4284 21486 4340
rect 24546 4284 24556 4340
rect 24612 4284 25676 4340
rect 25732 4284 25742 4340
rect 26002 4284 26012 4340
rect 26068 4284 27356 4340
rect 27412 4284 27422 4340
rect 32722 4284 32732 4340
rect 32788 4284 33628 4340
rect 33684 4284 33694 4340
rect 33852 4284 38668 4340
rect 39452 4340 39508 4396
rect 40348 4340 40404 4396
rect 42588 4340 42644 4396
rect 43652 4396 47292 4452
rect 47348 4396 47358 4452
rect 49746 4396 49756 4452
rect 49812 4396 53228 4452
rect 53284 4396 53294 4452
rect 53554 4396 53564 4452
rect 53620 4396 54796 4452
rect 54852 4396 54862 4452
rect 55234 4396 55244 4452
rect 55300 4396 56196 4452
rect 43652 4340 43708 4396
rect 56812 4340 56868 4508
rect 61292 4452 61348 4508
rect 73276 4452 73332 4508
rect 58706 4396 58716 4452
rect 58772 4396 59836 4452
rect 59892 4396 59902 4452
rect 60386 4396 60396 4452
rect 60452 4396 61348 4452
rect 62290 4396 62300 4452
rect 62356 4396 63532 4452
rect 63588 4396 68236 4452
rect 68292 4396 68302 4452
rect 69570 4396 69580 4452
rect 69636 4396 73332 4452
rect 39452 4284 40404 4340
rect 41346 4284 41356 4340
rect 41412 4284 41804 4340
rect 41860 4284 42364 4340
rect 42420 4284 42430 4340
rect 42588 4284 43708 4340
rect 44034 4284 44044 4340
rect 44100 4284 50092 4340
rect 50148 4284 50764 4340
rect 50820 4284 50830 4340
rect 51314 4284 51324 4340
rect 51380 4284 52108 4340
rect 52164 4284 52174 4340
rect 53666 4284 53676 4340
rect 53732 4284 55020 4340
rect 55076 4284 55412 4340
rect 55468 4284 55478 4340
rect 55794 4284 55804 4340
rect 55860 4284 56868 4340
rect 58034 4284 58044 4340
rect 58100 4284 61628 4340
rect 61684 4284 61694 4340
rect 67330 4284 67340 4340
rect 67396 4284 70924 4340
rect 70980 4284 72380 4340
rect 72436 4284 72446 4340
rect 33852 4228 33908 4284
rect 50764 4228 50820 4284
rect 9090 4172 9100 4228
rect 9156 4172 11116 4228
rect 11172 4172 12124 4228
rect 12180 4172 12190 4228
rect 13346 4172 13356 4228
rect 13412 4172 14924 4228
rect 14980 4172 14990 4228
rect 20402 4172 20412 4228
rect 20468 4172 21308 4228
rect 21364 4172 26236 4228
rect 26292 4172 26302 4228
rect 31378 4172 31388 4228
rect 31444 4172 33908 4228
rect 34402 4172 34412 4228
rect 34468 4172 36204 4228
rect 36260 4172 36270 4228
rect 37090 4172 37100 4228
rect 37156 4172 38668 4228
rect 38724 4172 39228 4228
rect 39284 4172 39294 4228
rect 50764 4172 51548 4228
rect 51604 4172 51614 4228
rect 53106 4172 53116 4228
rect 53172 4172 54124 4228
rect 54180 4172 54190 4228
rect 54786 4172 54796 4228
rect 54852 4172 55524 4228
rect 56690 4172 56700 4228
rect 56756 4172 57932 4228
rect 57988 4172 59500 4228
rect 59556 4172 60396 4228
rect 60452 4172 60462 4228
rect 63410 4172 63420 4228
rect 63476 4172 68348 4228
rect 68404 4172 68414 4228
rect 54124 4116 54180 4172
rect 11442 4060 11452 4116
rect 11508 4060 12012 4116
rect 12068 4060 15372 4116
rect 15428 4060 15438 4116
rect 24098 4060 24108 4116
rect 24164 4060 27020 4116
rect 27076 4060 27086 4116
rect 54124 4060 55244 4116
rect 55300 4060 55310 4116
rect 0 4004 800 4032
rect 55468 4004 55524 4172
rect 55906 4060 55916 4116
rect 55972 4060 63868 4116
rect 63924 4060 63934 4116
rect 67666 4060 67676 4116
rect 67732 4060 74172 4116
rect 74228 4060 74238 4116
rect 79200 4004 80000 4032
rect 0 3948 1932 4004
rect 1988 3948 1998 4004
rect 20178 3948 20188 4004
rect 20244 3948 21644 4004
rect 21700 3948 23996 4004
rect 24052 3948 27804 4004
rect 27860 3948 27870 4004
rect 40226 3948 40236 4004
rect 40292 3948 47404 4004
rect 47460 3948 47470 4004
rect 55468 3948 55636 4004
rect 57474 3948 57484 4004
rect 57540 3948 57820 4004
rect 57876 3948 58156 4004
rect 58212 3948 59164 4004
rect 59220 3948 59230 4004
rect 75506 3948 75516 4004
rect 75572 3948 80000 4004
rect 0 3920 800 3948
rect 10862 3892 10872 3948
rect 10928 3892 10976 3948
rect 11032 3892 11080 3948
rect 11136 3892 11146 3948
rect 30182 3892 30192 3948
rect 30248 3892 30296 3948
rect 30352 3892 30400 3948
rect 30456 3892 30466 3948
rect 49502 3892 49512 3948
rect 49568 3892 49616 3948
rect 49672 3892 49720 3948
rect 49776 3892 49786 3948
rect 55580 3892 55636 3948
rect 68822 3892 68832 3948
rect 68888 3892 68936 3948
rect 68992 3892 69040 3948
rect 69096 3892 69106 3948
rect 79200 3920 80000 3948
rect 19506 3836 19516 3892
rect 19572 3836 22876 3892
rect 22932 3836 24780 3892
rect 24836 3836 24846 3892
rect 55570 3836 55580 3892
rect 55636 3836 59724 3892
rect 59780 3836 59790 3892
rect 60722 3836 60732 3892
rect 60788 3836 67340 3892
rect 67396 3836 67406 3892
rect 74834 3836 74844 3892
rect 74900 3836 76748 3892
rect 76804 3836 77196 3892
rect 77252 3836 77262 3892
rect 11554 3724 11564 3780
rect 11620 3724 13356 3780
rect 13412 3724 13580 3780
rect 13636 3724 13646 3780
rect 15026 3724 15036 3780
rect 15092 3724 30044 3780
rect 30100 3724 30110 3780
rect 33506 3724 33516 3780
rect 33572 3724 34188 3780
rect 34244 3724 34254 3780
rect 39666 3724 39676 3780
rect 39732 3724 42924 3780
rect 42980 3724 45388 3780
rect 45444 3724 45454 3780
rect 59602 3724 59612 3780
rect 59668 3724 61292 3780
rect 61348 3724 61358 3780
rect 4946 3612 4956 3668
rect 5012 3612 9660 3668
rect 9716 3612 9726 3668
rect 10546 3612 10556 3668
rect 10612 3612 11452 3668
rect 11508 3612 11518 3668
rect 18386 3612 18396 3668
rect 18452 3612 22652 3668
rect 22708 3612 24444 3668
rect 24500 3612 24510 3668
rect 30146 3612 30156 3668
rect 30212 3612 32172 3668
rect 32228 3612 32238 3668
rect 41570 3612 41580 3668
rect 41636 3612 42812 3668
rect 42868 3612 50876 3668
rect 50932 3612 55468 3668
rect 55524 3612 55534 3668
rect 63522 3612 63532 3668
rect 63588 3612 64204 3668
rect 64260 3612 64270 3668
rect 70242 3612 70252 3668
rect 70308 3612 77308 3668
rect 77364 3612 77374 3668
rect 2146 3500 2156 3556
rect 2212 3500 2716 3556
rect 2772 3500 5628 3556
rect 5684 3500 5694 3556
rect 5852 3500 7196 3556
rect 7252 3500 7262 3556
rect 9986 3500 9996 3556
rect 10052 3500 11676 3556
rect 11732 3500 11742 3556
rect 14914 3500 14924 3556
rect 14980 3500 15708 3556
rect 15764 3500 17500 3556
rect 17556 3500 17566 3556
rect 17938 3500 17948 3556
rect 18004 3500 18844 3556
rect 18900 3500 19740 3556
rect 19796 3500 19806 3556
rect 20962 3500 20972 3556
rect 21028 3500 21868 3556
rect 21924 3500 22092 3556
rect 22148 3500 22158 3556
rect 24546 3500 24556 3556
rect 24612 3500 25004 3556
rect 25060 3500 25070 3556
rect 25890 3500 25900 3556
rect 25956 3500 28252 3556
rect 28308 3500 29260 3556
rect 29316 3500 29326 3556
rect 32498 3500 32508 3556
rect 32564 3500 34860 3556
rect 34916 3500 34926 3556
rect 35970 3500 35980 3556
rect 36036 3500 36764 3556
rect 36820 3500 37100 3556
rect 37156 3500 37166 3556
rect 38210 3500 38220 3556
rect 38276 3500 40124 3556
rect 40180 3500 44044 3556
rect 44100 3500 44110 3556
rect 47618 3500 47628 3556
rect 47684 3500 50988 3556
rect 51044 3500 51054 3556
rect 51650 3500 51660 3556
rect 51716 3500 52668 3556
rect 52724 3500 52734 3556
rect 59490 3500 59500 3556
rect 59556 3500 59948 3556
rect 60004 3500 60014 3556
rect 60162 3500 60172 3556
rect 60228 3500 62972 3556
rect 63028 3500 68348 3556
rect 68404 3500 68414 3556
rect 75506 3500 75516 3556
rect 75572 3500 77644 3556
rect 77700 3500 77710 3556
rect 5852 3444 5908 3500
rect 2818 3388 2828 3444
rect 2884 3388 5908 3444
rect 6738 3388 6748 3444
rect 6804 3388 6972 3444
rect 7028 3388 8204 3444
rect 8260 3388 8270 3444
rect 9090 3388 9100 3444
rect 9156 3388 10332 3444
rect 10388 3388 10398 3444
rect 12898 3388 12908 3444
rect 12964 3388 15036 3444
rect 15092 3388 15102 3444
rect 23538 3388 23548 3444
rect 23604 3388 26124 3444
rect 26180 3388 26348 3444
rect 26404 3388 26414 3444
rect 28578 3388 28588 3444
rect 28644 3388 30604 3444
rect 30660 3388 30670 3444
rect 31602 3388 31612 3444
rect 31668 3388 32396 3444
rect 32452 3388 33180 3444
rect 33236 3388 33246 3444
rect 36418 3388 36428 3444
rect 36484 3388 39452 3444
rect 39508 3388 40236 3444
rect 40292 3388 40302 3444
rect 41234 3388 41244 3444
rect 41300 3388 42028 3444
rect 42084 3388 42094 3444
rect 45266 3388 45276 3444
rect 45332 3388 47964 3444
rect 48020 3388 51772 3444
rect 51828 3388 51838 3444
rect 58146 3388 58156 3444
rect 58212 3388 58940 3444
rect 58996 3388 65660 3444
rect 65716 3388 65726 3444
rect 68674 3388 68684 3444
rect 68740 3388 70252 3444
rect 70308 3388 70318 3444
rect 70802 3388 70812 3444
rect 70868 3388 71372 3444
rect 71428 3388 77756 3444
rect 77812 3388 77822 3444
rect 7522 3276 7532 3332
rect 7588 3276 16268 3332
rect 16324 3276 25788 3332
rect 25844 3276 25854 3332
rect 28354 3276 28364 3332
rect 28420 3276 29596 3332
rect 29652 3276 29662 3332
rect 44930 3276 44940 3332
rect 44996 3276 47516 3332
rect 47572 3276 47582 3332
rect 48626 3276 48636 3332
rect 48692 3276 53564 3332
rect 53620 3276 53630 3332
rect 56802 3276 56812 3332
rect 56868 3276 58044 3332
rect 58100 3276 59612 3332
rect 59668 3276 60508 3332
rect 60564 3276 60574 3332
rect 61394 3276 61404 3332
rect 61460 3276 71932 3332
rect 71988 3276 71998 3332
rect 21410 3164 21420 3220
rect 21476 3164 28476 3220
rect 28532 3164 28542 3220
rect 42914 3164 42924 3220
rect 42980 3164 46284 3220
rect 46340 3164 48748 3220
rect 48804 3164 48814 3220
rect 20522 3108 20532 3164
rect 20588 3108 20636 3164
rect 20692 3108 20740 3164
rect 20796 3108 20806 3164
rect 39842 3108 39852 3164
rect 39908 3108 39956 3164
rect 40012 3108 40060 3164
rect 40116 3108 40126 3164
rect 59162 3108 59172 3164
rect 59228 3108 59276 3164
rect 59332 3108 59380 3164
rect 59436 3108 59446 3164
rect 78482 3108 78492 3164
rect 78548 3108 78596 3164
rect 78652 3108 78700 3164
rect 78756 3108 78766 3164
rect 45602 3052 45612 3108
rect 45668 3052 51324 3108
rect 51380 3052 51390 3108
rect 27122 2940 27132 2996
rect 27188 2940 48860 2996
rect 48916 2940 48926 2996
rect 59042 2940 59052 2996
rect 59108 2940 67004 2996
rect 67060 2940 67070 2996
rect 6514 2828 6524 2884
rect 6580 2828 24108 2884
rect 24164 2828 24174 2884
rect 24770 2828 24780 2884
rect 24836 2828 43596 2884
rect 43652 2828 43662 2884
rect 53778 2828 53788 2884
rect 53844 2828 55132 2884
rect 55188 2828 61180 2884
rect 61236 2828 61246 2884
rect 19058 2716 19068 2772
rect 19124 2716 35308 2772
rect 35364 2716 35374 2772
rect 37426 2716 37436 2772
rect 37492 2716 64316 2772
rect 64372 2716 64382 2772
rect 9762 2604 9772 2660
rect 9828 2604 57484 2660
rect 57540 2604 57550 2660
rect 29810 2492 29820 2548
rect 29876 2492 47180 2548
rect 47236 2492 47246 2548
rect 10658 2380 10668 2436
rect 10724 2380 30156 2436
rect 30212 2380 30222 2436
rect 29698 2268 29708 2324
rect 29764 2268 37436 2324
rect 37492 2268 37502 2324
rect 14690 2156 14700 2212
rect 14756 2156 36092 2212
rect 36148 2156 54012 2212
rect 54068 2156 54078 2212
rect 26450 2044 26460 2100
rect 26516 2044 40236 2100
rect 40292 2044 40302 2100
rect 17490 1596 17500 1652
rect 17556 1596 35084 1652
rect 35140 1596 35150 1652
rect 37650 1596 37660 1652
rect 37716 1596 54348 1652
rect 54404 1596 54414 1652
rect 0 1540 800 1568
rect 79200 1540 80000 1568
rect 0 1484 1820 1540
rect 1876 1484 1886 1540
rect 27234 1484 27244 1540
rect 27300 1484 43708 1540
rect 43764 1484 43774 1540
rect 43922 1484 43932 1540
rect 43988 1484 65100 1540
rect 65156 1484 65166 1540
rect 74834 1484 74844 1540
rect 74900 1484 80000 1540
rect 0 1456 800 1484
rect 79200 1456 80000 1484
rect 35298 1372 35308 1428
rect 35364 1372 65436 1428
rect 65492 1372 65502 1428
rect 16482 1260 16492 1316
rect 16548 1260 26908 1316
rect 26964 1260 26974 1316
rect 28802 1260 28812 1316
rect 28868 1260 56588 1316
rect 56644 1260 56654 1316
rect 25218 1148 25228 1204
rect 25284 1148 51212 1204
rect 51268 1148 51278 1204
rect 9538 1036 9548 1092
rect 9604 1036 55356 1092
rect 55412 1036 55422 1092
rect 14466 924 14476 980
rect 14532 924 37828 980
rect 43026 924 43036 980
rect 43092 924 56924 980
rect 56980 924 56990 980
rect 37772 868 37828 924
rect 11778 812 11788 868
rect 11844 812 37548 868
rect 37604 812 37614 868
rect 37772 812 46620 868
rect 46676 812 46686 868
<< via3 >>
rect 10872 36820 10928 36876
rect 10976 36820 11032 36876
rect 11080 36820 11136 36876
rect 30192 36820 30248 36876
rect 30296 36820 30352 36876
rect 30400 36820 30456 36876
rect 49512 36820 49568 36876
rect 49616 36820 49672 36876
rect 49720 36820 49776 36876
rect 68832 36820 68888 36876
rect 68936 36820 68992 36876
rect 69040 36820 69096 36876
rect 20532 36036 20588 36092
rect 20636 36036 20692 36092
rect 20740 36036 20796 36092
rect 39852 36036 39908 36092
rect 39956 36036 40012 36092
rect 40060 36036 40116 36092
rect 59172 36036 59228 36092
rect 59276 36036 59332 36092
rect 59380 36036 59436 36092
rect 78492 36036 78548 36092
rect 78596 36036 78652 36092
rect 78700 36036 78756 36092
rect 10872 35252 10928 35308
rect 10976 35252 11032 35308
rect 11080 35252 11136 35308
rect 30192 35252 30248 35308
rect 30296 35252 30352 35308
rect 30400 35252 30456 35308
rect 49512 35252 49568 35308
rect 49616 35252 49672 35308
rect 49720 35252 49776 35308
rect 68832 35252 68888 35308
rect 68936 35252 68992 35308
rect 69040 35252 69096 35308
rect 31276 35084 31332 35140
rect 31276 34748 31332 34804
rect 20532 34468 20588 34524
rect 20636 34468 20692 34524
rect 20740 34468 20796 34524
rect 39852 34468 39908 34524
rect 39956 34468 40012 34524
rect 40060 34468 40116 34524
rect 59172 34468 59228 34524
rect 59276 34468 59332 34524
rect 59380 34468 59436 34524
rect 78492 34468 78548 34524
rect 78596 34468 78652 34524
rect 78700 34468 78756 34524
rect 10872 33684 10928 33740
rect 10976 33684 11032 33740
rect 11080 33684 11136 33740
rect 30192 33684 30248 33740
rect 30296 33684 30352 33740
rect 30400 33684 30456 33740
rect 49512 33684 49568 33740
rect 49616 33684 49672 33740
rect 49720 33684 49776 33740
rect 68832 33684 68888 33740
rect 68936 33684 68992 33740
rect 69040 33684 69096 33740
rect 20532 32900 20588 32956
rect 20636 32900 20692 32956
rect 20740 32900 20796 32956
rect 39852 32900 39908 32956
rect 39956 32900 40012 32956
rect 40060 32900 40116 32956
rect 59172 32900 59228 32956
rect 59276 32900 59332 32956
rect 59380 32900 59436 32956
rect 78492 32900 78548 32956
rect 78596 32900 78652 32956
rect 78700 32900 78756 32956
rect 10872 32116 10928 32172
rect 10976 32116 11032 32172
rect 11080 32116 11136 32172
rect 30192 32116 30248 32172
rect 30296 32116 30352 32172
rect 30400 32116 30456 32172
rect 49512 32116 49568 32172
rect 49616 32116 49672 32172
rect 49720 32116 49776 32172
rect 68832 32116 68888 32172
rect 68936 32116 68992 32172
rect 69040 32116 69096 32172
rect 20532 31332 20588 31388
rect 20636 31332 20692 31388
rect 20740 31332 20796 31388
rect 39852 31332 39908 31388
rect 39956 31332 40012 31388
rect 40060 31332 40116 31388
rect 59172 31332 59228 31388
rect 59276 31332 59332 31388
rect 59380 31332 59436 31388
rect 78492 31332 78548 31388
rect 78596 31332 78652 31388
rect 78700 31332 78756 31388
rect 55468 30716 55524 30772
rect 10872 30548 10928 30604
rect 10976 30548 11032 30604
rect 11080 30548 11136 30604
rect 30192 30548 30248 30604
rect 30296 30548 30352 30604
rect 30400 30548 30456 30604
rect 49512 30548 49568 30604
rect 49616 30548 49672 30604
rect 49720 30548 49776 30604
rect 68832 30548 68888 30604
rect 68936 30548 68992 30604
rect 69040 30548 69096 30604
rect 55412 30492 55468 30548
rect 20532 29764 20588 29820
rect 20636 29764 20692 29820
rect 20740 29764 20796 29820
rect 39852 29764 39908 29820
rect 39956 29764 40012 29820
rect 40060 29764 40116 29820
rect 59172 29764 59228 29820
rect 59276 29764 59332 29820
rect 59380 29764 59436 29820
rect 78492 29764 78548 29820
rect 78596 29764 78652 29820
rect 78700 29764 78756 29820
rect 10872 28980 10928 29036
rect 10976 28980 11032 29036
rect 11080 28980 11136 29036
rect 30192 28980 30248 29036
rect 30296 28980 30352 29036
rect 30400 28980 30456 29036
rect 49512 28980 49568 29036
rect 49616 28980 49672 29036
rect 49720 28980 49776 29036
rect 68832 28980 68888 29036
rect 68936 28980 68992 29036
rect 69040 28980 69096 29036
rect 77980 28700 78036 28756
rect 77980 28252 78036 28308
rect 20532 28196 20588 28252
rect 20636 28196 20692 28252
rect 20740 28196 20796 28252
rect 39852 28196 39908 28252
rect 39956 28196 40012 28252
rect 40060 28196 40116 28252
rect 59172 28196 59228 28252
rect 59276 28196 59332 28252
rect 59380 28196 59436 28252
rect 78492 28196 78548 28252
rect 78596 28196 78652 28252
rect 78700 28196 78756 28252
rect 46844 27804 46900 27860
rect 46844 27468 46900 27524
rect 10872 27412 10928 27468
rect 10976 27412 11032 27468
rect 11080 27412 11136 27468
rect 30192 27412 30248 27468
rect 30296 27412 30352 27468
rect 30400 27412 30456 27468
rect 49512 27412 49568 27468
rect 49616 27412 49672 27468
rect 49720 27412 49776 27468
rect 68832 27412 68888 27468
rect 68936 27412 68992 27468
rect 69040 27412 69096 27468
rect 53788 27244 53844 27300
rect 20532 26628 20588 26684
rect 20636 26628 20692 26684
rect 20740 26628 20796 26684
rect 39852 26628 39908 26684
rect 39956 26628 40012 26684
rect 40060 26628 40116 26684
rect 59172 26628 59228 26684
rect 59276 26628 59332 26684
rect 59380 26628 59436 26684
rect 78492 26628 78548 26684
rect 78596 26628 78652 26684
rect 78700 26628 78756 26684
rect 53788 26572 53844 26628
rect 10872 25844 10928 25900
rect 10976 25844 11032 25900
rect 11080 25844 11136 25900
rect 30192 25844 30248 25900
rect 30296 25844 30352 25900
rect 30400 25844 30456 25900
rect 49512 25844 49568 25900
rect 49616 25844 49672 25900
rect 49720 25844 49776 25900
rect 68832 25844 68888 25900
rect 68936 25844 68992 25900
rect 69040 25844 69096 25900
rect 20532 25060 20588 25116
rect 20636 25060 20692 25116
rect 20740 25060 20796 25116
rect 39852 25060 39908 25116
rect 39956 25060 40012 25116
rect 40060 25060 40116 25116
rect 59172 25060 59228 25116
rect 59276 25060 59332 25116
rect 59380 25060 59436 25116
rect 78492 25060 78548 25116
rect 78596 25060 78652 25116
rect 78700 25060 78756 25116
rect 10872 24276 10928 24332
rect 10976 24276 11032 24332
rect 11080 24276 11136 24332
rect 30192 24276 30248 24332
rect 30296 24276 30352 24332
rect 30400 24276 30456 24332
rect 49512 24276 49568 24332
rect 49616 24276 49672 24332
rect 49720 24276 49776 24332
rect 68832 24276 68888 24332
rect 68936 24276 68992 24332
rect 69040 24276 69096 24332
rect 15148 24220 15204 24276
rect 60060 23548 60116 23604
rect 20532 23492 20588 23548
rect 20636 23492 20692 23548
rect 20740 23492 20796 23548
rect 39852 23492 39908 23548
rect 39956 23492 40012 23548
rect 40060 23492 40116 23548
rect 59172 23492 59228 23548
rect 59276 23492 59332 23548
rect 59380 23492 59436 23548
rect 78492 23492 78548 23548
rect 78596 23492 78652 23548
rect 78700 23492 78756 23548
rect 60060 23100 60116 23156
rect 10872 22708 10928 22764
rect 10976 22708 11032 22764
rect 11080 22708 11136 22764
rect 30192 22708 30248 22764
rect 30296 22708 30352 22764
rect 30400 22708 30456 22764
rect 49512 22708 49568 22764
rect 49616 22708 49672 22764
rect 49720 22708 49776 22764
rect 68832 22708 68888 22764
rect 68936 22708 68992 22764
rect 69040 22708 69096 22764
rect 65660 21980 65716 22036
rect 20532 21924 20588 21980
rect 20636 21924 20692 21980
rect 20740 21924 20796 21980
rect 39852 21924 39908 21980
rect 39956 21924 40012 21980
rect 40060 21924 40116 21980
rect 59172 21924 59228 21980
rect 59276 21924 59332 21980
rect 59380 21924 59436 21980
rect 78492 21924 78548 21980
rect 78596 21924 78652 21980
rect 78700 21924 78756 21980
rect 51884 21756 51940 21812
rect 51884 21532 51940 21588
rect 65660 21532 65716 21588
rect 10872 21140 10928 21196
rect 10976 21140 11032 21196
rect 11080 21140 11136 21196
rect 30192 21140 30248 21196
rect 30296 21140 30352 21196
rect 30400 21140 30456 21196
rect 49512 21140 49568 21196
rect 49616 21140 49672 21196
rect 49720 21140 49776 21196
rect 68832 21140 68888 21196
rect 68936 21140 68992 21196
rect 69040 21140 69096 21196
rect 15148 20860 15204 20916
rect 20532 20356 20588 20412
rect 20636 20356 20692 20412
rect 20740 20356 20796 20412
rect 39852 20356 39908 20412
rect 39956 20356 40012 20412
rect 40060 20356 40116 20412
rect 59172 20356 59228 20412
rect 59276 20356 59332 20412
rect 59380 20356 59436 20412
rect 78492 20356 78548 20412
rect 78596 20356 78652 20412
rect 78700 20356 78756 20412
rect 10872 19572 10928 19628
rect 10976 19572 11032 19628
rect 11080 19572 11136 19628
rect 30192 19572 30248 19628
rect 30296 19572 30352 19628
rect 30400 19572 30456 19628
rect 49512 19572 49568 19628
rect 49616 19572 49672 19628
rect 49720 19572 49776 19628
rect 18620 19404 18676 19460
rect 68832 19572 68888 19628
rect 68936 19572 68992 19628
rect 69040 19572 69096 19628
rect 20532 18788 20588 18844
rect 20636 18788 20692 18844
rect 20740 18788 20796 18844
rect 39852 18788 39908 18844
rect 39956 18788 40012 18844
rect 40060 18788 40116 18844
rect 59172 18788 59228 18844
rect 59276 18788 59332 18844
rect 59380 18788 59436 18844
rect 78492 18788 78548 18844
rect 78596 18788 78652 18844
rect 78700 18788 78756 18844
rect 10872 18004 10928 18060
rect 10976 18004 11032 18060
rect 11080 18004 11136 18060
rect 30192 18004 30248 18060
rect 30296 18004 30352 18060
rect 30400 18004 30456 18060
rect 49512 18004 49568 18060
rect 49616 18004 49672 18060
rect 49720 18004 49776 18060
rect 68832 18004 68888 18060
rect 68936 18004 68992 18060
rect 69040 18004 69096 18060
rect 20532 17220 20588 17276
rect 20636 17220 20692 17276
rect 20740 17220 20796 17276
rect 39852 17220 39908 17276
rect 39956 17220 40012 17276
rect 40060 17220 40116 17276
rect 59172 17220 59228 17276
rect 59276 17220 59332 17276
rect 59380 17220 59436 17276
rect 78492 17220 78548 17276
rect 78596 17220 78652 17276
rect 78700 17220 78756 17276
rect 18620 16604 18676 16660
rect 10872 16436 10928 16492
rect 10976 16436 11032 16492
rect 11080 16436 11136 16492
rect 30192 16436 30248 16492
rect 30296 16436 30352 16492
rect 30400 16436 30456 16492
rect 49512 16436 49568 16492
rect 49616 16436 49672 16492
rect 49720 16436 49776 16492
rect 68832 16436 68888 16492
rect 68936 16436 68992 16492
rect 69040 16436 69096 16492
rect 20532 15652 20588 15708
rect 20636 15652 20692 15708
rect 20740 15652 20796 15708
rect 32172 16044 32228 16100
rect 39852 15652 39908 15708
rect 39956 15652 40012 15708
rect 40060 15652 40116 15708
rect 59172 15652 59228 15708
rect 59276 15652 59332 15708
rect 59380 15652 59436 15708
rect 78492 15652 78548 15708
rect 78596 15652 78652 15708
rect 78700 15652 78756 15708
rect 37772 15596 37828 15652
rect 32172 15148 32228 15204
rect 37772 15148 37828 15204
rect 55356 15148 55412 15204
rect 10872 14868 10928 14924
rect 10976 14868 11032 14924
rect 11080 14868 11136 14924
rect 30192 14868 30248 14924
rect 30296 14868 30352 14924
rect 30400 14868 30456 14924
rect 49512 14868 49568 14924
rect 49616 14868 49672 14924
rect 49720 14868 49776 14924
rect 68832 14868 68888 14924
rect 68936 14868 68992 14924
rect 69040 14868 69096 14924
rect 20972 14476 21028 14532
rect 20532 14084 20588 14140
rect 20636 14084 20692 14140
rect 20740 14084 20796 14140
rect 39852 14084 39908 14140
rect 39956 14084 40012 14140
rect 40060 14084 40116 14140
rect 59172 14084 59228 14140
rect 59276 14084 59332 14140
rect 59380 14084 59436 14140
rect 78492 14084 78548 14140
rect 78596 14084 78652 14140
rect 78700 14084 78756 14140
rect 20972 13580 21028 13636
rect 18172 13468 18228 13524
rect 55356 13356 55412 13412
rect 10872 13300 10928 13356
rect 10976 13300 11032 13356
rect 11080 13300 11136 13356
rect 30192 13300 30248 13356
rect 30296 13300 30352 13356
rect 30400 13300 30456 13356
rect 49512 13300 49568 13356
rect 49616 13300 49672 13356
rect 49720 13300 49776 13356
rect 68832 13300 68888 13356
rect 68936 13300 68992 13356
rect 69040 13300 69096 13356
rect 18172 13020 18228 13076
rect 20532 12516 20588 12572
rect 20636 12516 20692 12572
rect 20740 12516 20796 12572
rect 39852 12516 39908 12572
rect 39956 12516 40012 12572
rect 40060 12516 40116 12572
rect 59172 12516 59228 12572
rect 59276 12516 59332 12572
rect 59380 12516 59436 12572
rect 78492 12516 78548 12572
rect 78596 12516 78652 12572
rect 78700 12516 78756 12572
rect 43596 12124 43652 12180
rect 10872 11732 10928 11788
rect 10976 11732 11032 11788
rect 11080 11732 11136 11788
rect 30192 11732 30248 11788
rect 30296 11732 30352 11788
rect 30400 11732 30456 11788
rect 49512 11732 49568 11788
rect 49616 11732 49672 11788
rect 49720 11732 49776 11788
rect 68832 11732 68888 11788
rect 68936 11732 68992 11788
rect 69040 11732 69096 11788
rect 43596 11676 43652 11732
rect 20532 10948 20588 11004
rect 20636 10948 20692 11004
rect 20740 10948 20796 11004
rect 39852 10948 39908 11004
rect 39956 10948 40012 11004
rect 40060 10948 40116 11004
rect 59172 10948 59228 11004
rect 59276 10948 59332 11004
rect 59380 10948 59436 11004
rect 78492 10948 78548 11004
rect 78596 10948 78652 11004
rect 78700 10948 78756 11004
rect 10872 10164 10928 10220
rect 10976 10164 11032 10220
rect 11080 10164 11136 10220
rect 30192 10164 30248 10220
rect 30296 10164 30352 10220
rect 30400 10164 30456 10220
rect 49512 10164 49568 10220
rect 49616 10164 49672 10220
rect 49720 10164 49776 10220
rect 68832 10164 68888 10220
rect 68936 10164 68992 10220
rect 69040 10164 69096 10220
rect 17948 10108 18004 10164
rect 24220 9996 24276 10052
rect 61516 9884 61572 9940
rect 15260 9660 15316 9716
rect 24220 9436 24276 9492
rect 20532 9380 20588 9436
rect 20636 9380 20692 9436
rect 20740 9380 20796 9436
rect 39852 9380 39908 9436
rect 39956 9380 40012 9436
rect 40060 9380 40116 9436
rect 59172 9380 59228 9436
rect 59276 9380 59332 9436
rect 59380 9380 59436 9436
rect 78492 9380 78548 9436
rect 78596 9380 78652 9436
rect 78700 9380 78756 9436
rect 17948 9324 18004 9380
rect 15260 9212 15316 9268
rect 61516 9100 61572 9156
rect 10872 8596 10928 8652
rect 10976 8596 11032 8652
rect 11080 8596 11136 8652
rect 30192 8596 30248 8652
rect 30296 8596 30352 8652
rect 30400 8596 30456 8652
rect 49512 8596 49568 8652
rect 49616 8596 49672 8652
rect 49720 8596 49776 8652
rect 68832 8596 68888 8652
rect 68936 8596 68992 8652
rect 69040 8596 69096 8652
rect 20532 7812 20588 7868
rect 20636 7812 20692 7868
rect 20740 7812 20796 7868
rect 39852 7812 39908 7868
rect 39956 7812 40012 7868
rect 40060 7812 40116 7868
rect 59172 7812 59228 7868
rect 59276 7812 59332 7868
rect 59380 7812 59436 7868
rect 78492 7812 78548 7868
rect 78596 7812 78652 7868
rect 78700 7812 78756 7868
rect 10872 7028 10928 7084
rect 10976 7028 11032 7084
rect 11080 7028 11136 7084
rect 30192 7028 30248 7084
rect 30296 7028 30352 7084
rect 30400 7028 30456 7084
rect 49512 7028 49568 7084
rect 49616 7028 49672 7084
rect 49720 7028 49776 7084
rect 68832 7028 68888 7084
rect 68936 7028 68992 7084
rect 69040 7028 69096 7084
rect 63868 6860 63924 6916
rect 55804 6636 55860 6692
rect 67228 6524 67284 6580
rect 20532 6244 20588 6300
rect 20636 6244 20692 6300
rect 20740 6244 20796 6300
rect 39852 6244 39908 6300
rect 39956 6244 40012 6300
rect 40060 6244 40116 6300
rect 67340 6300 67396 6356
rect 59172 6244 59228 6300
rect 59276 6244 59332 6300
rect 59380 6244 59436 6300
rect 78492 6244 78548 6300
rect 78596 6244 78652 6300
rect 78700 6244 78756 6300
rect 67228 6188 67284 6244
rect 55916 6076 55972 6132
rect 67452 6076 67508 6132
rect 56252 5964 56308 6020
rect 10872 5460 10928 5516
rect 10976 5460 11032 5516
rect 11080 5460 11136 5516
rect 30192 5460 30248 5516
rect 30296 5460 30352 5516
rect 30400 5460 30456 5516
rect 49512 5460 49568 5516
rect 49616 5460 49672 5516
rect 49720 5460 49776 5516
rect 68832 5460 68888 5516
rect 68936 5460 68992 5516
rect 69040 5460 69096 5516
rect 55804 5068 55860 5124
rect 55412 4956 55468 5012
rect 26852 4732 26908 4788
rect 31612 4732 31668 4788
rect 39676 4732 39732 4788
rect 20532 4676 20588 4732
rect 20636 4676 20692 4732
rect 20740 4676 20796 4732
rect 39852 4676 39908 4732
rect 39956 4676 40012 4732
rect 40060 4676 40116 4732
rect 59172 4676 59228 4732
rect 59276 4676 59332 4732
rect 59380 4676 59436 4732
rect 78492 4676 78548 4732
rect 78596 4676 78652 4732
rect 78700 4676 78756 4732
rect 55468 4620 55524 4676
rect 63868 4620 63924 4676
rect 55916 4508 55972 4564
rect 26908 4396 26964 4452
rect 31612 4396 31668 4452
rect 55412 4284 55468 4340
rect 55804 4284 55860 4340
rect 55916 4060 55972 4116
rect 10872 3892 10928 3948
rect 10976 3892 11032 3948
rect 11080 3892 11136 3948
rect 30192 3892 30248 3948
rect 30296 3892 30352 3948
rect 30400 3892 30456 3948
rect 49512 3892 49568 3948
rect 49616 3892 49672 3948
rect 49720 3892 49776 3948
rect 68832 3892 68888 3948
rect 68936 3892 68992 3948
rect 69040 3892 69096 3948
rect 39676 3724 39732 3780
rect 20532 3108 20588 3164
rect 20636 3108 20692 3164
rect 20740 3108 20796 3164
rect 39852 3108 39908 3164
rect 39956 3108 40012 3164
rect 40060 3108 40116 3164
rect 59172 3108 59228 3164
rect 59276 3108 59332 3164
rect 59380 3108 59436 3164
rect 78492 3108 78548 3164
rect 78596 3108 78652 3164
rect 78700 3108 78756 3164
<< metal4 >>
rect 10844 36876 11164 36908
rect 10844 36820 10872 36876
rect 10928 36820 10976 36876
rect 11032 36820 11080 36876
rect 11136 36820 11164 36876
rect 10844 35308 11164 36820
rect 10844 35252 10872 35308
rect 10928 35252 10976 35308
rect 11032 35252 11080 35308
rect 11136 35252 11164 35308
rect 10844 33740 11164 35252
rect 10844 33684 10872 33740
rect 10928 33684 10976 33740
rect 11032 33684 11080 33740
rect 11136 33684 11164 33740
rect 10844 32172 11164 33684
rect 10844 32116 10872 32172
rect 10928 32116 10976 32172
rect 11032 32116 11080 32172
rect 11136 32116 11164 32172
rect 10844 30604 11164 32116
rect 10844 30548 10872 30604
rect 10928 30548 10976 30604
rect 11032 30548 11080 30604
rect 11136 30548 11164 30604
rect 10844 29036 11164 30548
rect 10844 28980 10872 29036
rect 10928 28980 10976 29036
rect 11032 28980 11080 29036
rect 11136 28980 11164 29036
rect 10844 27468 11164 28980
rect 10844 27412 10872 27468
rect 10928 27412 10976 27468
rect 11032 27412 11080 27468
rect 11136 27412 11164 27468
rect 10844 25900 11164 27412
rect 10844 25844 10872 25900
rect 10928 25844 10976 25900
rect 11032 25844 11080 25900
rect 11136 25844 11164 25900
rect 10844 24332 11164 25844
rect 10844 24276 10872 24332
rect 10928 24276 10976 24332
rect 11032 24276 11080 24332
rect 11136 24276 11164 24332
rect 20504 36092 20824 36908
rect 20504 36036 20532 36092
rect 20588 36036 20636 36092
rect 20692 36036 20740 36092
rect 20796 36036 20824 36092
rect 20504 34524 20824 36036
rect 20504 34468 20532 34524
rect 20588 34468 20636 34524
rect 20692 34468 20740 34524
rect 20796 34468 20824 34524
rect 20504 32956 20824 34468
rect 20504 32900 20532 32956
rect 20588 32900 20636 32956
rect 20692 32900 20740 32956
rect 20796 32900 20824 32956
rect 20504 31388 20824 32900
rect 20504 31332 20532 31388
rect 20588 31332 20636 31388
rect 20692 31332 20740 31388
rect 20796 31332 20824 31388
rect 20504 29820 20824 31332
rect 20504 29764 20532 29820
rect 20588 29764 20636 29820
rect 20692 29764 20740 29820
rect 20796 29764 20824 29820
rect 20504 28252 20824 29764
rect 20504 28196 20532 28252
rect 20588 28196 20636 28252
rect 20692 28196 20740 28252
rect 20796 28196 20824 28252
rect 20504 26684 20824 28196
rect 20504 26628 20532 26684
rect 20588 26628 20636 26684
rect 20692 26628 20740 26684
rect 20796 26628 20824 26684
rect 20504 25116 20824 26628
rect 20504 25060 20532 25116
rect 20588 25060 20636 25116
rect 20692 25060 20740 25116
rect 20796 25060 20824 25116
rect 10844 22764 11164 24276
rect 10844 22708 10872 22764
rect 10928 22708 10976 22764
rect 11032 22708 11080 22764
rect 11136 22708 11164 22764
rect 10844 21196 11164 22708
rect 10844 21140 10872 21196
rect 10928 21140 10976 21196
rect 11032 21140 11080 21196
rect 11136 21140 11164 21196
rect 10844 19628 11164 21140
rect 15148 24276 15204 24286
rect 15148 20916 15204 24220
rect 15148 20850 15204 20860
rect 20504 23548 20824 25060
rect 20504 23492 20532 23548
rect 20588 23492 20636 23548
rect 20692 23492 20740 23548
rect 20796 23492 20824 23548
rect 20504 21980 20824 23492
rect 20504 21924 20532 21980
rect 20588 21924 20636 21980
rect 20692 21924 20740 21980
rect 20796 21924 20824 21980
rect 10844 19572 10872 19628
rect 10928 19572 10976 19628
rect 11032 19572 11080 19628
rect 11136 19572 11164 19628
rect 10844 18060 11164 19572
rect 20504 20412 20824 21924
rect 20504 20356 20532 20412
rect 20588 20356 20636 20412
rect 20692 20356 20740 20412
rect 20796 20356 20824 20412
rect 10844 18004 10872 18060
rect 10928 18004 10976 18060
rect 11032 18004 11080 18060
rect 11136 18004 11164 18060
rect 10844 16492 11164 18004
rect 18620 19460 18676 19470
rect 18620 16660 18676 19404
rect 18620 16594 18676 16604
rect 20504 18844 20824 20356
rect 20504 18788 20532 18844
rect 20588 18788 20636 18844
rect 20692 18788 20740 18844
rect 20796 18788 20824 18844
rect 20504 17276 20824 18788
rect 20504 17220 20532 17276
rect 20588 17220 20636 17276
rect 20692 17220 20740 17276
rect 20796 17220 20824 17276
rect 10844 16436 10872 16492
rect 10928 16436 10976 16492
rect 11032 16436 11080 16492
rect 11136 16436 11164 16492
rect 10844 14924 11164 16436
rect 10844 14868 10872 14924
rect 10928 14868 10976 14924
rect 11032 14868 11080 14924
rect 11136 14868 11164 14924
rect 10844 13356 11164 14868
rect 20504 15708 20824 17220
rect 20504 15652 20532 15708
rect 20588 15652 20636 15708
rect 20692 15652 20740 15708
rect 20796 15652 20824 15708
rect 20504 14140 20824 15652
rect 30164 36876 30484 36908
rect 30164 36820 30192 36876
rect 30248 36820 30296 36876
rect 30352 36820 30400 36876
rect 30456 36820 30484 36876
rect 30164 35308 30484 36820
rect 30164 35252 30192 35308
rect 30248 35252 30296 35308
rect 30352 35252 30400 35308
rect 30456 35252 30484 35308
rect 30164 33740 30484 35252
rect 39824 36092 40144 36908
rect 39824 36036 39852 36092
rect 39908 36036 39956 36092
rect 40012 36036 40060 36092
rect 40116 36036 40144 36092
rect 31276 35140 31332 35150
rect 31276 34804 31332 35084
rect 31276 34738 31332 34748
rect 30164 33684 30192 33740
rect 30248 33684 30296 33740
rect 30352 33684 30400 33740
rect 30456 33684 30484 33740
rect 30164 32172 30484 33684
rect 30164 32116 30192 32172
rect 30248 32116 30296 32172
rect 30352 32116 30400 32172
rect 30456 32116 30484 32172
rect 30164 30604 30484 32116
rect 30164 30548 30192 30604
rect 30248 30548 30296 30604
rect 30352 30548 30400 30604
rect 30456 30548 30484 30604
rect 30164 29036 30484 30548
rect 30164 28980 30192 29036
rect 30248 28980 30296 29036
rect 30352 28980 30400 29036
rect 30456 28980 30484 29036
rect 30164 27468 30484 28980
rect 30164 27412 30192 27468
rect 30248 27412 30296 27468
rect 30352 27412 30400 27468
rect 30456 27412 30484 27468
rect 30164 25900 30484 27412
rect 30164 25844 30192 25900
rect 30248 25844 30296 25900
rect 30352 25844 30400 25900
rect 30456 25844 30484 25900
rect 30164 24332 30484 25844
rect 30164 24276 30192 24332
rect 30248 24276 30296 24332
rect 30352 24276 30400 24332
rect 30456 24276 30484 24332
rect 30164 22764 30484 24276
rect 30164 22708 30192 22764
rect 30248 22708 30296 22764
rect 30352 22708 30400 22764
rect 30456 22708 30484 22764
rect 30164 21196 30484 22708
rect 30164 21140 30192 21196
rect 30248 21140 30296 21196
rect 30352 21140 30400 21196
rect 30456 21140 30484 21196
rect 30164 19628 30484 21140
rect 30164 19572 30192 19628
rect 30248 19572 30296 19628
rect 30352 19572 30400 19628
rect 30456 19572 30484 19628
rect 30164 18060 30484 19572
rect 30164 18004 30192 18060
rect 30248 18004 30296 18060
rect 30352 18004 30400 18060
rect 30456 18004 30484 18060
rect 30164 16492 30484 18004
rect 30164 16436 30192 16492
rect 30248 16436 30296 16492
rect 30352 16436 30400 16492
rect 30456 16436 30484 16492
rect 30164 14924 30484 16436
rect 39824 34524 40144 36036
rect 39824 34468 39852 34524
rect 39908 34468 39956 34524
rect 40012 34468 40060 34524
rect 40116 34468 40144 34524
rect 39824 32956 40144 34468
rect 39824 32900 39852 32956
rect 39908 32900 39956 32956
rect 40012 32900 40060 32956
rect 40116 32900 40144 32956
rect 39824 31388 40144 32900
rect 39824 31332 39852 31388
rect 39908 31332 39956 31388
rect 40012 31332 40060 31388
rect 40116 31332 40144 31388
rect 39824 29820 40144 31332
rect 39824 29764 39852 29820
rect 39908 29764 39956 29820
rect 40012 29764 40060 29820
rect 40116 29764 40144 29820
rect 39824 28252 40144 29764
rect 39824 28196 39852 28252
rect 39908 28196 39956 28252
rect 40012 28196 40060 28252
rect 40116 28196 40144 28252
rect 39824 26684 40144 28196
rect 49484 36876 49804 36908
rect 49484 36820 49512 36876
rect 49568 36820 49616 36876
rect 49672 36820 49720 36876
rect 49776 36820 49804 36876
rect 49484 35308 49804 36820
rect 49484 35252 49512 35308
rect 49568 35252 49616 35308
rect 49672 35252 49720 35308
rect 49776 35252 49804 35308
rect 49484 33740 49804 35252
rect 49484 33684 49512 33740
rect 49568 33684 49616 33740
rect 49672 33684 49720 33740
rect 49776 33684 49804 33740
rect 49484 32172 49804 33684
rect 49484 32116 49512 32172
rect 49568 32116 49616 32172
rect 49672 32116 49720 32172
rect 49776 32116 49804 32172
rect 49484 30604 49804 32116
rect 59144 36092 59464 36908
rect 59144 36036 59172 36092
rect 59228 36036 59276 36092
rect 59332 36036 59380 36092
rect 59436 36036 59464 36092
rect 59144 34524 59464 36036
rect 59144 34468 59172 34524
rect 59228 34468 59276 34524
rect 59332 34468 59380 34524
rect 59436 34468 59464 34524
rect 59144 32956 59464 34468
rect 59144 32900 59172 32956
rect 59228 32900 59276 32956
rect 59332 32900 59380 32956
rect 59436 32900 59464 32956
rect 59144 31388 59464 32900
rect 59144 31332 59172 31388
rect 59228 31332 59276 31388
rect 59332 31332 59380 31388
rect 59436 31332 59464 31388
rect 49484 30548 49512 30604
rect 49568 30548 49616 30604
rect 49672 30548 49720 30604
rect 49776 30548 49804 30604
rect 55468 30772 55524 30782
rect 55468 30558 55524 30716
rect 49484 29036 49804 30548
rect 55412 30548 55524 30558
rect 55468 30492 55524 30548
rect 55412 30482 55468 30492
rect 49484 28980 49512 29036
rect 49568 28980 49616 29036
rect 49672 28980 49720 29036
rect 49776 28980 49804 29036
rect 46844 27860 46900 27870
rect 46844 27524 46900 27804
rect 46844 27458 46900 27468
rect 49484 27468 49804 28980
rect 39824 26628 39852 26684
rect 39908 26628 39956 26684
rect 40012 26628 40060 26684
rect 40116 26628 40144 26684
rect 39824 25116 40144 26628
rect 39824 25060 39852 25116
rect 39908 25060 39956 25116
rect 40012 25060 40060 25116
rect 40116 25060 40144 25116
rect 39824 23548 40144 25060
rect 39824 23492 39852 23548
rect 39908 23492 39956 23548
rect 40012 23492 40060 23548
rect 40116 23492 40144 23548
rect 39824 21980 40144 23492
rect 39824 21924 39852 21980
rect 39908 21924 39956 21980
rect 40012 21924 40060 21980
rect 40116 21924 40144 21980
rect 39824 20412 40144 21924
rect 39824 20356 39852 20412
rect 39908 20356 39956 20412
rect 40012 20356 40060 20412
rect 40116 20356 40144 20412
rect 39824 18844 40144 20356
rect 39824 18788 39852 18844
rect 39908 18788 39956 18844
rect 40012 18788 40060 18844
rect 40116 18788 40144 18844
rect 39824 17276 40144 18788
rect 39824 17220 39852 17276
rect 39908 17220 39956 17276
rect 40012 17220 40060 17276
rect 40116 17220 40144 17276
rect 32172 16100 32228 16110
rect 32172 15204 32228 16044
rect 39824 15708 40144 17220
rect 32172 15138 32228 15148
rect 37772 15652 37828 15662
rect 37772 15204 37828 15596
rect 37772 15138 37828 15148
rect 39824 15652 39852 15708
rect 39908 15652 39956 15708
rect 40012 15652 40060 15708
rect 40116 15652 40144 15708
rect 30164 14868 30192 14924
rect 30248 14868 30296 14924
rect 30352 14868 30400 14924
rect 30456 14868 30484 14924
rect 20504 14084 20532 14140
rect 20588 14084 20636 14140
rect 20692 14084 20740 14140
rect 20796 14084 20824 14140
rect 10844 13300 10872 13356
rect 10928 13300 10976 13356
rect 11032 13300 11080 13356
rect 11136 13300 11164 13356
rect 10844 11788 11164 13300
rect 18172 13524 18228 13534
rect 18172 13076 18228 13468
rect 18172 13010 18228 13020
rect 10844 11732 10872 11788
rect 10928 11732 10976 11788
rect 11032 11732 11080 11788
rect 11136 11732 11164 11788
rect 10844 10220 11164 11732
rect 10844 10164 10872 10220
rect 10928 10164 10976 10220
rect 11032 10164 11080 10220
rect 11136 10164 11164 10220
rect 20504 12572 20824 14084
rect 20972 14532 21028 14542
rect 20972 13636 21028 14476
rect 20972 13570 21028 13580
rect 20504 12516 20532 12572
rect 20588 12516 20636 12572
rect 20692 12516 20740 12572
rect 20796 12516 20824 12572
rect 20504 11004 20824 12516
rect 20504 10948 20532 11004
rect 20588 10948 20636 11004
rect 20692 10948 20740 11004
rect 20796 10948 20824 11004
rect 10844 8652 11164 10164
rect 17948 10164 18004 10174
rect 15260 9716 15316 9726
rect 15260 9268 15316 9660
rect 17948 9380 18004 10108
rect 17948 9314 18004 9324
rect 20504 9436 20824 10948
rect 30164 13356 30484 14868
rect 30164 13300 30192 13356
rect 30248 13300 30296 13356
rect 30352 13300 30400 13356
rect 30456 13300 30484 13356
rect 30164 11788 30484 13300
rect 30164 11732 30192 11788
rect 30248 11732 30296 11788
rect 30352 11732 30400 11788
rect 30456 11732 30484 11788
rect 30164 10220 30484 11732
rect 30164 10164 30192 10220
rect 30248 10164 30296 10220
rect 30352 10164 30400 10220
rect 30456 10164 30484 10220
rect 20504 9380 20532 9436
rect 20588 9380 20636 9436
rect 20692 9380 20740 9436
rect 20796 9380 20824 9436
rect 24220 10052 24276 10062
rect 24220 9492 24276 9996
rect 24220 9426 24276 9436
rect 15260 9202 15316 9212
rect 10844 8596 10872 8652
rect 10928 8596 10976 8652
rect 11032 8596 11080 8652
rect 11136 8596 11164 8652
rect 10844 7084 11164 8596
rect 10844 7028 10872 7084
rect 10928 7028 10976 7084
rect 11032 7028 11080 7084
rect 11136 7028 11164 7084
rect 10844 5516 11164 7028
rect 10844 5460 10872 5516
rect 10928 5460 10976 5516
rect 11032 5460 11080 5516
rect 11136 5460 11164 5516
rect 10844 3948 11164 5460
rect 10844 3892 10872 3948
rect 10928 3892 10976 3948
rect 11032 3892 11080 3948
rect 11136 3892 11164 3948
rect 10844 3076 11164 3892
rect 20504 7868 20824 9380
rect 20504 7812 20532 7868
rect 20588 7812 20636 7868
rect 20692 7812 20740 7868
rect 20796 7812 20824 7868
rect 20504 6300 20824 7812
rect 20504 6244 20532 6300
rect 20588 6244 20636 6300
rect 20692 6244 20740 6300
rect 20796 6244 20824 6300
rect 20504 4732 20824 6244
rect 30164 8652 30484 10164
rect 30164 8596 30192 8652
rect 30248 8596 30296 8652
rect 30352 8596 30400 8652
rect 30456 8596 30484 8652
rect 30164 7084 30484 8596
rect 30164 7028 30192 7084
rect 30248 7028 30296 7084
rect 30352 7028 30400 7084
rect 30456 7028 30484 7084
rect 30164 5516 30484 7028
rect 30164 5460 30192 5516
rect 30248 5460 30296 5516
rect 30352 5460 30400 5516
rect 30456 5460 30484 5516
rect 20504 4676 20532 4732
rect 20588 4676 20636 4732
rect 20692 4676 20740 4732
rect 20796 4676 20824 4732
rect 26852 4788 26908 4798
rect 26908 4732 26964 4788
rect 26852 4722 26964 4732
rect 20504 3164 20824 4676
rect 26908 4452 26964 4722
rect 26908 4386 26964 4396
rect 20504 3108 20532 3164
rect 20588 3108 20636 3164
rect 20692 3108 20740 3164
rect 20796 3108 20824 3164
rect 20504 3076 20824 3108
rect 30164 3948 30484 5460
rect 39824 14140 40144 15652
rect 39824 14084 39852 14140
rect 39908 14084 39956 14140
rect 40012 14084 40060 14140
rect 40116 14084 40144 14140
rect 39824 12572 40144 14084
rect 39824 12516 39852 12572
rect 39908 12516 39956 12572
rect 40012 12516 40060 12572
rect 40116 12516 40144 12572
rect 39824 11004 40144 12516
rect 49484 27412 49512 27468
rect 49568 27412 49616 27468
rect 49672 27412 49720 27468
rect 49776 27412 49804 27468
rect 49484 25900 49804 27412
rect 59144 29820 59464 31332
rect 59144 29764 59172 29820
rect 59228 29764 59276 29820
rect 59332 29764 59380 29820
rect 59436 29764 59464 29820
rect 59144 28252 59464 29764
rect 59144 28196 59172 28252
rect 59228 28196 59276 28252
rect 59332 28196 59380 28252
rect 59436 28196 59464 28252
rect 53788 27300 53844 27310
rect 53788 26628 53844 27244
rect 53788 26562 53844 26572
rect 59144 26684 59464 28196
rect 59144 26628 59172 26684
rect 59228 26628 59276 26684
rect 59332 26628 59380 26684
rect 59436 26628 59464 26684
rect 49484 25844 49512 25900
rect 49568 25844 49616 25900
rect 49672 25844 49720 25900
rect 49776 25844 49804 25900
rect 49484 24332 49804 25844
rect 49484 24276 49512 24332
rect 49568 24276 49616 24332
rect 49672 24276 49720 24332
rect 49776 24276 49804 24332
rect 49484 22764 49804 24276
rect 49484 22708 49512 22764
rect 49568 22708 49616 22764
rect 49672 22708 49720 22764
rect 49776 22708 49804 22764
rect 49484 21196 49804 22708
rect 59144 25116 59464 26628
rect 59144 25060 59172 25116
rect 59228 25060 59276 25116
rect 59332 25060 59380 25116
rect 59436 25060 59464 25116
rect 59144 23548 59464 25060
rect 68804 36876 69124 36908
rect 68804 36820 68832 36876
rect 68888 36820 68936 36876
rect 68992 36820 69040 36876
rect 69096 36820 69124 36876
rect 68804 35308 69124 36820
rect 68804 35252 68832 35308
rect 68888 35252 68936 35308
rect 68992 35252 69040 35308
rect 69096 35252 69124 35308
rect 68804 33740 69124 35252
rect 68804 33684 68832 33740
rect 68888 33684 68936 33740
rect 68992 33684 69040 33740
rect 69096 33684 69124 33740
rect 68804 32172 69124 33684
rect 68804 32116 68832 32172
rect 68888 32116 68936 32172
rect 68992 32116 69040 32172
rect 69096 32116 69124 32172
rect 68804 30604 69124 32116
rect 68804 30548 68832 30604
rect 68888 30548 68936 30604
rect 68992 30548 69040 30604
rect 69096 30548 69124 30604
rect 68804 29036 69124 30548
rect 68804 28980 68832 29036
rect 68888 28980 68936 29036
rect 68992 28980 69040 29036
rect 69096 28980 69124 29036
rect 68804 27468 69124 28980
rect 78464 36092 78784 36908
rect 78464 36036 78492 36092
rect 78548 36036 78596 36092
rect 78652 36036 78700 36092
rect 78756 36036 78784 36092
rect 78464 34524 78784 36036
rect 78464 34468 78492 34524
rect 78548 34468 78596 34524
rect 78652 34468 78700 34524
rect 78756 34468 78784 34524
rect 78464 32956 78784 34468
rect 78464 32900 78492 32956
rect 78548 32900 78596 32956
rect 78652 32900 78700 32956
rect 78756 32900 78784 32956
rect 78464 31388 78784 32900
rect 78464 31332 78492 31388
rect 78548 31332 78596 31388
rect 78652 31332 78700 31388
rect 78756 31332 78784 31388
rect 78464 29820 78784 31332
rect 78464 29764 78492 29820
rect 78548 29764 78596 29820
rect 78652 29764 78700 29820
rect 78756 29764 78784 29820
rect 77980 28756 78036 28766
rect 77980 28308 78036 28700
rect 77980 28242 78036 28252
rect 78464 28252 78784 29764
rect 68804 27412 68832 27468
rect 68888 27412 68936 27468
rect 68992 27412 69040 27468
rect 69096 27412 69124 27468
rect 68804 25900 69124 27412
rect 68804 25844 68832 25900
rect 68888 25844 68936 25900
rect 68992 25844 69040 25900
rect 69096 25844 69124 25900
rect 68804 24332 69124 25844
rect 68804 24276 68832 24332
rect 68888 24276 68936 24332
rect 68992 24276 69040 24332
rect 69096 24276 69124 24332
rect 59144 23492 59172 23548
rect 59228 23492 59276 23548
rect 59332 23492 59380 23548
rect 59436 23492 59464 23548
rect 59144 21980 59464 23492
rect 60060 23604 60116 23614
rect 60060 23156 60116 23548
rect 60060 23090 60116 23100
rect 68804 22764 69124 24276
rect 68804 22708 68832 22764
rect 68888 22708 68936 22764
rect 68992 22708 69040 22764
rect 69096 22708 69124 22764
rect 59144 21924 59172 21980
rect 59228 21924 59276 21980
rect 59332 21924 59380 21980
rect 59436 21924 59464 21980
rect 51884 21812 51940 21822
rect 51884 21588 51940 21756
rect 51884 21522 51940 21532
rect 49484 21140 49512 21196
rect 49568 21140 49616 21196
rect 49672 21140 49720 21196
rect 49776 21140 49804 21196
rect 49484 19628 49804 21140
rect 49484 19572 49512 19628
rect 49568 19572 49616 19628
rect 49672 19572 49720 19628
rect 49776 19572 49804 19628
rect 49484 18060 49804 19572
rect 49484 18004 49512 18060
rect 49568 18004 49616 18060
rect 49672 18004 49720 18060
rect 49776 18004 49804 18060
rect 49484 16492 49804 18004
rect 49484 16436 49512 16492
rect 49568 16436 49616 16492
rect 49672 16436 49720 16492
rect 49776 16436 49804 16492
rect 49484 14924 49804 16436
rect 59144 20412 59464 21924
rect 65660 22036 65716 22046
rect 65660 21588 65716 21980
rect 65660 21522 65716 21532
rect 59144 20356 59172 20412
rect 59228 20356 59276 20412
rect 59332 20356 59380 20412
rect 59436 20356 59464 20412
rect 59144 18844 59464 20356
rect 59144 18788 59172 18844
rect 59228 18788 59276 18844
rect 59332 18788 59380 18844
rect 59436 18788 59464 18844
rect 59144 17276 59464 18788
rect 59144 17220 59172 17276
rect 59228 17220 59276 17276
rect 59332 17220 59380 17276
rect 59436 17220 59464 17276
rect 59144 15708 59464 17220
rect 59144 15652 59172 15708
rect 59228 15652 59276 15708
rect 59332 15652 59380 15708
rect 59436 15652 59464 15708
rect 49484 14868 49512 14924
rect 49568 14868 49616 14924
rect 49672 14868 49720 14924
rect 49776 14868 49804 14924
rect 49484 13356 49804 14868
rect 49484 13300 49512 13356
rect 49568 13300 49616 13356
rect 49672 13300 49720 13356
rect 49776 13300 49804 13356
rect 55356 15204 55412 15214
rect 55356 13412 55412 15148
rect 55356 13346 55412 13356
rect 59144 14140 59464 15652
rect 59144 14084 59172 14140
rect 59228 14084 59276 14140
rect 59332 14084 59380 14140
rect 59436 14084 59464 14140
rect 43596 12180 43652 12190
rect 43596 11732 43652 12124
rect 43596 11666 43652 11676
rect 49484 11788 49804 13300
rect 49484 11732 49512 11788
rect 49568 11732 49616 11788
rect 49672 11732 49720 11788
rect 49776 11732 49804 11788
rect 39824 10948 39852 11004
rect 39908 10948 39956 11004
rect 40012 10948 40060 11004
rect 40116 10948 40144 11004
rect 39824 9436 40144 10948
rect 39824 9380 39852 9436
rect 39908 9380 39956 9436
rect 40012 9380 40060 9436
rect 40116 9380 40144 9436
rect 39824 7868 40144 9380
rect 39824 7812 39852 7868
rect 39908 7812 39956 7868
rect 40012 7812 40060 7868
rect 40116 7812 40144 7868
rect 39824 6300 40144 7812
rect 39824 6244 39852 6300
rect 39908 6244 39956 6300
rect 40012 6244 40060 6300
rect 40116 6244 40144 6300
rect 31612 4788 31668 4798
rect 31612 4452 31668 4732
rect 31612 4386 31668 4396
rect 39676 4788 39732 4798
rect 30164 3892 30192 3948
rect 30248 3892 30296 3948
rect 30352 3892 30400 3948
rect 30456 3892 30484 3948
rect 30164 3076 30484 3892
rect 39676 3780 39732 4732
rect 39676 3714 39732 3724
rect 39824 4732 40144 6244
rect 39824 4676 39852 4732
rect 39908 4676 39956 4732
rect 40012 4676 40060 4732
rect 40116 4676 40144 4732
rect 39824 3164 40144 4676
rect 39824 3108 39852 3164
rect 39908 3108 39956 3164
rect 40012 3108 40060 3164
rect 40116 3108 40144 3164
rect 39824 3076 40144 3108
rect 49484 10220 49804 11732
rect 49484 10164 49512 10220
rect 49568 10164 49616 10220
rect 49672 10164 49720 10220
rect 49776 10164 49804 10220
rect 49484 8652 49804 10164
rect 49484 8596 49512 8652
rect 49568 8596 49616 8652
rect 49672 8596 49720 8652
rect 49776 8596 49804 8652
rect 49484 7084 49804 8596
rect 49484 7028 49512 7084
rect 49568 7028 49616 7084
rect 49672 7028 49720 7084
rect 49776 7028 49804 7084
rect 49484 5516 49804 7028
rect 59144 12572 59464 14084
rect 59144 12516 59172 12572
rect 59228 12516 59276 12572
rect 59332 12516 59380 12572
rect 59436 12516 59464 12572
rect 59144 11004 59464 12516
rect 59144 10948 59172 11004
rect 59228 10948 59276 11004
rect 59332 10948 59380 11004
rect 59436 10948 59464 11004
rect 59144 9436 59464 10948
rect 68804 21196 69124 22708
rect 68804 21140 68832 21196
rect 68888 21140 68936 21196
rect 68992 21140 69040 21196
rect 69096 21140 69124 21196
rect 68804 19628 69124 21140
rect 68804 19572 68832 19628
rect 68888 19572 68936 19628
rect 68992 19572 69040 19628
rect 69096 19572 69124 19628
rect 68804 18060 69124 19572
rect 68804 18004 68832 18060
rect 68888 18004 68936 18060
rect 68992 18004 69040 18060
rect 69096 18004 69124 18060
rect 68804 16492 69124 18004
rect 68804 16436 68832 16492
rect 68888 16436 68936 16492
rect 68992 16436 69040 16492
rect 69096 16436 69124 16492
rect 68804 14924 69124 16436
rect 68804 14868 68832 14924
rect 68888 14868 68936 14924
rect 68992 14868 69040 14924
rect 69096 14868 69124 14924
rect 68804 13356 69124 14868
rect 68804 13300 68832 13356
rect 68888 13300 68936 13356
rect 68992 13300 69040 13356
rect 69096 13300 69124 13356
rect 68804 11788 69124 13300
rect 68804 11732 68832 11788
rect 68888 11732 68936 11788
rect 68992 11732 69040 11788
rect 69096 11732 69124 11788
rect 68804 10220 69124 11732
rect 68804 10164 68832 10220
rect 68888 10164 68936 10220
rect 68992 10164 69040 10220
rect 69096 10164 69124 10220
rect 59144 9380 59172 9436
rect 59228 9380 59276 9436
rect 59332 9380 59380 9436
rect 59436 9380 59464 9436
rect 59144 7868 59464 9380
rect 61516 9940 61572 9950
rect 61516 9156 61572 9884
rect 61516 9090 61572 9100
rect 59144 7812 59172 7868
rect 59228 7812 59276 7868
rect 59332 7812 59380 7868
rect 59436 7812 59464 7868
rect 49484 5460 49512 5516
rect 49568 5460 49616 5516
rect 49672 5460 49720 5516
rect 49776 5460 49804 5516
rect 49484 3948 49804 5460
rect 55804 6692 55860 6702
rect 55804 5124 55860 6636
rect 59144 6300 59464 7812
rect 68804 8652 69124 10164
rect 68804 8596 68832 8652
rect 68888 8596 68936 8652
rect 68992 8596 69040 8652
rect 69096 8596 69124 8652
rect 68804 7084 69124 8596
rect 68804 7028 68832 7084
rect 68888 7028 68936 7084
rect 68992 7028 69040 7084
rect 69096 7028 69124 7084
rect 59144 6244 59172 6300
rect 59228 6244 59276 6300
rect 59332 6244 59380 6300
rect 59436 6244 59464 6300
rect 55916 6132 55972 6142
rect 55972 6076 56308 6132
rect 55916 6066 55972 6076
rect 56252 6020 56308 6076
rect 56252 5954 56308 5964
rect 55804 5058 55860 5068
rect 55412 5012 55468 5022
rect 55468 4956 55524 5012
rect 55412 4946 55524 4956
rect 55468 4676 55524 4946
rect 55468 4610 55524 4620
rect 59144 4732 59464 6244
rect 59144 4676 59172 4732
rect 59228 4676 59276 4732
rect 59332 4676 59380 4732
rect 59436 4676 59464 4732
rect 55916 4564 55972 4574
rect 55412 4340 55468 4350
rect 55804 4340 55860 4350
rect 55468 4284 55804 4340
rect 55412 4274 55468 4284
rect 55804 4274 55860 4284
rect 55916 4116 55972 4508
rect 55916 4050 55972 4060
rect 49484 3892 49512 3948
rect 49568 3892 49616 3948
rect 49672 3892 49720 3948
rect 49776 3892 49804 3948
rect 49484 3076 49804 3892
rect 59144 3164 59464 4676
rect 63868 6916 63924 6926
rect 63868 4676 63924 6860
rect 67228 6580 67284 6590
rect 67228 6244 67284 6524
rect 67228 6178 67284 6188
rect 67340 6356 67396 6366
rect 67340 6132 67396 6300
rect 67452 6132 67508 6142
rect 67340 6076 67452 6132
rect 67452 6066 67508 6076
rect 63868 4610 63924 4620
rect 68804 5516 69124 7028
rect 68804 5460 68832 5516
rect 68888 5460 68936 5516
rect 68992 5460 69040 5516
rect 69096 5460 69124 5516
rect 59144 3108 59172 3164
rect 59228 3108 59276 3164
rect 59332 3108 59380 3164
rect 59436 3108 59464 3164
rect 59144 3076 59464 3108
rect 68804 3948 69124 5460
rect 68804 3892 68832 3948
rect 68888 3892 68936 3948
rect 68992 3892 69040 3948
rect 69096 3892 69124 3948
rect 68804 3076 69124 3892
rect 78464 28196 78492 28252
rect 78548 28196 78596 28252
rect 78652 28196 78700 28252
rect 78756 28196 78784 28252
rect 78464 26684 78784 28196
rect 78464 26628 78492 26684
rect 78548 26628 78596 26684
rect 78652 26628 78700 26684
rect 78756 26628 78784 26684
rect 78464 25116 78784 26628
rect 78464 25060 78492 25116
rect 78548 25060 78596 25116
rect 78652 25060 78700 25116
rect 78756 25060 78784 25116
rect 78464 23548 78784 25060
rect 78464 23492 78492 23548
rect 78548 23492 78596 23548
rect 78652 23492 78700 23548
rect 78756 23492 78784 23548
rect 78464 21980 78784 23492
rect 78464 21924 78492 21980
rect 78548 21924 78596 21980
rect 78652 21924 78700 21980
rect 78756 21924 78784 21980
rect 78464 20412 78784 21924
rect 78464 20356 78492 20412
rect 78548 20356 78596 20412
rect 78652 20356 78700 20412
rect 78756 20356 78784 20412
rect 78464 18844 78784 20356
rect 78464 18788 78492 18844
rect 78548 18788 78596 18844
rect 78652 18788 78700 18844
rect 78756 18788 78784 18844
rect 78464 17276 78784 18788
rect 78464 17220 78492 17276
rect 78548 17220 78596 17276
rect 78652 17220 78700 17276
rect 78756 17220 78784 17276
rect 78464 15708 78784 17220
rect 78464 15652 78492 15708
rect 78548 15652 78596 15708
rect 78652 15652 78700 15708
rect 78756 15652 78784 15708
rect 78464 14140 78784 15652
rect 78464 14084 78492 14140
rect 78548 14084 78596 14140
rect 78652 14084 78700 14140
rect 78756 14084 78784 14140
rect 78464 12572 78784 14084
rect 78464 12516 78492 12572
rect 78548 12516 78596 12572
rect 78652 12516 78700 12572
rect 78756 12516 78784 12572
rect 78464 11004 78784 12516
rect 78464 10948 78492 11004
rect 78548 10948 78596 11004
rect 78652 10948 78700 11004
rect 78756 10948 78784 11004
rect 78464 9436 78784 10948
rect 78464 9380 78492 9436
rect 78548 9380 78596 9436
rect 78652 9380 78700 9436
rect 78756 9380 78784 9436
rect 78464 7868 78784 9380
rect 78464 7812 78492 7868
rect 78548 7812 78596 7868
rect 78652 7812 78700 7868
rect 78756 7812 78784 7868
rect 78464 6300 78784 7812
rect 78464 6244 78492 6300
rect 78548 6244 78596 6300
rect 78652 6244 78700 6300
rect 78756 6244 78784 6300
rect 78464 4732 78784 6244
rect 78464 4676 78492 4732
rect 78548 4676 78596 4732
rect 78652 4676 78700 4732
rect 78756 4676 78784 4732
rect 78464 3164 78784 4676
rect 78464 3108 78492 3164
rect 78548 3108 78596 3164
rect 78652 3108 78700 3164
rect 78756 3108 78784 3164
rect 78464 3076 78784 3108
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1387__I Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 1904 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1388__I
timestamp 1669390400
transform 1 0 36176 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1389__I
timestamp 1669390400
transform -1 0 21728 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1390__I
timestamp 1669390400
transform 1 0 22624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1391__I
timestamp 1669390400
transform 1 0 22624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1392__A1
timestamp 1669390400
transform -1 0 19824 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1392__A2
timestamp 1669390400
transform 1 0 20048 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1394__I
timestamp 1669390400
transform 1 0 20160 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1395__I
timestamp 1669390400
transform 1 0 20272 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1396__I
timestamp 1669390400
transform -1 0 21952 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1397__I
timestamp 1669390400
transform 1 0 22960 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1398__I
timestamp 1669390400
transform 1 0 24752 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1399__A1
timestamp 1669390400
transform 1 0 17024 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1399__A2
timestamp 1669390400
transform 1 0 17472 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1400__I
timestamp 1669390400
transform -1 0 44464 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1401__I
timestamp 1669390400
transform 1 0 16128 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1402__I
timestamp 1669390400
transform 1 0 15680 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1403__I
timestamp 1669390400
transform 1 0 25536 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1404__A1
timestamp 1669390400
transform -1 0 17024 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1404__A2
timestamp 1669390400
transform 1 0 16464 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1406__A1
timestamp 1669390400
transform 1 0 21952 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1406__A2
timestamp 1669390400
transform 1 0 24528 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1408__A1
timestamp 1669390400
transform 1 0 21392 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1408__A2
timestamp 1669390400
transform -1 0 22512 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1408__A3
timestamp 1669390400
transform 1 0 21840 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1412__I
timestamp 1669390400
transform 1 0 16240 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1413__I
timestamp 1669390400
transform 1 0 14784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1414__A1
timestamp 1669390400
transform 1 0 15904 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1414__A2
timestamp 1669390400
transform -1 0 15456 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1418__A1
timestamp 1669390400
transform -1 0 17136 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1418__A2
timestamp 1669390400
transform -1 0 16800 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1419__A1
timestamp 1669390400
transform 1 0 16128 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1419__A2
timestamp 1669390400
transform 1 0 17360 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1420__I
timestamp 1669390400
transform -1 0 8288 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1421__I
timestamp 1669390400
transform 1 0 23520 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1422__A1
timestamp 1669390400
transform 1 0 20720 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1422__A2
timestamp 1669390400
transform 1 0 20832 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1429__A1
timestamp 1669390400
transform 1 0 12656 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1429__A2
timestamp 1669390400
transform -1 0 13888 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1430__I
timestamp 1669390400
transform -1 0 47152 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1431__I
timestamp 1669390400
transform 1 0 49392 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1432__A1
timestamp 1669390400
transform 1 0 15568 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1432__A2
timestamp 1669390400
transform -1 0 16240 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1434__A1
timestamp 1669390400
transform -1 0 15680 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1434__A2
timestamp 1669390400
transform -1 0 13776 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1437__A1
timestamp 1669390400
transform 1 0 20496 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1437__A2
timestamp 1669390400
transform -1 0 21168 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1438__A1
timestamp 1669390400
transform 1 0 21952 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1438__A2
timestamp 1669390400
transform 1 0 21504 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1438__B1
timestamp 1669390400
transform 1 0 22400 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1438__B2
timestamp 1669390400
transform 1 0 21504 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1440__A1
timestamp 1669390400
transform 1 0 17696 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1440__A2
timestamp 1669390400
transform 1 0 17248 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1441__I
timestamp 1669390400
transform 1 0 14672 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1442__I
timestamp 1669390400
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1443__A1
timestamp 1669390400
transform -1 0 22400 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1443__A2
timestamp 1669390400
transform 1 0 19936 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1445__A1
timestamp 1669390400
transform 1 0 17136 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1445__A2
timestamp 1669390400
transform 1 0 17584 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1452__A1
timestamp 1669390400
transform -1 0 16128 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1452__A2
timestamp 1669390400
transform 1 0 16128 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1453__A1
timestamp 1669390400
transform 1 0 16352 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1453__A2
timestamp 1669390400
transform 1 0 16576 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1455__I
timestamp 1669390400
transform -1 0 58464 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1456__I
timestamp 1669390400
transform -1 0 11872 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1457__A1
timestamp 1669390400
transform 1 0 9632 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1457__A2
timestamp 1669390400
transform 1 0 9184 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1458__A1
timestamp 1669390400
transform -1 0 12096 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1458__A2
timestamp 1669390400
transform 1 0 12880 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1461__A1
timestamp 1669390400
transform 1 0 20048 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1461__A2
timestamp 1669390400
transform 1 0 19488 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1462__A1
timestamp 1669390400
transform 1 0 22848 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1462__A2
timestamp 1669390400
transform 1 0 24080 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1462__B1
timestamp 1669390400
transform 1 0 22288 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1462__B2
timestamp 1669390400
transform 1 0 21952 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1464__A1
timestamp 1669390400
transform 1 0 18480 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1464__A2
timestamp 1669390400
transform 1 0 18032 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1465__I
timestamp 1669390400
transform 1 0 5376 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1466__I
timestamp 1669390400
transform 1 0 48608 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1467__A1
timestamp 1669390400
transform 1 0 21280 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1467__A2
timestamp 1669390400
transform 1 0 19600 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1469__A1
timestamp 1669390400
transform 1 0 12544 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1469__A2
timestamp 1669390400
transform 1 0 12096 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1475__A1
timestamp 1669390400
transform -1 0 11088 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1475__A2
timestamp 1669390400
transform -1 0 11536 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1478__A1
timestamp 1669390400
transform 1 0 17248 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1479__A1
timestamp 1669390400
transform -1 0 11872 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1479__A2
timestamp 1669390400
transform 1 0 11984 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1482__I
timestamp 1669390400
transform 1 0 7056 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1483__A1
timestamp 1669390400
transform 1 0 7952 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1483__A2
timestamp 1669390400
transform -1 0 7168 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1485__A1
timestamp 1669390400
transform 1 0 13328 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1485__A2
timestamp 1669390400
transform 1 0 12880 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1487__A1
timestamp 1669390400
transform 1 0 19152 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1487__A2
timestamp 1669390400
transform 1 0 19600 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1488__A1
timestamp 1669390400
transform 1 0 20832 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1488__A2
timestamp 1669390400
transform 1 0 24528 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1488__B1
timestamp 1669390400
transform -1 0 23744 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1488__B2
timestamp 1669390400
transform 1 0 23072 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1490__A1
timestamp 1669390400
transform 1 0 17136 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1490__A2
timestamp 1669390400
transform 1 0 16128 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1491__I
timestamp 1669390400
transform 1 0 9632 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1492__A1
timestamp 1669390400
transform -1 0 16352 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1492__A2
timestamp 1669390400
transform 1 0 15232 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1495__A1
timestamp 1669390400
transform -1 0 9856 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1495__A2
timestamp 1669390400
transform 1 0 12096 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1497__A1
timestamp 1669390400
transform 1 0 14448 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1497__A2
timestamp 1669390400
transform 1 0 12880 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1500__A3
timestamp 1669390400
transform 1 0 11872 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1505__A1
timestamp 1669390400
transform 1 0 15568 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1508__A1
timestamp 1669390400
transform 1 0 12432 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1508__A2
timestamp 1669390400
transform 1 0 12544 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1511__I
timestamp 1669390400
transform 1 0 2464 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1512__A1
timestamp 1669390400
transform -1 0 15232 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1512__A2
timestamp 1669390400
transform 1 0 12880 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1512__B1
timestamp 1669390400
transform 1 0 12432 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1512__B2
timestamp 1669390400
transform -1 0 14784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1513__A1
timestamp 1669390400
transform 1 0 4816 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1513__A2
timestamp 1669390400
transform 1 0 4368 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1516__A1
timestamp 1669390400
transform -1 0 4928 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1517__A1
timestamp 1669390400
transform 1 0 5040 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1520__A1
timestamp 1669390400
transform -1 0 15904 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1520__A2
timestamp 1669390400
transform -1 0 18816 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1521__A1
timestamp 1669390400
transform 1 0 19376 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1521__A2
timestamp 1669390400
transform 1 0 19712 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1521__B1
timestamp 1669390400
transform -1 0 17136 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1521__B2
timestamp 1669390400
transform 1 0 19152 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1523__A1
timestamp 1669390400
transform -1 0 16240 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1523__A2
timestamp 1669390400
transform 1 0 15232 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1524__I
timestamp 1669390400
transform 1 0 8400 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1525__I
timestamp 1669390400
transform 1 0 67424 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1526__A1
timestamp 1669390400
transform 1 0 19600 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1526__A2
timestamp 1669390400
transform 1 0 19936 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1528__A1
timestamp 1669390400
transform -1 0 8288 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1528__A2
timestamp 1669390400
transform -1 0 7840 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1529__A1
timestamp 1669390400
transform -1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1529__A2
timestamp 1669390400
transform 1 0 9184 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1530__A1
timestamp 1669390400
transform 1 0 9632 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1530__A2
timestamp 1669390400
transform 1 0 11760 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1530__A3
timestamp 1669390400
transform 1 0 12208 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1530__A4
timestamp 1669390400
transform 1 0 11312 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1531__A1
timestamp 1669390400
transform 1 0 21840 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1531__A2
timestamp 1669390400
transform 1 0 23968 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1531__B1
timestamp 1669390400
transform 1 0 24416 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1531__B2
timestamp 1669390400
transform 1 0 23968 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1532__A2
timestamp 1669390400
transform -1 0 8736 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1535__A1
timestamp 1669390400
transform 1 0 7952 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1536__A1
timestamp 1669390400
transform 1 0 7728 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1538__A3
timestamp 1669390400
transform -1 0 8512 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1541__I
timestamp 1669390400
transform 1 0 9632 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1542__A1
timestamp 1669390400
transform -1 0 2240 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1542__A2
timestamp 1669390400
transform -1 0 2240 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1543__A1
timestamp 1669390400
transform 1 0 6048 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1543__A2
timestamp 1669390400
transform -1 0 6720 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1544__A2
timestamp 1669390400
transform 1 0 5040 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1548__A1
timestamp 1669390400
transform -1 0 6272 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1548__A2
timestamp 1669390400
transform 1 0 7728 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1550__A1
timestamp 1669390400
transform -1 0 8400 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1550__A2
timestamp 1669390400
transform -1 0 7952 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1551__A1
timestamp 1669390400
transform 1 0 8624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1551__A2
timestamp 1669390400
transform 1 0 9856 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1552__A1
timestamp 1669390400
transform 1 0 12768 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1552__A2
timestamp 1669390400
transform 1 0 11760 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1554__A1
timestamp 1669390400
transform 1 0 19152 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1554__A2
timestamp 1669390400
transform 1 0 16128 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1555__I
timestamp 1669390400
transform 1 0 46816 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1556__A1
timestamp 1669390400
transform 1 0 21504 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1556__A2
timestamp 1669390400
transform 1 0 20608 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1556__B1
timestamp 1669390400
transform 1 0 20384 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1556__B2
timestamp 1669390400
transform 1 0 20832 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1558__A1
timestamp 1669390400
transform 1 0 16128 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1558__A2
timestamp 1669390400
transform 1 0 15680 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1559__I
timestamp 1669390400
transform 1 0 28448 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1560__I
timestamp 1669390400
transform 1 0 15568 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1561__A1
timestamp 1669390400
transform -1 0 22624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1561__A2
timestamp 1669390400
transform 1 0 17808 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1565__A3
timestamp 1669390400
transform 1 0 4928 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1567__A1
timestamp 1669390400
transform 1 0 9520 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1567__A2
timestamp 1669390400
transform -1 0 8288 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1568__A2
timestamp 1669390400
transform -1 0 8288 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1569__A2
timestamp 1669390400
transform 1 0 9856 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1574__A1
timestamp 1669390400
transform 1 0 8960 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1576__A1
timestamp 1669390400
transform 1 0 10304 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1578__A1
timestamp 1669390400
transform 1 0 20384 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1578__A2
timestamp 1669390400
transform -1 0 18256 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1578__A3
timestamp 1669390400
transform 1 0 16912 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1579__A1
timestamp 1669390400
transform 1 0 15120 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1581__A1
timestamp 1669390400
transform 1 0 16464 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1582__A1
timestamp 1669390400
transform 1 0 9632 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1583__A1
timestamp 1669390400
transform 1 0 14336 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1585__A2
timestamp 1669390400
transform 1 0 20496 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1590__I
timestamp 1669390400
transform -1 0 28224 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1591__I
timestamp 1669390400
transform -1 0 24864 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1592__A1
timestamp 1669390400
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1593__A1
timestamp 1669390400
transform -1 0 24640 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1594__A2
timestamp 1669390400
transform 1 0 5600 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1595__A2
timestamp 1669390400
transform 1 0 7056 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1597__A2
timestamp 1669390400
transform -1 0 3136 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1600__A1
timestamp 1669390400
transform 1 0 11088 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1600__A2
timestamp 1669390400
transform 1 0 11536 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1601__A1
timestamp 1669390400
transform 1 0 8960 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1601__A2
timestamp 1669390400
transform 1 0 7952 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1604__A1
timestamp 1669390400
transform 1 0 2464 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1604__A2
timestamp 1669390400
transform 1 0 5600 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1605__A1
timestamp 1669390400
transform 1 0 5600 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1605__A2
timestamp 1669390400
transform 1 0 6048 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1606__A1
timestamp 1669390400
transform 1 0 8176 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1606__A2
timestamp 1669390400
transform -1 0 6720 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1612__A1
timestamp 1669390400
transform 1 0 10528 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1612__A2
timestamp 1669390400
transform 1 0 10416 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1613__A1
timestamp 1669390400
transform 1 0 14112 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1613__A2
timestamp 1669390400
transform 1 0 14336 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1615__A1
timestamp 1669390400
transform -1 0 17360 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1615__A2
timestamp 1669390400
transform 1 0 16688 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1616__A1
timestamp 1669390400
transform 1 0 16688 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1616__A2
timestamp 1669390400
transform -1 0 16016 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1616__B1
timestamp 1669390400
transform 1 0 16240 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1616__B2
timestamp 1669390400
transform 1 0 17136 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1618__A1
timestamp 1669390400
transform 1 0 16128 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1618__A2
timestamp 1669390400
transform 1 0 15680 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1619__I
timestamp 1669390400
transform 1 0 30912 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1620__A1
timestamp 1669390400
transform 1 0 17808 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1620__A2
timestamp 1669390400
transform -1 0 22176 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1623__A1
timestamp 1669390400
transform -1 0 21056 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1624__A3
timestamp 1669390400
transform 1 0 15456 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1625__A1
timestamp 1669390400
transform 1 0 13888 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1626__A2
timestamp 1669390400
transform -1 0 22960 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1630__A2
timestamp 1669390400
transform -1 0 23520 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1631__A1
timestamp 1669390400
transform 1 0 24304 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1631__A2
timestamp 1669390400
transform -1 0 22064 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1632__A1
timestamp 1669390400
transform 1 0 22736 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1632__A2
timestamp 1669390400
transform -1 0 22512 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1633__A2
timestamp 1669390400
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1640__A2
timestamp 1669390400
transform -1 0 25088 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1643__A1
timestamp 1669390400
transform -1 0 25984 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1643__A3
timestamp 1669390400
transform -1 0 26432 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1644__A1
timestamp 1669390400
transform 1 0 12880 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1645__A2
timestamp 1669390400
transform 1 0 22960 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1649__A1
timestamp 1669390400
transform 1 0 25984 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1650__I
timestamp 1669390400
transform 1 0 58464 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1651__I
timestamp 1669390400
transform 1 0 58464 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1652__A1
timestamp 1669390400
transform -1 0 27440 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1652__A2
timestamp 1669390400
transform -1 0 28224 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1653__A1
timestamp 1669390400
transform 1 0 25984 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1653__A2
timestamp 1669390400
transform 1 0 25536 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1653__A4
timestamp 1669390400
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1656__A1
timestamp 1669390400
transform -1 0 26992 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1657__A2
timestamp 1669390400
transform -1 0 12208 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1658__A2
timestamp 1669390400
transform 1 0 15232 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1660__A1
timestamp 1669390400
transform 1 0 6384 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1660__A2
timestamp 1669390400
transform 1 0 6160 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1662__A1
timestamp 1669390400
transform 1 0 5040 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1662__A2
timestamp 1669390400
transform 1 0 4592 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1663__A1
timestamp 1669390400
transform 1 0 10416 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1663__A2
timestamp 1669390400
transform 1 0 9184 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1666__A1
timestamp 1669390400
transform 1 0 5264 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1666__A2
timestamp 1669390400
transform 1 0 5712 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1667__A1
timestamp 1669390400
transform 1 0 4928 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1668__A1
timestamp 1669390400
transform -1 0 2464 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1668__A2
timestamp 1669390400
transform 1 0 4928 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1673__A1
timestamp 1669390400
transform -1 0 22848 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1674__A1
timestamp 1669390400
transform 1 0 14560 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1674__A2
timestamp 1669390400
transform 1 0 12320 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1675__A1
timestamp 1669390400
transform 1 0 15232 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1675__A2
timestamp 1669390400
transform 1 0 14336 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1677__A1
timestamp 1669390400
transform 1 0 19824 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1677__A2
timestamp 1669390400
transform -1 0 21728 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1678__I
timestamp 1669390400
transform 1 0 15904 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1679__A1
timestamp 1669390400
transform -1 0 17136 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1679__A2
timestamp 1669390400
transform 1 0 15680 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1679__B1
timestamp 1669390400
transform 1 0 16464 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1679__B2
timestamp 1669390400
transform -1 0 16352 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1681__A1
timestamp 1669390400
transform -1 0 17136 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1681__A2
timestamp 1669390400
transform 1 0 17584 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1682__I
timestamp 1669390400
transform 1 0 40768 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1683__I
timestamp 1669390400
transform 1 0 64624 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1684__A1
timestamp 1669390400
transform 1 0 22848 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1684__A2
timestamp 1669390400
transform 1 0 23296 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1687__A1
timestamp 1669390400
transform 1 0 23296 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1688__A1
timestamp 1669390400
transform 1 0 22176 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1689__A1
timestamp 1669390400
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1689__A2
timestamp 1669390400
transform -1 0 25424 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1693__A2
timestamp 1669390400
transform 1 0 23968 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1695__A1
timestamp 1669390400
transform 1 0 29568 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1699__A1
timestamp 1669390400
transform 1 0 29792 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1700__A1
timestamp 1669390400
transform 1 0 25200 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1700__A2
timestamp 1669390400
transform -1 0 24976 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1707__I
timestamp 1669390400
transform 1 0 64624 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1708__A1
timestamp 1669390400
transform 1 0 25648 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1708__A2
timestamp 1669390400
transform -1 0 26320 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1709__A1
timestamp 1669390400
transform 1 0 28224 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1709__A2
timestamp 1669390400
transform -1 0 29680 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1711__A1
timestamp 1669390400
transform 1 0 25536 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1711__B1
timestamp 1669390400
transform 1 0 28224 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1711__B2
timestamp 1669390400
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1715__A1
timestamp 1669390400
transform 1 0 29568 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1718__A1
timestamp 1669390400
transform 1 0 23520 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1719__A1
timestamp 1669390400
transform 1 0 3696 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1719__A2
timestamp 1669390400
transform -1 0 1904 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1720__A2
timestamp 1669390400
transform 1 0 5264 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1723__A1
timestamp 1669390400
transform 1 0 11872 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1723__A2
timestamp 1669390400
transform 1 0 15232 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1726__A1
timestamp 1669390400
transform 1 0 2800 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1726__A2
timestamp 1669390400
transform -1 0 1904 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1727__A1
timestamp 1669390400
transform -1 0 2576 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1727__A2
timestamp 1669390400
transform -1 0 2128 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1728__A1
timestamp 1669390400
transform -1 0 2128 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1733__A1
timestamp 1669390400
transform 1 0 23744 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1734__A1
timestamp 1669390400
transform 1 0 14784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1734__A2
timestamp 1669390400
transform 1 0 14336 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1735__A1
timestamp 1669390400
transform 1 0 14784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1735__A2
timestamp 1669390400
transform 1 0 15232 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1737__A1
timestamp 1669390400
transform 1 0 21504 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1737__A2
timestamp 1669390400
transform 1 0 21056 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1738__A1
timestamp 1669390400
transform -1 0 21728 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1738__A2
timestamp 1669390400
transform 1 0 19824 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1738__B1
timestamp 1669390400
transform 1 0 22848 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1738__B2
timestamp 1669390400
transform -1 0 20720 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1740__A1
timestamp 1669390400
transform -1 0 16240 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1740__A2
timestamp 1669390400
transform 1 0 16464 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1741__I
timestamp 1669390400
transform 1 0 69328 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1742__I
timestamp 1669390400
transform 1 0 66080 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1743__A1
timestamp 1669390400
transform 1 0 20048 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1743__A2
timestamp 1669390400
transform 1 0 20496 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1746__A1
timestamp 1669390400
transform -1 0 24752 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1747__A1
timestamp 1669390400
transform -1 0 25536 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1748__A1
timestamp 1669390400
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1748__A2
timestamp 1669390400
transform 1 0 29344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1750__A1
timestamp 1669390400
transform 1 0 32032 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1754__A1
timestamp 1669390400
transform 1 0 30688 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1763__A1
timestamp 1669390400
transform 1 0 46144 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1763__A2
timestamp 1669390400
transform 1 0 46592 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1767__A1
timestamp 1669390400
transform 1 0 32816 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1768__A1
timestamp 1669390400
transform 1 0 32144 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1769__A1
timestamp 1669390400
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1769__A2
timestamp 1669390400
transform -1 0 30688 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1774__I
timestamp 1669390400
transform 1 0 66528 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1775__I
timestamp 1669390400
transform 1 0 64512 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1776__A1
timestamp 1669390400
transform 1 0 30016 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1776__A2
timestamp 1669390400
transform -1 0 31248 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1779__A1
timestamp 1669390400
transform 1 0 25872 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1779__A2
timestamp 1669390400
transform -1 0 26992 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1780__A1
timestamp 1669390400
transform 1 0 24192 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1780__A2
timestamp 1669390400
transform 1 0 26768 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1784__A1
timestamp 1669390400
transform -1 0 31696 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1788__A1
timestamp 1669390400
transform -1 0 25872 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1789__A1
timestamp 1669390400
transform 1 0 5600 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1789__A2
timestamp 1669390400
transform 1 0 5824 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1791__A1
timestamp 1669390400
transform 1 0 15568 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1791__A2
timestamp 1669390400
transform 1 0 15120 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1794__A1
timestamp 1669390400
transform 1 0 3696 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1794__A2
timestamp 1669390400
transform 1 0 1904 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1795__A1
timestamp 1669390400
transform 1 0 8960 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1795__A2
timestamp 1669390400
transform 1 0 7728 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1800__A1
timestamp 1669390400
transform 1 0 26656 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1801__A1
timestamp 1669390400
transform 1 0 11760 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1801__A2
timestamp 1669390400
transform -1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1802__A1
timestamp 1669390400
transform 1 0 15680 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1802__A2
timestamp 1669390400
transform 1 0 16128 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1804__A1
timestamp 1669390400
transform 1 0 20608 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1804__A2
timestamp 1669390400
transform 1 0 21616 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1805__A1
timestamp 1669390400
transform -1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1805__A2
timestamp 1669390400
transform 1 0 21952 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1805__B1
timestamp 1669390400
transform 1 0 22848 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1805__B2
timestamp 1669390400
transform 1 0 22400 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1807__A1
timestamp 1669390400
transform 1 0 16688 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1807__A2
timestamp 1669390400
transform 1 0 16240 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1808__I
timestamp 1669390400
transform 1 0 30912 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1809__I
timestamp 1669390400
transform 1 0 20944 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1810__A1
timestamp 1669390400
transform -1 0 24528 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1810__A2
timestamp 1669390400
transform 1 0 22288 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1813__A1
timestamp 1669390400
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1814__A1
timestamp 1669390400
transform -1 0 27552 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1815__A2
timestamp 1669390400
transform -1 0 34496 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1815__A3
timestamp 1669390400
transform 1 0 33824 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1816__A1
timestamp 1669390400
transform -1 0 36960 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1824__A1
timestamp 1669390400
transform 1 0 34272 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1827__A1
timestamp 1669390400
transform 1 0 33824 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1827__A2
timestamp 1669390400
transform 1 0 33376 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1828__A1
timestamp 1669390400
transform 1 0 36064 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1828__A2
timestamp 1669390400
transform 1 0 37408 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1832__A1
timestamp 1669390400
transform 1 0 27440 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1834__A1
timestamp 1669390400
transform -1 0 2016 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1834__A2
timestamp 1669390400
transform -1 0 2240 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1837__A1
timestamp 1669390400
transform 1 0 11984 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1837__A2
timestamp 1669390400
transform 1 0 12432 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1838__A1
timestamp 1669390400
transform 1 0 12880 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1838__A2
timestamp 1669390400
transform -1 0 15232 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1838__B1
timestamp 1669390400
transform -1 0 14784 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1838__B2
timestamp 1669390400
transform 1 0 14336 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1840__A1
timestamp 1669390400
transform 1 0 8848 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1840__A2
timestamp 1669390400
transform -1 0 9520 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1841__A1
timestamp 1669390400
transform 1 0 9744 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1841__A2
timestamp 1669390400
transform -1 0 7280 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1846__A1
timestamp 1669390400
transform -1 0 26544 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1847__A1
timestamp 1669390400
transform 1 0 15456 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1847__A2
timestamp 1669390400
transform -1 0 12656 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1848__A1
timestamp 1669390400
transform 1 0 15344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1848__A2
timestamp 1669390400
transform 1 0 15792 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1850__A1
timestamp 1669390400
transform 1 0 17584 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1850__A2
timestamp 1669390400
transform 1 0 16576 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1851__A1
timestamp 1669390400
transform -1 0 20832 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1851__A2
timestamp 1669390400
transform -1 0 16688 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1851__B1
timestamp 1669390400
transform -1 0 17136 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1851__B2
timestamp 1669390400
transform 1 0 17584 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1853__A1
timestamp 1669390400
transform 1 0 19488 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1853__A2
timestamp 1669390400
transform 1 0 19040 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1854__I
timestamp 1669390400
transform -1 0 64176 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1855__I
timestamp 1669390400
transform 1 0 61824 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1856__A1
timestamp 1669390400
transform 1 0 25648 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1856__A2
timestamp 1669390400
transform 1 0 25536 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1857__A3
timestamp 1669390400
transform 1 0 19936 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1860__A1
timestamp 1669390400
transform 1 0 28112 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1860__A3
timestamp 1669390400
transform -1 0 28112 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1861__A1
timestamp 1669390400
transform 1 0 35504 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1861__A2
timestamp 1669390400
transform 1 0 35056 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1862__A1
timestamp 1669390400
transform 1 0 30912 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1862__A2
timestamp 1669390400
transform 1 0 32368 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1867__I
timestamp 1669390400
transform 1 0 66528 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1868__I
timestamp 1669390400
transform 1 0 65296 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1869__A1
timestamp 1669390400
transform 1 0 39088 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1869__A2
timestamp 1669390400
transform 1 0 41216 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1869__B1
timestamp 1669390400
transform 1 0 40768 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1869__B2
timestamp 1669390400
transform 1 0 38640 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1870__A1
timestamp 1669390400
transform 1 0 38528 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1870__A2
timestamp 1669390400
transform -1 0 39424 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1870__A3
timestamp 1669390400
transform 1 0 41664 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1870__A4
timestamp 1669390400
transform 1 0 42112 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1873__A1
timestamp 1669390400
transform 1 0 25872 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1874__A1
timestamp 1669390400
transform -1 0 25200 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1874__A2
timestamp 1669390400
transform -1 0 25648 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1875__A1
timestamp 1669390400
transform 1 0 24416 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1875__B1
timestamp 1669390400
transform 1 0 27888 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1875__B2
timestamp 1669390400
transform 1 0 24864 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1877__A1
timestamp 1669390400
transform 1 0 28560 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1877__A2
timestamp 1669390400
transform 1 0 28112 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1878__A1
timestamp 1669390400
transform 1 0 27104 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1878__A2
timestamp 1669390400
transform 1 0 26880 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1882__A1
timestamp 1669390400
transform 1 0 33824 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1885__A1
timestamp 1669390400
transform -1 0 39088 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1889__A1
timestamp 1669390400
transform 1 0 39200 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1896__A1
timestamp 1669390400
transform 1 0 41664 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1898__A1
timestamp 1669390400
transform -1 0 33824 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1900__A1
timestamp 1669390400
transform -1 0 36176 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1900__A2
timestamp 1669390400
transform -1 0 35728 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1907__I
timestamp 1669390400
transform 1 0 71568 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1908__A1
timestamp 1669390400
transform 1 0 39536 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1908__A2
timestamp 1669390400
transform 1 0 41552 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1909__A1
timestamp 1669390400
transform 1 0 39424 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1909__A2
timestamp 1669390400
transform 1 0 40656 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1910__A1
timestamp 1669390400
transform 1 0 38976 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1910__A2
timestamp 1669390400
transform -1 0 41664 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1913__A1
timestamp 1669390400
transform 1 0 26320 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1913__A2
timestamp 1669390400
transform 1 0 28560 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1914__A1
timestamp 1669390400
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1914__B1
timestamp 1669390400
transform 1 0 25872 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1914__B2
timestamp 1669390400
transform 1 0 24416 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1916__A1
timestamp 1669390400
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1916__A2
timestamp 1669390400
transform 1 0 29008 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1917__A1
timestamp 1669390400
transform -1 0 32256 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1917__A2
timestamp 1669390400
transform 1 0 29680 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1921__A1
timestamp 1669390400
transform -1 0 32704 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1923__A2
timestamp 1669390400
transform -1 0 27440 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1924__A2
timestamp 1669390400
transform 1 0 30240 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1925__A1
timestamp 1669390400
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1926__A1
timestamp 1669390400
transform -1 0 10752 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1926__A2
timestamp 1669390400
transform 1 0 10976 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1929__A1
timestamp 1669390400
transform 1 0 17584 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1929__A2
timestamp 1669390400
transform 1 0 16800 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1932__A1
timestamp 1669390400
transform 1 0 6608 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1932__A2
timestamp 1669390400
transform -1 0 5936 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1933__A1
timestamp 1669390400
transform 1 0 8848 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1933__A2
timestamp 1669390400
transform -1 0 11200 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1940__A1
timestamp 1669390400
transform 1 0 11984 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1940__A2
timestamp 1669390400
transform 1 0 12768 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1941__A1
timestamp 1669390400
transform 1 0 17024 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1941__A2
timestamp 1669390400
transform -1 0 15568 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1943__A1
timestamp 1669390400
transform -1 0 21728 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1943__A2
timestamp 1669390400
transform -1 0 23296 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1944__A1
timestamp 1669390400
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1944__A2
timestamp 1669390400
transform 1 0 24416 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1944__B1
timestamp 1669390400
transform 1 0 24752 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1944__B2
timestamp 1669390400
transform 1 0 25984 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1946__A1
timestamp 1669390400
transform 1 0 22848 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1946__A2
timestamp 1669390400
transform -1 0 25536 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1947__I
timestamp 1669390400
transform 1 0 63504 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1948__A1
timestamp 1669390400
transform 1 0 41888 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1948__A2
timestamp 1669390400
transform 1 0 42672 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1949__A3
timestamp 1669390400
transform 1 0 26432 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1953__A1
timestamp 1669390400
transform -1 0 25536 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1954__A1
timestamp 1669390400
transform 1 0 37184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1954__A2
timestamp 1669390400
transform 1 0 35952 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1955__A2
timestamp 1669390400
transform -1 0 38192 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1956__A3
timestamp 1669390400
transform -1 0 41440 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1963__A1
timestamp 1669390400
transform 1 0 50512 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1966__A1
timestamp 1669390400
transform 1 0 53088 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1970__A2
timestamp 1669390400
transform 1 0 38528 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1971__A2
timestamp 1669390400
transform 1 0 39984 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1973__I
timestamp 1669390400
transform 1 0 68320 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1974__A1
timestamp 1669390400
transform 1 0 43120 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1974__A2
timestamp 1669390400
transform 1 0 45472 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1975__A1
timestamp 1669390400
transform 1 0 35056 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1983__A1
timestamp 1669390400
transform 1 0 35504 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1983__A2
timestamp 1669390400
transform 1 0 35952 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1984__A2
timestamp 1669390400
transform 1 0 38080 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1984__B
timestamp 1669390400
transform -1 0 36960 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1991__A1
timestamp 1669390400
transform 1 0 38640 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1991__A2
timestamp 1669390400
transform 1 0 40992 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1992__A1
timestamp 1669390400
transform 1 0 40880 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1992__A2
timestamp 1669390400
transform -1 0 42784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1994__A1
timestamp 1669390400
transform -1 0 37856 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1994__A2
timestamp 1669390400
transform 1 0 38976 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1994__B1
timestamp 1669390400
transform 1 0 39088 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1994__B2
timestamp 1669390400
transform 1 0 38080 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1997__A1
timestamp 1669390400
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1997__A2
timestamp 1669390400
transform 1 0 30016 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2000__A1
timestamp 1669390400
transform 1 0 26656 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2000__A2
timestamp 1669390400
transform 1 0 28112 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2001__A1
timestamp 1669390400
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2001__A2
timestamp 1669390400
transform 1 0 29568 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2005__A1
timestamp 1669390400
transform 1 0 33712 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2008__A1
timestamp 1669390400
transform -1 0 25088 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2009__A1
timestamp 1669390400
transform 1 0 10416 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2009__A2
timestamp 1669390400
transform 1 0 10864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2010__A2
timestamp 1669390400
transform 1 0 5600 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2011__A1
timestamp 1669390400
transform 1 0 19152 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2011__A2
timestamp 1669390400
transform 1 0 18928 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2013__A2
timestamp 1669390400
transform -1 0 16912 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2014__A1
timestamp 1669390400
transform 1 0 7952 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2014__A2
timestamp 1669390400
transform -1 0 7728 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2015__A1
timestamp 1669390400
transform 1 0 11312 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2015__A2
timestamp 1669390400
transform 1 0 10864 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2016__A1
timestamp 1669390400
transform 1 0 7392 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2017__A1
timestamp 1669390400
transform -1 0 4592 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2021__A1
timestamp 1669390400
transform -1 0 34160 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2021__A2
timestamp 1669390400
transform 1 0 33824 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2022__A1
timestamp 1669390400
transform 1 0 17472 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2022__A2
timestamp 1669390400
transform -1 0 17136 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2023__A1
timestamp 1669390400
transform -1 0 13888 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2023__A2
timestamp 1669390400
transform -1 0 17584 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2024__A2
timestamp 1669390400
transform -1 0 42224 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2025__I
timestamp 1669390400
transform -1 0 54880 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2026__A1
timestamp 1669390400
transform -1 0 27776 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2026__A2
timestamp 1669390400
transform 1 0 26992 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2026__B1
timestamp 1669390400
transform -1 0 27328 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2026__B2
timestamp 1669390400
transform -1 0 28224 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2027__A1
timestamp 1669390400
transform -1 0 23520 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2027__A2
timestamp 1669390400
transform -1 0 26320 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2028__A1
timestamp 1669390400
transform -1 0 38304 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2028__A2
timestamp 1669390400
transform -1 0 36512 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2029__I
timestamp 1669390400
transform -1 0 54432 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2030__A1
timestamp 1669390400
transform 1 0 31248 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2030__A2
timestamp 1669390400
transform -1 0 29008 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2031__A1
timestamp 1669390400
transform 1 0 30016 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2031__A2
timestamp 1669390400
transform -1 0 30688 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2035__A1
timestamp 1669390400
transform 1 0 24640 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2037__A2
timestamp 1669390400
transform 1 0 36736 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2040__A2
timestamp 1669390400
transform 1 0 44352 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2041__A1
timestamp 1669390400
transform 1 0 45360 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2045__I
timestamp 1669390400
transform 1 0 61264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2046__A1
timestamp 1669390400
transform 1 0 44912 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2046__A2
timestamp 1669390400
transform 1 0 45360 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2050__A1
timestamp 1669390400
transform 1 0 33824 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2054__A1
timestamp 1669390400
transform -1 0 45472 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2056__A2
timestamp 1669390400
transform 1 0 38416 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2056__B
timestamp 1669390400
transform -1 0 36512 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2061__A1
timestamp 1669390400
transform 1 0 6048 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2063__A1
timestamp 1669390400
transform 1 0 38080 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2063__A2
timestamp 1669390400
transform -1 0 38752 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2064__A1
timestamp 1669390400
transform 1 0 38640 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2064__A2
timestamp 1669390400
transform -1 0 40208 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2067__A1
timestamp 1669390400
transform 1 0 29120 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2067__A2
timestamp 1669390400
transform 1 0 29568 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2070__A1
timestamp 1669390400
transform 1 0 33600 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2070__A2
timestamp 1669390400
transform -1 0 34272 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2071__A1
timestamp 1669390400
transform -1 0 33376 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2071__A2
timestamp 1669390400
transform 1 0 33488 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2074__A1
timestamp 1669390400
transform 1 0 36176 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2075__A2
timestamp 1669390400
transform 1 0 31472 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2077__A1
timestamp 1669390400
transform -1 0 21728 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2078__A2
timestamp 1669390400
transform 1 0 61264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2079__A1
timestamp 1669390400
transform -1 0 9408 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2080__A2
timestamp 1669390400
transform -1 0 9968 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2081__A1
timestamp 1669390400
transform 1 0 28336 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2081__A2
timestamp 1669390400
transform 1 0 27888 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2082__A1
timestamp 1669390400
transform -1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2083__A2
timestamp 1669390400
transform -1 0 12992 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2083__B2
timestamp 1669390400
transform -1 0 13440 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2084__A1
timestamp 1669390400
transform 1 0 26656 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2084__A2
timestamp 1669390400
transform -1 0 26432 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2085__A1
timestamp 1669390400
transform 1 0 27104 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2085__A2
timestamp 1669390400
transform 1 0 26320 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2086__A1
timestamp 1669390400
transform 1 0 27440 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2087__A2
timestamp 1669390400
transform -1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2091__A2
timestamp 1669390400
transform -1 0 58464 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2092__A1
timestamp 1669390400
transform 1 0 36848 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2092__A2
timestamp 1669390400
transform 1 0 37296 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2093__A1
timestamp 1669390400
transform 1 0 32256 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2093__A2
timestamp 1669390400
transform 1 0 37744 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2094__A2
timestamp 1669390400
transform 1 0 48720 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2095__A1
timestamp 1669390400
transform 1 0 43344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2095__A2
timestamp 1669390400
transform 1 0 42448 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2095__B1
timestamp 1669390400
transform 1 0 42896 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2095__B2
timestamp 1669390400
transform 1 0 42560 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2096__A1
timestamp 1669390400
transform 1 0 41440 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2096__B2
timestamp 1669390400
transform 1 0 40992 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2097__A1
timestamp 1669390400
transform 1 0 50624 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2097__A2
timestamp 1669390400
transform 1 0 50176 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2098__A1
timestamp 1669390400
transform -1 0 53984 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2098__A2
timestamp 1669390400
transform 1 0 57120 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2100__A2
timestamp 1669390400
transform -1 0 38752 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2102__A1
timestamp 1669390400
transform 1 0 31248 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2103__A1
timestamp 1669390400
transform -1 0 30240 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2104__A1
timestamp 1669390400
transform -1 0 33040 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2106__A2
timestamp 1669390400
transform 1 0 43008 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2110__I
timestamp 1669390400
transform 1 0 48272 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2111__A2
timestamp 1669390400
transform 1 0 43792 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2116__A1
timestamp 1669390400
transform -1 0 50736 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2117__A1
timestamp 1669390400
transform 1 0 45360 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2118__A1
timestamp 1669390400
transform 1 0 48048 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2122__A1
timestamp 1669390400
transform -1 0 47376 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2122__A2
timestamp 1669390400
transform -1 0 47824 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2128__A1
timestamp 1669390400
transform 1 0 48608 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2129__A2
timestamp 1669390400
transform 1 0 44800 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2131__A1
timestamp 1669390400
transform 1 0 35728 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2132__A1
timestamp 1669390400
transform 1 0 34048 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2137__A1
timestamp 1669390400
transform 1 0 43344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2138__A1
timestamp 1669390400
transform 1 0 46816 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2140__A1
timestamp 1669390400
transform 1 0 33824 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2144__A1
timestamp 1669390400
transform 1 0 35616 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2146__A2
timestamp 1669390400
transform -1 0 12096 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2148__I
timestamp 1669390400
transform 1 0 65296 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2149__A1
timestamp 1669390400
transform 1 0 37632 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2149__A2
timestamp 1669390400
transform -1 0 38080 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2149__B1
timestamp 1669390400
transform 1 0 39536 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2149__B2
timestamp 1669390400
transform -1 0 37632 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2150__A1
timestamp 1669390400
transform -1 0 39312 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2150__A2
timestamp 1669390400
transform 1 0 40880 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2153__A1
timestamp 1669390400
transform 1 0 30464 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2153__A2
timestamp 1669390400
transform 1 0 30240 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2155__A1
timestamp 1669390400
transform 1 0 34496 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2155__A2
timestamp 1669390400
transform -1 0 36064 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2156__A1
timestamp 1669390400
transform 1 0 35168 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2156__A2
timestamp 1669390400
transform 1 0 35840 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2159__A1
timestamp 1669390400
transform -1 0 37744 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2161__A1
timestamp 1669390400
transform -1 0 37744 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2163__A1
timestamp 1669390400
transform 1 0 31920 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2164__A1
timestamp 1669390400
transform -1 0 32032 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2165__A1
timestamp 1669390400
transform 1 0 29456 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2165__A2
timestamp 1669390400
transform 1 0 29904 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2166__A1
timestamp 1669390400
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2167__A1
timestamp 1669390400
transform 1 0 25760 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2168__A1
timestamp 1669390400
transform 1 0 36736 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2168__A2
timestamp 1669390400
transform 1 0 37408 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2169__A1
timestamp 1669390400
transform -1 0 34496 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2170__A1
timestamp 1669390400
transform 1 0 34160 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2170__B2
timestamp 1669390400
transform 1 0 37856 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2171__A1
timestamp 1669390400
transform 1 0 32256 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2171__A2
timestamp 1669390400
transform -1 0 33264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2172__A1
timestamp 1669390400
transform 1 0 26992 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2172__A2
timestamp 1669390400
transform 1 0 29456 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2173__A2
timestamp 1669390400
transform -1 0 29680 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2177__A2
timestamp 1669390400
transform 1 0 38080 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2179__A1
timestamp 1669390400
transform 1 0 33824 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2179__A2
timestamp 1669390400
transform 1 0 34272 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2180__A1
timestamp 1669390400
transform -1 0 34944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2180__A2
timestamp 1669390400
transform -1 0 35840 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2182__A1
timestamp 1669390400
transform 1 0 57568 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2182__A2
timestamp 1669390400
transform 1 0 58016 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2183__I
timestamp 1669390400
transform 1 0 60368 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2184__A1
timestamp 1669390400
transform 1 0 43456 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2184__A2
timestamp 1669390400
transform 1 0 46816 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2184__B1
timestamp 1669390400
transform 1 0 44688 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2184__B2
timestamp 1669390400
transform 1 0 47264 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2185__A1
timestamp 1669390400
transform -1 0 45472 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2186__A1
timestamp 1669390400
transform 1 0 55552 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2186__A2
timestamp 1669390400
transform 1 0 53312 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2187__A1
timestamp 1669390400
transform -1 0 52192 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2187__A2
timestamp 1669390400
transform 1 0 56672 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2192__A1
timestamp 1669390400
transform -1 0 38752 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2193__A1
timestamp 1669390400
transform -1 0 38640 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2195__A1
timestamp 1669390400
transform 1 0 42896 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2196__A2
timestamp 1669390400
transform -1 0 45920 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2202__A1
timestamp 1669390400
transform 1 0 41888 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2203__A2
timestamp 1669390400
transform 1 0 45360 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2203__B
timestamp 1669390400
transform 1 0 44464 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2204__A1
timestamp 1669390400
transform 1 0 37184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2207__A2
timestamp 1669390400
transform 1 0 44688 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2208__A1
timestamp 1669390400
transform 1 0 39088 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2210__A1
timestamp 1669390400
transform 1 0 39648 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2214__A1
timestamp 1669390400
transform -1 0 37184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2214__A2
timestamp 1669390400
transform 1 0 36736 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2216__A1
timestamp 1669390400
transform 1 0 50736 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2216__A2
timestamp 1669390400
transform 1 0 53312 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2217__A1
timestamp 1669390400
transform 1 0 49392 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2217__A2
timestamp 1669390400
transform 1 0 48944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2217__A3
timestamp 1669390400
transform 1 0 50624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2217__A4
timestamp 1669390400
transform 1 0 50288 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2218__A1
timestamp 1669390400
transform 1 0 50624 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2218__A2
timestamp 1669390400
transform 1 0 52304 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2218__B1
timestamp 1669390400
transform 1 0 52304 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2218__B2
timestamp 1669390400
transform 1 0 51520 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2221__A2
timestamp 1669390400
transform 1 0 42112 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2222__A2
timestamp 1669390400
transform 1 0 41552 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2224__A1
timestamp 1669390400
transform 1 0 39312 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2225__A1
timestamp 1669390400
transform 1 0 29456 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2225__A2
timestamp 1669390400
transform 1 0 29904 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2227__A1
timestamp 1669390400
transform 1 0 34944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2227__A2
timestamp 1669390400
transform -1 0 36960 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2230__A1
timestamp 1669390400
transform 1 0 34944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2230__A2
timestamp 1669390400
transform 1 0 36176 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2231__A1
timestamp 1669390400
transform 1 0 30240 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2231__A2
timestamp 1669390400
transform 1 0 30912 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2232__A2
timestamp 1669390400
transform -1 0 31136 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2235__A1
timestamp 1669390400
transform 1 0 41440 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2238__A1
timestamp 1669390400
transform 1 0 39536 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2238__A2
timestamp 1669390400
transform 1 0 39984 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2239__A1
timestamp 1669390400
transform -1 0 35392 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2239__A2
timestamp 1669390400
transform 1 0 37856 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2240__A3
timestamp 1669390400
transform 1 0 40656 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2241__A1
timestamp 1669390400
transform 1 0 52864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2241__A2
timestamp 1669390400
transform 1 0 52416 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2242__A1
timestamp 1669390400
transform 1 0 48272 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2242__A2
timestamp 1669390400
transform 1 0 47376 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2242__B1
timestamp 1669390400
transform 1 0 47824 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2242__B2
timestamp 1669390400
transform 1 0 45360 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2244__A1
timestamp 1669390400
transform 1 0 51968 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2244__A2
timestamp 1669390400
transform 1 0 52080 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2245__A1
timestamp 1669390400
transform 1 0 59696 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2245__A2
timestamp 1669390400
transform 1 0 59248 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2251__A1
timestamp 1669390400
transform -1 0 42672 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2258__A1
timestamp 1669390400
transform 1 0 47264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2274__A2
timestamp 1669390400
transform 1 0 44912 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2277__A1
timestamp 1669390400
transform 1 0 42448 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2278__A1
timestamp 1669390400
transform 1 0 44576 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2280__A1
timestamp 1669390400
transform 1 0 43568 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2283__A1
timestamp 1669390400
transform -1 0 45584 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2284__A1
timestamp 1669390400
transform 1 0 45584 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2286__I
timestamp 1669390400
transform 1 0 40992 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2289__A1
timestamp 1669390400
transform 1 0 51184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2289__A2
timestamp 1669390400
transform 1 0 51632 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2290__A1
timestamp 1669390400
transform 1 0 47264 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2290__A2
timestamp 1669390400
transform 1 0 49840 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2291__A1
timestamp 1669390400
transform 1 0 53648 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2291__A2
timestamp 1669390400
transform 1 0 54992 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2292__A2
timestamp 1669390400
transform -1 0 52080 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2296__A1
timestamp 1669390400
transform 1 0 52640 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2297__A1
timestamp 1669390400
transform -1 0 53200 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2300__A1
timestamp 1669390400
transform 1 0 57904 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2300__A2
timestamp 1669390400
transform 1 0 58352 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2301__A1
timestamp 1669390400
transform -1 0 42784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2301__A2
timestamp 1669390400
transform 1 0 43904 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2304__A1
timestamp 1669390400
transform 1 0 37408 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2304__A2
timestamp 1669390400
transform 1 0 38304 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2305__A2
timestamp 1669390400
transform 1 0 40544 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2306__A2
timestamp 1669390400
transform 1 0 42112 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2307__A1
timestamp 1669390400
transform 1 0 55888 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2307__A2
timestamp 1669390400
transform 1 0 56896 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2308__A1
timestamp 1669390400
transform 1 0 69216 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2309__A1
timestamp 1669390400
transform 1 0 58016 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2309__A2
timestamp 1669390400
transform 1 0 58464 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2311__A1
timestamp 1669390400
transform 1 0 54992 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2312__A1
timestamp 1669390400
transform 1 0 50960 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2315__A1
timestamp 1669390400
transform 1 0 51520 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2315__A2
timestamp 1669390400
transform 1 0 50288 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2316__A1
timestamp 1669390400
transform 1 0 43568 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2316__A2
timestamp 1669390400
transform 1 0 44016 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2317__A1
timestamp 1669390400
transform 1 0 48720 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2317__A3
timestamp 1669390400
transform 1 0 49952 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2318__A1
timestamp 1669390400
transform 1 0 53312 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2318__A2
timestamp 1669390400
transform 1 0 53760 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2319__I
timestamp 1669390400
transform -1 0 55552 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2320__I
timestamp 1669390400
transform 1 0 55552 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2321__A1
timestamp 1669390400
transform 1 0 49728 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2321__A2
timestamp 1669390400
transform 1 0 50960 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2321__B1
timestamp 1669390400
transform 1 0 50960 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2321__B2
timestamp 1669390400
transform 1 0 49280 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2322__B1
timestamp 1669390400
transform 1 0 52528 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2323__A1
timestamp 1669390400
transform 1 0 57344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2323__A2
timestamp 1669390400
transform 1 0 57792 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2324__A1
timestamp 1669390400
transform 1 0 59136 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2324__A2
timestamp 1669390400
transform 1 0 58688 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2343__A1
timestamp 1669390400
transform 1 0 56112 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2344__A1
timestamp 1669390400
transform 1 0 54880 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2348__A1
timestamp 1669390400
transform 1 0 54768 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2349__A1
timestamp 1669390400
transform 1 0 52416 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2350__A1
timestamp 1669390400
transform 1 0 60592 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2350__A2
timestamp 1669390400
transform 1 0 62272 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2350__B1
timestamp 1669390400
transform -1 0 62048 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2350__B2
timestamp 1669390400
transform -1 0 61376 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2351__A1
timestamp 1669390400
transform 1 0 60256 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2351__A2
timestamp 1669390400
transform 1 0 60704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2351__A3
timestamp 1669390400
transform 1 0 62608 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2351__A4
timestamp 1669390400
transform 1 0 63056 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2352__A2
timestamp 1669390400
transform 1 0 63616 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2353__A2
timestamp 1669390400
transform 1 0 54544 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2354__A2
timestamp 1669390400
transform 1 0 57344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2357__A1
timestamp 1669390400
transform 1 0 62384 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2362__A1
timestamp 1669390400
transform 1 0 68432 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2363__A1
timestamp 1669390400
transform 1 0 55776 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2363__A2
timestamp 1669390400
transform -1 0 58464 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2366__A1
timestamp 1669390400
transform 1 0 49616 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2366__A2
timestamp 1669390400
transform 1 0 49168 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2367__A1
timestamp 1669390400
transform 1 0 49392 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2367__A2
timestamp 1669390400
transform 1 0 49168 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2368__A1
timestamp 1669390400
transform 1 0 52304 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2368__A2
timestamp 1669390400
transform -1 0 49616 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2369__A1
timestamp 1669390400
transform 1 0 66976 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2369__A2
timestamp 1669390400
transform -1 0 66304 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2370__A1
timestamp 1669390400
transform 1 0 66752 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2370__A2
timestamp 1669390400
transform 1 0 69552 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2371__A1
timestamp 1669390400
transform 1 0 68320 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2373__A1
timestamp 1669390400
transform 1 0 64736 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2377__A1
timestamp 1669390400
transform 1 0 60592 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2377__A2
timestamp 1669390400
transform -1 0 59808 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2378__A1
timestamp 1669390400
transform 1 0 54208 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2378__A2
timestamp 1669390400
transform 1 0 53536 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2378__B1
timestamp 1669390400
transform 1 0 53760 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2378__B2
timestamp 1669390400
transform 1 0 53536 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2380__A1
timestamp 1669390400
transform 1 0 60032 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2380__A2
timestamp 1669390400
transform 1 0 60480 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2381__A2
timestamp 1669390400
transform 1 0 64848 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2384__A1
timestamp 1669390400
transform 1 0 62832 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2384__A2
timestamp 1669390400
transform 1 0 62496 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2385__A1
timestamp 1669390400
transform 1 0 65744 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2385__A2
timestamp 1669390400
transform 1 0 65744 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2386__A1
timestamp 1669390400
transform 1 0 58800 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2386__A2
timestamp 1669390400
transform -1 0 61152 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2390__A1
timestamp 1669390400
transform -1 0 59024 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2408__A2
timestamp 1669390400
transform 1 0 54880 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2411__A2
timestamp 1669390400
transform 1 0 54208 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2416__A1
timestamp 1669390400
transform 1 0 61936 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2418__A1
timestamp 1669390400
transform -1 0 60592 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2421__A1
timestamp 1669390400
transform 1 0 63952 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2423__A1
timestamp 1669390400
transform 1 0 65296 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2423__A2
timestamp 1669390400
transform -1 0 65968 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2423__A3
timestamp 1669390400
transform 1 0 64288 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2424__A1
timestamp 1669390400
transform 1 0 65296 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2431__A2
timestamp 1669390400
transform 1 0 64624 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2432__A1
timestamp 1669390400
transform 1 0 60144 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2432__A2
timestamp 1669390400
transform 1 0 57792 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2432__B1
timestamp 1669390400
transform 1 0 57344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2432__B2
timestamp 1669390400
transform 1 0 55216 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2434__A2
timestamp 1669390400
transform -1 0 64736 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2435__A1
timestamp 1669390400
transform -1 0 59584 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2435__A2
timestamp 1669390400
transform -1 0 59136 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2436__A3
timestamp 1669390400
transform -1 0 70336 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2437__A1
timestamp 1669390400
transform 1 0 78064 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2437__A2
timestamp 1669390400
transform 1 0 77616 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2438__A1
timestamp 1669390400
transform 1 0 68432 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2438__A2
timestamp 1669390400
transform 1 0 70560 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2439__A1
timestamp 1669390400
transform 1 0 66976 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2439__A2
timestamp 1669390400
transform -1 0 64400 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2440__A1
timestamp 1669390400
transform 1 0 70560 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2440__A2
timestamp 1669390400
transform 1 0 69216 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2444__A1
timestamp 1669390400
transform -1 0 75600 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2445__A1
timestamp 1669390400
transform 1 0 69776 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2445__A2
timestamp 1669390400
transform 1 0 72240 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2446__A1
timestamp 1669390400
transform 1 0 70000 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2449__A1
timestamp 1669390400
transform 1 0 63504 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2450__A1
timestamp 1669390400
transform 1 0 74032 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2450__A2
timestamp 1669390400
transform 1 0 73808 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2451__A1
timestamp 1669390400
transform 1 0 73696 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2451__A2
timestamp 1669390400
transform 1 0 72240 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2454__A1
timestamp 1669390400
transform 1 0 75824 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2457__A2
timestamp 1669390400
transform 1 0 69216 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2467__A1
timestamp 1669390400
transform 1 0 63840 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2467__A2
timestamp 1669390400
transform 1 0 63392 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2467__A3
timestamp 1669390400
transform -1 0 63168 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2467__A4
timestamp 1669390400
transform -1 0 64512 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2469__A2
timestamp 1669390400
transform -1 0 68880 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2472__A1
timestamp 1669390400
transform 1 0 77504 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2474__A1
timestamp 1669390400
transform -1 0 75488 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2475__A1
timestamp 1669390400
transform 1 0 77840 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2477__A1
timestamp 1669390400
transform -1 0 74256 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2477__A2
timestamp 1669390400
transform -1 0 74816 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2479__A2
timestamp 1669390400
transform -1 0 60032 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2480__A1
timestamp 1669390400
transform 1 0 63392 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2480__A2
timestamp 1669390400
transform 1 0 61376 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2480__B1
timestamp 1669390400
transform 1 0 64400 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2481__A2
timestamp 1669390400
transform -1 0 63952 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2482__A1
timestamp 1669390400
transform 1 0 69664 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2482__A2
timestamp 1669390400
transform -1 0 65520 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2483__A1
timestamp 1669390400
transform 1 0 63840 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2483__A2
timestamp 1669390400
transform 1 0 64176 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2484__A1
timestamp 1669390400
transform 1 0 74032 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2484__A3
timestamp 1669390400
transform 1 0 74368 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2485__A1
timestamp 1669390400
transform -1 0 73920 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2486__A1
timestamp 1669390400
transform 1 0 69776 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2486__A2
timestamp 1669390400
transform 1 0 70224 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2487__A1
timestamp 1669390400
transform 1 0 73472 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2487__A2
timestamp 1669390400
transform 1 0 73584 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2488__A1
timestamp 1669390400
transform 1 0 66304 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2488__A2
timestamp 1669390400
transform -1 0 68208 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2489__A3
timestamp 1669390400
transform 1 0 73136 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2495__A1
timestamp 1669390400
transform 1 0 73248 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2496__A1
timestamp 1669390400
transform 1 0 70448 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2496__A2
timestamp 1669390400
transform 1 0 70896 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2497__A1
timestamp 1669390400
transform -1 0 69552 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2497__A2
timestamp 1669390400
transform 1 0 70784 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2498__A2
timestamp 1669390400
transform 1 0 69552 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2499__A1
timestamp 1669390400
transform 1 0 69776 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2499__A2
timestamp 1669390400
transform 1 0 72352 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2513__A2
timestamp 1669390400
transform -1 0 55104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2519__A1
timestamp 1669390400
transform 1 0 78064 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2530__A1
timestamp 1669390400
transform 1 0 74144 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2532__A1
timestamp 1669390400
transform 1 0 64624 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2532__A2
timestamp 1669390400
transform 1 0 66864 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2533__A1
timestamp 1669390400
transform 1 0 73248 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2533__A2
timestamp 1669390400
transform -1 0 72464 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2534__A1
timestamp 1669390400
transform 1 0 72576 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2534__A2
timestamp 1669390400
transform 1 0 73024 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2535__A1
timestamp 1669390400
transform 1 0 66528 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2535__A2
timestamp 1669390400
transform 1 0 66080 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2536__A1
timestamp 1669390400
transform -1 0 59920 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2536__A2
timestamp 1669390400
transform 1 0 58576 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2537__A1
timestamp 1669390400
transform 1 0 64848 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2537__A2
timestamp 1669390400
transform 1 0 67984 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2537__A3
timestamp 1669390400
transform 1 0 64176 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2538__A1
timestamp 1669390400
transform 1 0 71680 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2539__A1
timestamp 1669390400
transform 1 0 66080 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2539__A2
timestamp 1669390400
transform 1 0 64624 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2540__A1
timestamp 1669390400
transform 1 0 65744 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2540__A2
timestamp 1669390400
transform 1 0 67760 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2541__A1
timestamp 1669390400
transform 1 0 67872 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2541__A2
timestamp 1669390400
transform 1 0 68320 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2542__A1
timestamp 1669390400
transform -1 0 64848 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2544__A1
timestamp 1669390400
transform 1 0 74032 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2545__A1
timestamp 1669390400
transform 1 0 71232 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2545__A2
timestamp 1669390400
transform 1 0 70784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2547__A2
timestamp 1669390400
transform 1 0 73248 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2548__A2
timestamp 1669390400
transform 1 0 70672 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2549__A1
timestamp 1669390400
transform 1 0 67760 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2549__A2
timestamp 1669390400
transform 1 0 68208 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2551__A1
timestamp 1669390400
transform 1 0 70784 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2554__A1
timestamp 1669390400
transform 1 0 77952 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2555__A1
timestamp 1669390400
transform -1 0 73584 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2560__A2
timestamp 1669390400
transform 1 0 63056 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2565__A1
timestamp 1669390400
transform 1 0 77952 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2566__A1
timestamp 1669390400
transform -1 0 74032 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2567__I
timestamp 1669390400
transform 1 0 70336 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2571__A1
timestamp 1669390400
transform 1 0 74480 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2573__A1
timestamp 1669390400
transform 1 0 68544 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2575__A1
timestamp 1669390400
transform 1 0 60592 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2575__A2
timestamp 1669390400
transform 1 0 59472 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2576__A1
timestamp 1669390400
transform -1 0 63280 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2576__A2
timestamp 1669390400
transform -1 0 63728 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2577__A1
timestamp 1669390400
transform 1 0 66640 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2577__A2
timestamp 1669390400
transform 1 0 65744 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2577__B2
timestamp 1669390400
transform 1 0 67088 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2578__A1
timestamp 1669390400
transform 1 0 60256 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2578__A2
timestamp 1669390400
transform 1 0 60704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2579__A1
timestamp 1669390400
transform 1 0 56784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2579__A2
timestamp 1669390400
transform 1 0 60368 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2580__A1
timestamp 1669390400
transform 1 0 61264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2581__A1
timestamp 1669390400
transform -1 0 70672 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2582__A1
timestamp 1669390400
transform 1 0 63168 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2582__A2
timestamp 1669390400
transform 1 0 65296 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2583__A1
timestamp 1669390400
transform 1 0 63728 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2583__A2
timestamp 1669390400
transform 1 0 64176 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2584__A1
timestamp 1669390400
transform 1 0 66976 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2584__A2
timestamp 1669390400
transform 1 0 64736 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2588__A1
timestamp 1669390400
transform -1 0 67536 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2589__A1
timestamp 1669390400
transform 1 0 67872 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2590__A1
timestamp 1669390400
transform 1 0 68992 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2590__A2
timestamp 1669390400
transform 1 0 72688 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2590__A3
timestamp 1669390400
transform 1 0 69664 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2594__A1
timestamp 1669390400
transform 1 0 74368 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2597__A1
timestamp 1669390400
transform 1 0 77056 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2601__A2
timestamp 1669390400
transform 1 0 74480 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2602__A1
timestamp 1669390400
transform 1 0 67312 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2602__A2
timestamp 1669390400
transform 1 0 67760 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2605__B
timestamp 1669390400
transform 1 0 56000 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2606__C
timestamp 1669390400
transform -1 0 52528 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2608__B2
timestamp 1669390400
transform 1 0 63840 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2609__A1
timestamp 1669390400
transform 1 0 62608 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2609__A2
timestamp 1669390400
transform 1 0 59696 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2609__A3
timestamp 1669390400
transform 1 0 64288 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2612__I
timestamp 1669390400
transform 1 0 68768 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2613__A2
timestamp 1669390400
transform 1 0 68208 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2615__A1
timestamp 1669390400
transform 1 0 60592 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2615__A2
timestamp 1669390400
transform 1 0 60144 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2615__A3
timestamp 1669390400
transform 1 0 63840 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2616__I
timestamp 1669390400
transform -1 0 68768 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2617__B
timestamp 1669390400
transform -1 0 69552 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2617__C
timestamp 1669390400
transform 1 0 69776 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2621__A1
timestamp 1669390400
transform 1 0 63392 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2621__A2
timestamp 1669390400
transform 1 0 63840 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2624__A1
timestamp 1669390400
transform 1 0 70560 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2626__A1
timestamp 1669390400
transform 1 0 56896 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2626__A2
timestamp 1669390400
transform 1 0 58128 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2627__A1
timestamp 1669390400
transform -1 0 60032 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2628__A1
timestamp 1669390400
transform 1 0 59920 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2629__A1
timestamp 1669390400
transform 1 0 59024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2629__A2
timestamp 1669390400
transform 1 0 60144 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2630__A1
timestamp 1669390400
transform 1 0 59024 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2630__A2
timestamp 1669390400
transform 1 0 56448 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2634__A1
timestamp 1669390400
transform 1 0 67424 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2634__A2
timestamp 1669390400
transform 1 0 67872 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2635__A1
timestamp 1669390400
transform 1 0 67312 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2635__A2
timestamp 1669390400
transform 1 0 67760 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2638__A1
timestamp 1669390400
transform 1 0 69776 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2640__A1
timestamp 1669390400
transform 1 0 76832 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2644__A1
timestamp 1669390400
transform 1 0 73248 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2645__A2
timestamp 1669390400
transform 1 0 77840 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2646__A2
timestamp 1669390400
transform -1 0 77728 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2646__B
timestamp 1669390400
transform -1 0 74256 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2648__I
timestamp 1669390400
transform 1 0 67200 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2652__A2
timestamp 1669390400
transform -1 0 76832 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2660__A1
timestamp 1669390400
transform 1 0 68992 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2661__A1
timestamp 1669390400
transform 1 0 63280 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2661__A2
timestamp 1669390400
transform 1 0 64624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2661__B1
timestamp 1669390400
transform 1 0 64176 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2661__B2
timestamp 1669390400
transform -1 0 63952 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2662__A1
timestamp 1669390400
transform 1 0 64624 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2662__A2
timestamp 1669390400
transform 1 0 65968 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2666__A1
timestamp 1669390400
transform 1 0 59920 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2666__A2
timestamp 1669390400
transform 1 0 59472 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2668__A1
timestamp 1669390400
transform 1 0 58800 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2668__A2
timestamp 1669390400
transform 1 0 59808 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2669__A1
timestamp 1669390400
transform 1 0 57344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2669__A2
timestamp 1669390400
transform 1 0 55888 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2671__A1
timestamp 1669390400
transform 1 0 59024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2671__A2
timestamp 1669390400
transform 1 0 56224 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2671__B1
timestamp 1669390400
transform 1 0 56672 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2671__B2
timestamp 1669390400
transform 1 0 58576 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2680__A1
timestamp 1669390400
transform 1 0 74032 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2685__A1
timestamp 1669390400
transform 1 0 77952 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2687__A2
timestamp 1669390400
transform 1 0 74144 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2688__A1
timestamp 1669390400
transform -1 0 76720 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2698__A1
timestamp 1669390400
transform 1 0 60256 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2698__A2
timestamp 1669390400
transform 1 0 60704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2699__A1
timestamp 1669390400
transform -1 0 56336 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2699__A2
timestamp 1669390400
transform 1 0 55776 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2710__A2
timestamp 1669390400
transform 1 0 72016 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2721__A1
timestamp 1669390400
transform 1 0 72016 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2725__A1
timestamp 1669390400
transform -1 0 53536 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2725__A2
timestamp 1669390400
transform 1 0 55328 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2726__A1
timestamp 1669390400
transform 1 0 53536 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2726__A2
timestamp 1669390400
transform 1 0 53760 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2727__A1
timestamp 1669390400
transform -1 0 56784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2727__A2
timestamp 1669390400
transform 1 0 56224 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2735__A1
timestamp 1669390400
transform 1 0 60368 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2735__A2
timestamp 1669390400
transform 1 0 60816 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2739__I
timestamp 1669390400
transform 1 0 62496 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2748__A1
timestamp 1669390400
transform 1 0 68544 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2751__A2
timestamp 1669390400
transform 1 0 70000 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2751__A3
timestamp 1669390400
transform 1 0 72688 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2760__A1
timestamp 1669390400
transform 1 0 51744 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2760__A2
timestamp 1669390400
transform 1 0 52192 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2763__A1
timestamp 1669390400
transform -1 0 52864 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2763__A2
timestamp 1669390400
transform -1 0 52416 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2774__A2
timestamp 1669390400
transform 1 0 71792 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2779__A1
timestamp 1669390400
transform 1 0 57232 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2779__A2
timestamp 1669390400
transform 1 0 56336 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2784__A1
timestamp 1669390400
transform -1 0 55440 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2785__A1
timestamp 1669390400
transform 1 0 57568 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2791__A1
timestamp 1669390400
transform -1 0 63952 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2795__A1
timestamp 1669390400
transform 1 0 67088 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2796__A1
timestamp 1669390400
transform 1 0 57680 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2796__A2
timestamp 1669390400
transform 1 0 59248 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2797__A1
timestamp 1669390400
transform 1 0 58240 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2797__A2
timestamp 1669390400
transform -1 0 59248 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2801__A2
timestamp 1669390400
transform -1 0 18816 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2804__A1
timestamp 1669390400
transform 1 0 23408 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2804__A2
timestamp 1669390400
transform 1 0 25200 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2804__B1
timestamp 1669390400
transform 1 0 24192 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2804__B2
timestamp 1669390400
transform 1 0 21504 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2806__CLK
timestamp 1669390400
transform 1 0 5600 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2807__I
timestamp 1669390400
transform 1 0 74928 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2808__I
timestamp 1669390400
transform 1 0 77952 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2809__I
timestamp 1669390400
transform 1 0 77952 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2810__I
timestamp 1669390400
transform 1 0 77616 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2811__I
timestamp 1669390400
transform 1 0 78064 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2812__I
timestamp 1669390400
transform -1 0 73696 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2813__I
timestamp 1669390400
transform 1 0 78064 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2814__I
timestamp 1669390400
transform 1 0 77952 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2815__I
timestamp 1669390400
transform 1 0 73248 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2816__I
timestamp 1669390400
transform 1 0 78064 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2817__I
timestamp 1669390400
transform -1 0 74032 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2818__I
timestamp 1669390400
transform 1 0 77952 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2819__I
timestamp 1669390400
transform 1 0 75600 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2820__I
timestamp 1669390400
transform 1 0 74032 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2821__I
timestamp 1669390400
transform -1 0 72464 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2822__I
timestamp 1669390400
transform 1 0 71680 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2823__I
timestamp 1669390400
transform -1 0 4592 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2824__I
timestamp 1669390400
transform 1 0 4816 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2825__I
timestamp 1669390400
transform -1 0 2576 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2826__I
timestamp 1669390400
transform -1 0 2352 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2827__I
timestamp 1669390400
transform -1 0 2016 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2828__I
timestamp 1669390400
transform -1 0 2464 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2829__I
timestamp 1669390400
transform -1 0 2352 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2830__I
timestamp 1669390400
transform -1 0 4704 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2831__I
timestamp 1669390400
transform -1 0 2464 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2832__I
timestamp 1669390400
transform 1 0 3472 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2833__I
timestamp 1669390400
transform 1 0 3584 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2834__I
timestamp 1669390400
transform 1 0 3584 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2835__I
timestamp 1669390400
transform 1 0 3584 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2836__I
timestamp 1669390400
transform 1 0 4368 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2837__I
timestamp 1669390400
transform 1 0 4816 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2838__I
timestamp 1669390400
transform 1 0 5264 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1669390400
transform -1 0 8736 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1669390400
transform -1 0 31696 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1669390400
transform -1 0 32592 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1669390400
transform -1 0 36064 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1669390400
transform -1 0 37856 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1669390400
transform 1 0 42000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1669390400
transform -1 0 43232 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1669390400
transform -1 0 11648 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1669390400
transform 1 0 19936 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1669390400
transform 1 0 17920 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input11_I
timestamp 1669390400
transform -1 0 18032 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input12_I
timestamp 1669390400
transform -1 0 21056 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input13_I
timestamp 1669390400
transform 1 0 25088 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input14_I
timestamp 1669390400
transform -1 0 23632 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input15_I
timestamp 1669390400
transform -1 0 25984 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input16_I
timestamp 1669390400
transform -1 0 28672 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input17_I
timestamp 1669390400
transform 1 0 51744 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input18_I
timestamp 1669390400
transform 1 0 73920 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input19_I
timestamp 1669390400
transform 1 0 77280 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input20_I
timestamp 1669390400
transform 1 0 77728 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input21_I
timestamp 1669390400
transform 1 0 77168 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input22_I
timestamp 1669390400
transform -1 0 74592 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input23_I
timestamp 1669390400
transform -1 0 74704 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input24_I
timestamp 1669390400
transform 1 0 53760 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input25_I
timestamp 1669390400
transform 1 0 53312 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input26_I
timestamp 1669390400
transform -1 0 52640 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input27_I
timestamp 1669390400
transform 1 0 61264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input28_I
timestamp 1669390400
transform -1 0 56000 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input29_I
timestamp 1669390400
transform 1 0 65632 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input30_I
timestamp 1669390400
transform 1 0 68320 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input31_I
timestamp 1669390400
transform 1 0 68208 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input32_I
timestamp 1669390400
transform -1 0 64624 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input33_I
timestamp 1669390400
transform -1 0 6832 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output34_I
timestamp 1669390400
transform 1 0 6048 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output35_I
timestamp 1669390400
transform 1 0 27888 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output36_I
timestamp 1669390400
transform -1 0 28672 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output37_I
timestamp 1669390400
transform 1 0 32592 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output38_I
timestamp 1669390400
transform -1 0 33600 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output39_I
timestamp 1669390400
transform 1 0 38080 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output40_I
timestamp 1669390400
transform 1 0 40544 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output41_I
timestamp 1669390400
transform 1 0 43008 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output42_I
timestamp 1669390400
transform 1 0 45360 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output43_I
timestamp 1669390400
transform 1 0 47936 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output44_I
timestamp 1669390400
transform 1 0 49168 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output45_I
timestamp 1669390400
transform 1 0 5600 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output46_I
timestamp 1669390400
transform 1 0 52528 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output47_I
timestamp 1669390400
transform 1 0 53312 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output48_I
timestamp 1669390400
transform 1 0 58128 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output49_I
timestamp 1669390400
transform 1 0 60480 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output50_I
timestamp 1669390400
transform 1 0 61264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output51_I
timestamp 1669390400
transform 1 0 67872 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output52_I
timestamp 1669390400
transform 1 0 68320 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output53_I
timestamp 1669390400
transform 1 0 68992 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output54_I
timestamp 1669390400
transform 1 0 71232 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output55_I
timestamp 1669390400
transform -1 0 73248 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output56_I
timestamp 1669390400
transform 1 0 8512 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output57_I
timestamp 1669390400
transform -1 0 74368 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output58_I
timestamp 1669390400
transform -1 0 74480 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output59_I
timestamp 1669390400
transform 1 0 10416 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output60_I
timestamp 1669390400
transform 1 0 12320 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output61_I
timestamp 1669390400
transform 1 0 13664 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output62_I
timestamp 1669390400
transform -1 0 14448 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output63_I
timestamp 1669390400
transform -1 0 15904 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output64_I
timestamp 1669390400
transform 1 0 21840 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output65_I
timestamp 1669390400
transform 1 0 25200 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output68_I
timestamp 1669390400
transform 1 0 78064 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output76_I
timestamp 1669390400
transform 1 0 77392 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output77_I
timestamp 1669390400
transform 1 0 77840 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output78_I
timestamp 1669390400
transform -1 0 74592 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output79_I
timestamp 1669390400
transform -1 0 75600 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output80_I
timestamp 1669390400
transform -1 0 77392 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output81_I
timestamp 1669390400
transform 1 0 74368 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output82_I
timestamp 1669390400
transform -1 0 77392 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output97_I
timestamp 1669390400
transform 1 0 6496 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2 Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 1568 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4 Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 1792 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34
timestamp 1669390400
transform 1 0 5152 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37
timestamp 1669390400
transform 1 0 5488 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40 Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 5824 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44
timestamp 1669390400
transform 1 0 6272 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46
timestamp 1669390400
transform 1 0 6496 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49
timestamp 1669390400
transform 1 0 6832 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67
timestamp 1669390400
transform 1 0 8848 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69
timestamp 1669390400
transform 1 0 9072 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72
timestamp 1669390400
transform 1 0 9408 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_87
timestamp 1669390400
transform 1 0 11088 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_97
timestamp 1669390400
transform 1 0 12208 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_101
timestamp 1669390400
transform 1 0 12656 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_104
timestamp 1669390400
transform 1 0 12992 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_107
timestamp 1669390400
transform 1 0 13328 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_116
timestamp 1669390400
transform 1 0 14336 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_130
timestamp 1669390400
transform 1 0 15904 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_138
timestamp 1669390400
transform 1 0 16800 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_142
timestamp 1669390400
transform 1 0 17248 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_145
timestamp 1669390400
transform 1 0 17584 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_149
timestamp 1669390400
transform 1 0 18032 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_159
timestamp 1669390400
transform 1 0 19152 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_173
timestamp 1669390400
transform 1 0 20720 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_177
timestamp 1669390400
transform 1 0 21168 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_179
timestamp 1669390400
transform 1 0 21392 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_182
timestamp 1669390400
transform 1 0 21728 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_192
timestamp 1669390400
transform 1 0 22848 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_196
timestamp 1669390400
transform 1 0 23296 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_199
timestamp 1669390400
transform 1 0 23632 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_209
timestamp 1669390400
transform 1 0 24752 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_212
timestamp 1669390400
transform 1 0 25088 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_216
timestamp 1669390400
transform 1 0 25536 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_220
timestamp 1669390400
transform 1 0 25984 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_228
timestamp 1669390400
transform 1 0 26880 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_232
timestamp 1669390400
transform 1 0 27328 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_236
timestamp 1669390400
transform 1 0 27776 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_240
timestamp 1669390400
transform 1 0 28224 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_244
timestamp 1669390400
transform 1 0 28672 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_247
timestamp 1669390400
transform 1 0 29008 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_254
timestamp 1669390400
transform 1 0 29792 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_258
timestamp 1669390400
transform 1 0 30240 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_266
timestamp 1669390400
transform 1 0 31136 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_268
timestamp 1669390400
transform 1 0 31360 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_271
timestamp 1669390400
transform 1 0 31696 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_275
timestamp 1669390400
transform 1 0 32144 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_279
timestamp 1669390400
transform 1 0 32592 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_282
timestamp 1669390400
transform 1 0 32928 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_289
timestamp 1669390400
transform 1 0 33712 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_296
timestamp 1669390400
transform 1 0 34496 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_304
timestamp 1669390400
transform 1 0 35392 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_310
timestamp 1669390400
transform 1 0 36064 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_314
timestamp 1669390400
transform 1 0 36512 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_317
timestamp 1669390400
transform 1 0 36848 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_324
timestamp 1669390400
transform 1 0 37632 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_330
timestamp 1669390400
transform 1 0 38304 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_334
timestamp 1669390400
transform 1 0 38752 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_342
timestamp 1669390400
transform 1 0 39648 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_349
timestamp 1669390400
transform 1 0 40432 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_352
timestamp 1669390400
transform 1 0 40768 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_354
timestamp 1669390400
transform 1 0 40992 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_361
timestamp 1669390400
transform 1 0 41776 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_365
timestamp 1669390400
transform 1 0 42224 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_374
timestamp 1669390400
transform 1 0 43232 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_384
timestamp 1669390400
transform 1 0 44352 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_387
timestamp 1669390400
transform 1 0 44688 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_398
timestamp 1669390400
transform 1 0 45920 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_408
timestamp 1669390400
transform 1 0 47040 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_418
timestamp 1669390400
transform 1 0 48160 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_422
timestamp 1669390400
transform 1 0 48608 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_448
timestamp 1669390400
transform 1 0 51520 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_452
timestamp 1669390400
transform 1 0 51968 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_454
timestamp 1669390400
transform 1 0 52192 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_457
timestamp 1669390400
transform 1 0 52528 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_466
timestamp 1669390400
transform 1 0 53536 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_476
timestamp 1669390400
transform 1 0 54656 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_486
timestamp 1669390400
transform 1 0 55776 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_492
timestamp 1669390400
transform 1 0 56448 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_498
timestamp 1669390400
transform 1 0 57120 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_508
timestamp 1669390400
transform 1 0 58240 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_516
timestamp 1669390400
transform 1 0 59136 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_523
timestamp 1669390400
transform 1 0 59920 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_527
timestamp 1669390400
transform 1 0 60368 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_553
timestamp 1669390400
transform 1 0 63280 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_557
timestamp 1669390400
transform 1 0 63728 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_559
timestamp 1669390400
transform 1 0 63952 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_562
timestamp 1669390400
transform 1 0 64288 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_572
timestamp 1669390400
transform 1 0 65408 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_576
timestamp 1669390400
transform 1 0 65856 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_584
timestamp 1669390400
transform 1 0 66752 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_594
timestamp 1669390400
transform 1 0 67872 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_597
timestamp 1669390400
transform 1 0 68208 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_600
timestamp 1669390400
transform 1 0 68544 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_618
timestamp 1669390400
transform 1 0 70560 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_620
timestamp 1669390400
transform 1 0 70784 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_627
timestamp 1669390400
transform 1 0 71568 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_629
timestamp 1669390400
transform 1 0 71792 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_632
timestamp 1669390400
transform 1 0 72128 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_635
timestamp 1669390400
transform 1 0 72464 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_639
timestamp 1669390400
transform 1 0 72912 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_646
timestamp 1669390400
transform 1 0 73696 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_664
timestamp 1669390400
transform 1 0 75712 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_667
timestamp 1669390400
transform 1 0 76048 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_676
timestamp 1669390400
transform 1 0 77056 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_680
timestamp 1669390400
transform 1 0 77504 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_684
timestamp 1669390400
transform 1 0 77952 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_2
timestamp 1669390400
transform 1 0 1568 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_17
timestamp 1669390400
transform 1 0 3248 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_25
timestamp 1669390400
transform 1 0 4144 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_29 Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 4592 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_61
timestamp 1669390400
transform 1 0 8176 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_63
timestamp 1669390400
transform 1 0 8400 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_66
timestamp 1669390400
transform 1 0 8736 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_70
timestamp 1669390400
transform 1 0 9184 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_73
timestamp 1669390400
transform 1 0 9520 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_79
timestamp 1669390400
transform 1 0 10192 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_94
timestamp 1669390400
transform 1 0 11872 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_104
timestamp 1669390400
transform 1 0 12992 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_108
timestamp 1669390400
transform 1 0 13440 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_112
timestamp 1669390400
transform 1 0 13888 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_137
timestamp 1669390400
transform 1 0 16688 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_141
timestamp 1669390400
transform 1 0 17136 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_144
timestamp 1669390400
transform 1 0 17472 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_154
timestamp 1669390400
transform 1 0 18592 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_156
timestamp 1669390400
transform 1 0 18816 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_159
timestamp 1669390400
transform 1 0 19152 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_174
timestamp 1669390400
transform 1 0 20832 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_181
timestamp 1669390400
transform 1 0 21616 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_188
timestamp 1669390400
transform 1 0 22400 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_194
timestamp 1669390400
transform 1 0 23072 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_198
timestamp 1669390400
transform 1 0 23520 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_205
timestamp 1669390400
transform 1 0 24304 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_212
timestamp 1669390400
transform 1 0 25088 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_215
timestamp 1669390400
transform 1 0 25424 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_226
timestamp 1669390400
transform 1 0 26656 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_237
timestamp 1669390400
transform 1 0 27888 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_239
timestamp 1669390400
transform 1 0 28112 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_264
timestamp 1669390400
transform 1 0 30912 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_266
timestamp 1669390400
transform 1 0 31136 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_269
timestamp 1669390400
transform 1 0 31472 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_283
timestamp 1669390400
transform 1 0 33040 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_286
timestamp 1669390400
transform 1 0 33376 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_300
timestamp 1669390400
transform 1 0 34944 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_302
timestamp 1669390400
transform 1 0 35168 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_308
timestamp 1669390400
transform 1 0 35840 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_322
timestamp 1669390400
transform 1 0 37408 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_329
timestamp 1669390400
transform 1 0 38192 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_344
timestamp 1669390400
transform 1 0 39872 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_351
timestamp 1669390400
transform 1 0 40656 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_357
timestamp 1669390400
transform 1 0 41328 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_367
timestamp 1669390400
transform 1 0 42448 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_371
timestamp 1669390400
transform 1 0 42896 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_373
timestamp 1669390400
transform 1 0 43120 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_408
timestamp 1669390400
transform 1 0 47040 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_415
timestamp 1669390400
transform 1 0 47824 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_419
timestamp 1669390400
transform 1 0 48272 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_425
timestamp 1669390400
transform 1 0 48944 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_428
timestamp 1669390400
transform 1 0 49280 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_430
timestamp 1669390400
transform 1 0 49504 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_437
timestamp 1669390400
transform 1 0 50288 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_444
timestamp 1669390400
transform 1 0 51072 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_451
timestamp 1669390400
transform 1 0 51856 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_463
timestamp 1669390400
transform 1 0 53200 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_465
timestamp 1669390400
transform 1 0 53424 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_474
timestamp 1669390400
transform 1 0 54432 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_482
timestamp 1669390400
transform 1 0 55328 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_486
timestamp 1669390400
transform 1 0 55776 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_494
timestamp 1669390400
transform 1 0 56672 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_496
timestamp 1669390400
transform 1 0 56896 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_499
timestamp 1669390400
transform 1 0 57232 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_501
timestamp 1669390400
transform 1 0 57456 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_511
timestamp 1669390400
transform 1 0 58576 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_518
timestamp 1669390400
transform 1 0 59360 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_525
timestamp 1669390400
transform 1 0 60144 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_529
timestamp 1669390400
transform 1 0 60592 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_543
timestamp 1669390400
transform 1 0 62160 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_561
timestamp 1669390400
transform 1 0 64176 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_565
timestamp 1669390400
transform 1 0 64624 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_567
timestamp 1669390400
transform 1 0 64848 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_570
timestamp 1669390400
transform 1 0 65184 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_595
timestamp 1669390400
transform 1 0 67984 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_599
timestamp 1669390400
transform 1 0 68432 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_627
timestamp 1669390400
transform 1 0 71568 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_634
timestamp 1669390400
transform 1 0 72352 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_638
timestamp 1669390400
transform 1 0 72800 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_641
timestamp 1669390400
transform 1 0 73136 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_644
timestamp 1669390400
transform 1 0 73472 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_654
timestamp 1669390400
transform 1 0 74592 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_670
timestamp 1669390400
transform 1 0 76384 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_678
timestamp 1669390400
transform 1 0 77280 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_686
timestamp 1669390400
transform 1 0 78176 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_2
timestamp 1669390400
transform 1 0 1568 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_17
timestamp 1669390400
transform 1 0 3248 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_25
timestamp 1669390400
transform 1 0 4144 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_29
timestamp 1669390400
transform 1 0 4592 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_33
timestamp 1669390400
transform 1 0 5040 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_37 Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 5488 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_53
timestamp 1669390400
transform 1 0 7280 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_57
timestamp 1669390400
transform 1 0 7728 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_61
timestamp 1669390400
transform 1 0 8176 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_68
timestamp 1669390400
transform 1 0 8960 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_72
timestamp 1669390400
transform 1 0 9408 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_74
timestamp 1669390400
transform 1 0 9632 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_77
timestamp 1669390400
transform 1 0 9968 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_91
timestamp 1669390400
transform 1 0 11536 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_98
timestamp 1669390400
transform 1 0 12320 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_102
timestamp 1669390400
transform 1 0 12768 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_105
timestamp 1669390400
transform 1 0 13104 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_108
timestamp 1669390400
transform 1 0 13440 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_117
timestamp 1669390400
transform 1 0 14448 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_119
timestamp 1669390400
transform 1 0 14672 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_128
timestamp 1669390400
transform 1 0 15680 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_132
timestamp 1669390400
transform 1 0 16128 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_138
timestamp 1669390400
transform 1 0 16800 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_142
timestamp 1669390400
transform 1 0 17248 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_146
timestamp 1669390400
transform 1 0 17696 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_150
timestamp 1669390400
transform 1 0 18144 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_157
timestamp 1669390400
transform 1 0 18928 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_161
timestamp 1669390400
transform 1 0 19376 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_163
timestamp 1669390400
transform 1 0 19600 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_172
timestamp 1669390400
transform 1 0 20608 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_176
timestamp 1669390400
transform 1 0 21056 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_179
timestamp 1669390400
transform 1 0 21392 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_193
timestamp 1669390400
transform 1 0 22960 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_197
timestamp 1669390400
transform 1 0 23408 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_222
timestamp 1669390400
transform 1 0 26208 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_226
timestamp 1669390400
transform 1 0 26656 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_228
timestamp 1669390400
transform 1 0 26880 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_231
timestamp 1669390400
transform 1 0 27216 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_235
timestamp 1669390400
transform 1 0 27664 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_239
timestamp 1669390400
transform 1 0 28112 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_243
timestamp 1669390400
transform 1 0 28560 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_247
timestamp 1669390400
transform 1 0 29008 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_250
timestamp 1669390400
transform 1 0 29344 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_257
timestamp 1669390400
transform 1 0 30128 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_259
timestamp 1669390400
transform 1 0 30352 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_265
timestamp 1669390400
transform 1 0 31024 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_269
timestamp 1669390400
transform 1 0 31472 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_271
timestamp 1669390400
transform 1 0 31696 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_274
timestamp 1669390400
transform 1 0 32032 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_278
timestamp 1669390400
transform 1 0 32480 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_288
timestamp 1669390400
transform 1 0 33600 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_290
timestamp 1669390400
transform 1 0 33824 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_293
timestamp 1669390400
transform 1 0 34160 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_318
timestamp 1669390400
transform 1 0 36960 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_321
timestamp 1669390400
transform 1 0 37296 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_323
timestamp 1669390400
transform 1 0 37520 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_326
timestamp 1669390400
transform 1 0 37856 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_330
timestamp 1669390400
transform 1 0 38304 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_340
timestamp 1669390400
transform 1 0 39424 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_352
timestamp 1669390400
transform 1 0 40768 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_356
timestamp 1669390400
transform 1 0 41216 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_360
timestamp 1669390400
transform 1 0 41664 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_364
timestamp 1669390400
transform 1 0 42112 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_366
timestamp 1669390400
transform 1 0 42336 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_369
timestamp 1669390400
transform 1 0 42672 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_373
timestamp 1669390400
transform 1 0 43120 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_377
timestamp 1669390400
transform 1 0 43568 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_379
timestamp 1669390400
transform 1 0 43792 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_389
timestamp 1669390400
transform 1 0 44912 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_392
timestamp 1669390400
transform 1 0 45248 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_398
timestamp 1669390400
transform 1 0 45920 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_405
timestamp 1669390400
transform 1 0 46704 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_409
timestamp 1669390400
transform 1 0 47152 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_434
timestamp 1669390400
transform 1 0 49952 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_460
timestamp 1669390400
transform 1 0 52864 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_463
timestamp 1669390400
transform 1 0 53200 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_469
timestamp 1669390400
transform 1 0 53872 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_473
timestamp 1669390400
transform 1 0 54320 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_479
timestamp 1669390400
transform 1 0 54992 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_489
timestamp 1669390400
transform 1 0 56112 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_496
timestamp 1669390400
transform 1 0 56896 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_500
timestamp 1669390400
transform 1 0 57344 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_504
timestamp 1669390400
transform 1 0 57792 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_508
timestamp 1669390400
transform 1 0 58240 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_515
timestamp 1669390400
transform 1 0 59024 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_519
timestamp 1669390400
transform 1 0 59472 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_523
timestamp 1669390400
transform 1 0 59920 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_525
timestamp 1669390400
transform 1 0 60144 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_531
timestamp 1669390400
transform 1 0 60816 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_534
timestamp 1669390400
transform 1 0 61152 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_537
timestamp 1669390400
transform 1 0 61488 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_539
timestamp 1669390400
transform 1 0 61712 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_548
timestamp 1669390400
transform 1 0 62720 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_555
timestamp 1669390400
transform 1 0 63504 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_565
timestamp 1669390400
transform 1 0 64624 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_569
timestamp 1669390400
transform 1 0 65072 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_576
timestamp 1669390400
transform 1 0 65856 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_583
timestamp 1669390400
transform 1 0 66640 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_587
timestamp 1669390400
transform 1 0 67088 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_601
timestamp 1669390400
transform 1 0 68656 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_605
timestamp 1669390400
transform 1 0 69104 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_608
timestamp 1669390400
transform 1 0 69440 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_612
timestamp 1669390400
transform 1 0 69888 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_616
timestamp 1669390400
transform 1 0 70336 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_620
timestamp 1669390400
transform 1 0 70784 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_624
timestamp 1669390400
transform 1 0 71232 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_638
timestamp 1669390400
transform 1 0 72800 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_642
timestamp 1669390400
transform 1 0 73248 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_646
timestamp 1669390400
transform 1 0 73696 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_650
timestamp 1669390400
transform 1 0 74144 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_654
timestamp 1669390400
transform 1 0 74592 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_658
timestamp 1669390400
transform 1 0 75040 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_672
timestamp 1669390400
transform 1 0 76608 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_676
timestamp 1669390400
transform 1 0 77056 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_679
timestamp 1669390400
transform 1 0 77392 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_683
timestamp 1669390400
transform 1 0 77840 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_687
timestamp 1669390400
transform 1 0 78288 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_2
timestamp 1669390400
transform 1 0 1568 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_6
timestamp 1669390400
transform 1 0 2016 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_8
timestamp 1669390400
transform 1 0 2240 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_11
timestamp 1669390400
transform 1 0 2576 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_26
timestamp 1669390400
transform 1 0 4256 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_52
timestamp 1669390400
transform 1 0 7168 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_56
timestamp 1669390400
transform 1 0 7616 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_60
timestamp 1669390400
transform 1 0 8064 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_70
timestamp 1669390400
transform 1 0 9184 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_73
timestamp 1669390400
transform 1 0 9520 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_84
timestamp 1669390400
transform 1 0 10752 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_88
timestamp 1669390400
transform 1 0 11200 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_92
timestamp 1669390400
transform 1 0 11648 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_96
timestamp 1669390400
transform 1 0 12096 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_121
timestamp 1669390400
transform 1 0 14896 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_127
timestamp 1669390400
transform 1 0 15568 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_134
timestamp 1669390400
transform 1 0 16352 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_140
timestamp 1669390400
transform 1 0 17024 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_144
timestamp 1669390400
transform 1 0 17472 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_147
timestamp 1669390400
transform 1 0 17808 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_156
timestamp 1669390400
transform 1 0 18816 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_160
timestamp 1669390400
transform 1 0 19264 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_164
timestamp 1669390400
transform 1 0 19712 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_168 Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 20160 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_176
timestamp 1669390400
transform 1 0 21056 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_188
timestamp 1669390400
transform 1 0 22400 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_190
timestamp 1669390400
transform 1 0 22624 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_201
timestamp 1669390400
transform 1 0 23856 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_205
timestamp 1669390400
transform 1 0 24304 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_208
timestamp 1669390400
transform 1 0 24640 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_212
timestamp 1669390400
transform 1 0 25088 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_215
timestamp 1669390400
transform 1 0 25424 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_219
timestamp 1669390400
transform 1 0 25872 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_223
timestamp 1669390400
transform 1 0 26320 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_249
timestamp 1669390400
transform 1 0 29232 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_253
timestamp 1669390400
transform 1 0 29680 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_262
timestamp 1669390400
transform 1 0 30688 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_266
timestamp 1669390400
transform 1 0 31136 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_282
timestamp 1669390400
transform 1 0 32928 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_286
timestamp 1669390400
transform 1 0 33376 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_292
timestamp 1669390400
transform 1 0 34048 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_296
timestamp 1669390400
transform 1 0 34496 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_306
timestamp 1669390400
transform 1 0 35616 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_315
timestamp 1669390400
transform 1 0 36624 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_319
timestamp 1669390400
transform 1 0 37072 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_323
timestamp 1669390400
transform 1 0 37520 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_327
timestamp 1669390400
transform 1 0 37968 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_331
timestamp 1669390400
transform 1 0 38416 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_334
timestamp 1669390400
transform 1 0 38752 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_348
timestamp 1669390400
transform 1 0 40320 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_354
timestamp 1669390400
transform 1 0 40992 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_357
timestamp 1669390400
transform 1 0 41328 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_366
timestamp 1669390400
transform 1 0 42336 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_370
timestamp 1669390400
transform 1 0 42784 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_374
timestamp 1669390400
transform 1 0 43232 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_378
timestamp 1669390400
transform 1 0 43680 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_393
timestamp 1669390400
transform 1 0 45360 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_404
timestamp 1669390400
transform 1 0 46592 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_408
timestamp 1669390400
transform 1 0 47040 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_412
timestamp 1669390400
transform 1 0 47488 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_414
timestamp 1669390400
transform 1 0 47712 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_425
timestamp 1669390400
transform 1 0 48944 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_428
timestamp 1669390400
transform 1 0 49280 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_434
timestamp 1669390400
transform 1 0 49952 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_438
timestamp 1669390400
transform 1 0 50400 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_442
timestamp 1669390400
transform 1 0 50848 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_444
timestamp 1669390400
transform 1 0 51072 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_450
timestamp 1669390400
transform 1 0 51744 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_454
timestamp 1669390400
transform 1 0 52192 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_458
timestamp 1669390400
transform 1 0 52640 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_462
timestamp 1669390400
transform 1 0 53088 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_466
timestamp 1669390400
transform 1 0 53536 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_470
timestamp 1669390400
transform 1 0 53984 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_472
timestamp 1669390400
transform 1 0 54208 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_481
timestamp 1669390400
transform 1 0 55216 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_492
timestamp 1669390400
transform 1 0 56448 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_496
timestamp 1669390400
transform 1 0 56896 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_499
timestamp 1669390400
transform 1 0 57232 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_501
timestamp 1669390400
transform 1 0 57456 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_507
timestamp 1669390400
transform 1 0 58128 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_519
timestamp 1669390400
transform 1 0 59472 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_545
timestamp 1669390400
transform 1 0 62384 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_552
timestamp 1669390400
transform 1 0 63168 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_559
timestamp 1669390400
transform 1 0 63952 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_563
timestamp 1669390400
transform 1 0 64400 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_567
timestamp 1669390400
transform 1 0 64848 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_570
timestamp 1669390400
transform 1 0 65184 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_579
timestamp 1669390400
transform 1 0 66192 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_586
timestamp 1669390400
transform 1 0 66976 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_598
timestamp 1669390400
transform 1 0 68320 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_605
timestamp 1669390400
transform 1 0 69104 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_609
timestamp 1669390400
transform 1 0 69552 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_613
timestamp 1669390400
transform 1 0 70000 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_617
timestamp 1669390400
transform 1 0 70448 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_621
timestamp 1669390400
transform 1 0 70896 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_625
timestamp 1669390400
transform 1 0 71344 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_638
timestamp 1669390400
transform 1 0 72800 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_641
timestamp 1669390400
transform 1 0 73136 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_644
timestamp 1669390400
transform 1 0 73472 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_648
timestamp 1669390400
transform 1 0 73920 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_654
timestamp 1669390400
transform 1 0 74592 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_668
timestamp 1669390400
transform 1 0 76160 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_682
timestamp 1669390400
transform 1 0 77728 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_686
timestamp 1669390400
transform 1 0 78176 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_2
timestamp 1669390400
transform 1 0 1568 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_17
timestamp 1669390400
transform 1 0 3248 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_23
timestamp 1669390400
transform 1 0 3920 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_25
timestamp 1669390400
transform 1 0 4144 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_31
timestamp 1669390400
transform 1 0 4816 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_37
timestamp 1669390400
transform 1 0 5488 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_40
timestamp 1669390400
transform 1 0 5824 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_44
timestamp 1669390400
transform 1 0 6272 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_60
timestamp 1669390400
transform 1 0 8064 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_62
timestamp 1669390400
transform 1 0 8288 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_65
timestamp 1669390400
transform 1 0 8624 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_69
timestamp 1669390400
transform 1 0 9072 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_76
timestamp 1669390400
transform 1 0 9856 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_83
timestamp 1669390400
transform 1 0 10640 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_87
timestamp 1669390400
transform 1 0 11088 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_91
timestamp 1669390400
transform 1 0 11536 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_97
timestamp 1669390400
transform 1 0 12208 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_104
timestamp 1669390400
transform 1 0 12992 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_108
timestamp 1669390400
transform 1 0 13440 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_119
timestamp 1669390400
transform 1 0 14672 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_129
timestamp 1669390400
transform 1 0 15792 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_138
timestamp 1669390400
transform 1 0 16800 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_164
timestamp 1669390400
transform 1 0 19712 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_168
timestamp 1669390400
transform 1 0 20160 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_176
timestamp 1669390400
transform 1 0 21056 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_179
timestamp 1669390400
transform 1 0 21392 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_192
timestamp 1669390400
transform 1 0 22848 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_196
timestamp 1669390400
transform 1 0 23296 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_207
timestamp 1669390400
transform 1 0 24528 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_209
timestamp 1669390400
transform 1 0 24752 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_215
timestamp 1669390400
transform 1 0 25424 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_217
timestamp 1669390400
transform 1 0 25648 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_220
timestamp 1669390400
transform 1 0 25984 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_224
timestamp 1669390400
transform 1 0 26432 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_231
timestamp 1669390400
transform 1 0 27216 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_243
timestamp 1669390400
transform 1 0 28560 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_247
timestamp 1669390400
transform 1 0 29008 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_250
timestamp 1669390400
transform 1 0 29344 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_253
timestamp 1669390400
transform 1 0 29680 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_255
timestamp 1669390400
transform 1 0 29904 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_258
timestamp 1669390400
transform 1 0 30240 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_262
timestamp 1669390400
transform 1 0 30688 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_268
timestamp 1669390400
transform 1 0 31360 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_283
timestamp 1669390400
transform 1 0 33040 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_291
timestamp 1669390400
transform 1 0 33936 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_295
timestamp 1669390400
transform 1 0 34384 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_307
timestamp 1669390400
transform 1 0 35728 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_314
timestamp 1669390400
transform 1 0 36512 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_318
timestamp 1669390400
transform 1 0 36960 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_321
timestamp 1669390400
transform 1 0 37296 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_324
timestamp 1669390400
transform 1 0 37632 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_328
timestamp 1669390400
transform 1 0 38080 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_336
timestamp 1669390400
transform 1 0 38976 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_338
timestamp 1669390400
transform 1 0 39200 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_352
timestamp 1669390400
transform 1 0 40768 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_359
timestamp 1669390400
transform 1 0 41552 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_365
timestamp 1669390400
transform 1 0 42224 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_379
timestamp 1669390400
transform 1 0 43792 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_385
timestamp 1669390400
transform 1 0 44464 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_389
timestamp 1669390400
transform 1 0 44912 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_392
timestamp 1669390400
transform 1 0 45248 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_395
timestamp 1669390400
transform 1 0 45584 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_405
timestamp 1669390400
transform 1 0 46704 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_409
timestamp 1669390400
transform 1 0 47152 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_413
timestamp 1669390400
transform 1 0 47600 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_417
timestamp 1669390400
transform 1 0 48048 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_421
timestamp 1669390400
transform 1 0 48496 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_425
timestamp 1669390400
transform 1 0 48944 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_431
timestamp 1669390400
transform 1 0 49616 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_438
timestamp 1669390400
transform 1 0 50400 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_440
timestamp 1669390400
transform 1 0 50624 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_451
timestamp 1669390400
transform 1 0 51856 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_455
timestamp 1669390400
transform 1 0 52304 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_459
timestamp 1669390400
transform 1 0 52752 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_463
timestamp 1669390400
transform 1 0 53200 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_466
timestamp 1669390400
transform 1 0 53536 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_470
timestamp 1669390400
transform 1 0 53984 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_479
timestamp 1669390400
transform 1 0 54992 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_491
timestamp 1669390400
transform 1 0 56336 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_498
timestamp 1669390400
transform 1 0 57120 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_502
timestamp 1669390400
transform 1 0 57568 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_506
timestamp 1669390400
transform 1 0 58016 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_510
timestamp 1669390400
transform 1 0 58464 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_514
timestamp 1669390400
transform 1 0 58912 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_523
timestamp 1669390400
transform 1 0 59920 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_527
timestamp 1669390400
transform 1 0 60368 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_531
timestamp 1669390400
transform 1 0 60816 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_534
timestamp 1669390400
transform 1 0 61152 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_537
timestamp 1669390400
transform 1 0 61488 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_552
timestamp 1669390400
transform 1 0 63168 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_556
timestamp 1669390400
transform 1 0 63616 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_560
timestamp 1669390400
transform 1 0 64064 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_567
timestamp 1669390400
transform 1 0 64848 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_584
timestamp 1669390400
transform 1 0 66752 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_588
timestamp 1669390400
transform 1 0 67200 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_600
timestamp 1669390400
transform 1 0 68544 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_602
timestamp 1669390400
transform 1 0 68768 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_605
timestamp 1669390400
transform 1 0 69104 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_629
timestamp 1669390400
transform 1 0 71792 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_639
timestamp 1669390400
transform 1 0 72912 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_643
timestamp 1669390400
transform 1 0 73360 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_647
timestamp 1669390400
transform 1 0 73808 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_651
timestamp 1669390400
transform 1 0 74256 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_655
timestamp 1669390400
transform 1 0 74704 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_670
timestamp 1669390400
transform 1 0 76384 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_676
timestamp 1669390400
transform 1 0 77056 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_685
timestamp 1669390400
transform 1 0 78064 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_687
timestamp 1669390400
transform 1 0 78288 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_2
timestamp 1669390400
transform 1 0 1568 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_5
timestamp 1669390400
transform 1 0 1904 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_9
timestamp 1669390400
transform 1 0 2352 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_17
timestamp 1669390400
transform 1 0 3248 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_31
timestamp 1669390400
transform 1 0 4816 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_41
timestamp 1669390400
transform 1 0 5936 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_47
timestamp 1669390400
transform 1 0 6608 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_55
timestamp 1669390400
transform 1 0 7504 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_70
timestamp 1669390400
transform 1 0 9184 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_73
timestamp 1669390400
transform 1 0 9520 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_79
timestamp 1669390400
transform 1 0 10192 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_83
timestamp 1669390400
transform 1 0 10640 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_87
timestamp 1669390400
transform 1 0 11088 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_95
timestamp 1669390400
transform 1 0 11984 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_99
timestamp 1669390400
transform 1 0 12432 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_101
timestamp 1669390400
transform 1 0 12656 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_104
timestamp 1669390400
transform 1 0 12992 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_116
timestamp 1669390400
transform 1 0 14336 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_123
timestamp 1669390400
transform 1 0 15120 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_127
timestamp 1669390400
transform 1 0 15568 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_131
timestamp 1669390400
transform 1 0 16016 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_135
timestamp 1669390400
transform 1 0 16464 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_139
timestamp 1669390400
transform 1 0 16912 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_141
timestamp 1669390400
transform 1 0 17136 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_144
timestamp 1669390400
transform 1 0 17472 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_147
timestamp 1669390400
transform 1 0 17808 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_161
timestamp 1669390400
transform 1 0 19376 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_177
timestamp 1669390400
transform 1 0 21168 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_181
timestamp 1669390400
transform 1 0 21616 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_183
timestamp 1669390400
transform 1 0 21840 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_197
timestamp 1669390400
transform 1 0 23408 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_204
timestamp 1669390400
transform 1 0 24192 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_208
timestamp 1669390400
transform 1 0 24640 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_211
timestamp 1669390400
transform 1 0 24976 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_215
timestamp 1669390400
transform 1 0 25424 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_218
timestamp 1669390400
transform 1 0 25760 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_222
timestamp 1669390400
transform 1 0 26208 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_228
timestamp 1669390400
transform 1 0 26880 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_232
timestamp 1669390400
transform 1 0 27328 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_242
timestamp 1669390400
transform 1 0 28448 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_249
timestamp 1669390400
transform 1 0 29232 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_253
timestamp 1669390400
transform 1 0 29680 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_257
timestamp 1669390400
transform 1 0 30128 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_261
timestamp 1669390400
transform 1 0 30576 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_263
timestamp 1669390400
transform 1 0 30800 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_266
timestamp 1669390400
transform 1 0 31136 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_273
timestamp 1669390400
transform 1 0 31920 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_283
timestamp 1669390400
transform 1 0 33040 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_286
timestamp 1669390400
transform 1 0 33376 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_302
timestamp 1669390400
transform 1 0 35168 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_333
timestamp 1669390400
transform 1 0 38640 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_337
timestamp 1669390400
transform 1 0 39088 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_341
timestamp 1669390400
transform 1 0 39536 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_351
timestamp 1669390400
transform 1 0 40656 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_357
timestamp 1669390400
transform 1 0 41328 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_373
timestamp 1669390400
transform 1 0 43120 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_381
timestamp 1669390400
transform 1 0 44016 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_390
timestamp 1669390400
transform 1 0 45024 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_394
timestamp 1669390400
transform 1 0 45472 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_415
timestamp 1669390400
transform 1 0 47824 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_422
timestamp 1669390400
transform 1 0 48608 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_428
timestamp 1669390400
transform 1 0 49280 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_453
timestamp 1669390400
transform 1 0 52080 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_464
timestamp 1669390400
transform 1 0 53312 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_468
timestamp 1669390400
transform 1 0 53760 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_496
timestamp 1669390400
transform 1 0 56896 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_499
timestamp 1669390400
transform 1 0 57232 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_502
timestamp 1669390400
transform 1 0 57568 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_506
timestamp 1669390400
transform 1 0 58016 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_510
timestamp 1669390400
transform 1 0 58464 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_514
timestamp 1669390400
transform 1 0 58912 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_518
timestamp 1669390400
transform 1 0 59360 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_522
timestamp 1669390400
transform 1 0 59808 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_526
timestamp 1669390400
transform 1 0 60256 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_530
timestamp 1669390400
transform 1 0 60704 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_534
timestamp 1669390400
transform 1 0 61152 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_538
timestamp 1669390400
transform 1 0 61600 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_542
timestamp 1669390400
transform 1 0 62048 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_546
timestamp 1669390400
transform 1 0 62496 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_555
timestamp 1669390400
transform 1 0 63504 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_559
timestamp 1669390400
transform 1 0 63952 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_563
timestamp 1669390400
transform 1 0 64400 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_567
timestamp 1669390400
transform 1 0 64848 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_570
timestamp 1669390400
transform 1 0 65184 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_576
timestamp 1669390400
transform 1 0 65856 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_580
timestamp 1669390400
transform 1 0 66304 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_584
timestamp 1669390400
transform 1 0 66752 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_593
timestamp 1669390400
transform 1 0 67760 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_597
timestamp 1669390400
transform 1 0 68208 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_601
timestamp 1669390400
transform 1 0 68656 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_605
timestamp 1669390400
transform 1 0 69104 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_616
timestamp 1669390400
transform 1 0 70336 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_620
timestamp 1669390400
transform 1 0 70784 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_624
timestamp 1669390400
transform 1 0 71232 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_638
timestamp 1669390400
transform 1 0 72800 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_641
timestamp 1669390400
transform 1 0 73136 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_644
timestamp 1669390400
transform 1 0 73472 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_648
timestamp 1669390400
transform 1 0 73920 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_652
timestamp 1669390400
transform 1 0 74368 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_656
timestamp 1669390400
transform 1 0 74816 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_663
timestamp 1669390400
transform 1 0 75600 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_677
timestamp 1669390400
transform 1 0 77168 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_685
timestamp 1669390400
transform 1 0 78064 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_687
timestamp 1669390400
transform 1 0 78288 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_2
timestamp 1669390400
transform 1 0 1568 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_8
timestamp 1669390400
transform 1 0 2240 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_12
timestamp 1669390400
transform 1 0 2688 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_19
timestamp 1669390400
transform 1 0 3472 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_33
timestamp 1669390400
transform 1 0 5040 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_37
timestamp 1669390400
transform 1 0 5488 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_41
timestamp 1669390400
transform 1 0 5936 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_45
timestamp 1669390400
transform 1 0 6384 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_49
timestamp 1669390400
transform 1 0 6832 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_53
timestamp 1669390400
transform 1 0 7280 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_63
timestamp 1669390400
transform 1 0 8400 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_73
timestamp 1669390400
transform 1 0 9520 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_80
timestamp 1669390400
transform 1 0 10304 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_84
timestamp 1669390400
transform 1 0 10752 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_88
timestamp 1669390400
transform 1 0 11200 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_104
timestamp 1669390400
transform 1 0 12992 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_108
timestamp 1669390400
transform 1 0 13440 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_132
timestamp 1669390400
transform 1 0 16128 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_138
timestamp 1669390400
transform 1 0 16800 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_145
timestamp 1669390400
transform 1 0 17584 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_160
timestamp 1669390400
transform 1 0 19264 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_170
timestamp 1669390400
transform 1 0 20384 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_174
timestamp 1669390400
transform 1 0 20832 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_176
timestamp 1669390400
transform 1 0 21056 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_179
timestamp 1669390400
transform 1 0 21392 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_182
timestamp 1669390400
transform 1 0 21728 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_192
timestamp 1669390400
transform 1 0 22848 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_206
timestamp 1669390400
transform 1 0 24416 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_210
timestamp 1669390400
transform 1 0 24864 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_214
timestamp 1669390400
transform 1 0 25312 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_222
timestamp 1669390400
transform 1 0 26208 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_225
timestamp 1669390400
transform 1 0 26544 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_232
timestamp 1669390400
transform 1 0 27328 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_247
timestamp 1669390400
transform 1 0 29008 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_250
timestamp 1669390400
transform 1 0 29344 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_253
timestamp 1669390400
transform 1 0 29680 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_255
timestamp 1669390400
transform 1 0 29904 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_264
timestamp 1669390400
transform 1 0 30912 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_278
timestamp 1669390400
transform 1 0 32480 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_282
timestamp 1669390400
transform 1 0 32928 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_285
timestamp 1669390400
transform 1 0 33264 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_293
timestamp 1669390400
transform 1 0 34160 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_297
timestamp 1669390400
transform 1 0 34608 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_300
timestamp 1669390400
transform 1 0 34944 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_304
timestamp 1669390400
transform 1 0 35392 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_308
timestamp 1669390400
transform 1 0 35840 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_318
timestamp 1669390400
transform 1 0 36960 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_321
timestamp 1669390400
transform 1 0 37296 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_332
timestamp 1669390400
transform 1 0 38528 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_348
timestamp 1669390400
transform 1 0 40320 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_350
timestamp 1669390400
transform 1 0 40544 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_353
timestamp 1669390400
transform 1 0 40880 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_378
timestamp 1669390400
transform 1 0 43680 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_386
timestamp 1669390400
transform 1 0 44576 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_392
timestamp 1669390400
transform 1 0 45248 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_408
timestamp 1669390400
transform 1 0 47040 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_418
timestamp 1669390400
transform 1 0 48160 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_425
timestamp 1669390400
transform 1 0 48944 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_429
timestamp 1669390400
transform 1 0 49392 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_433
timestamp 1669390400
transform 1 0 49840 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_435
timestamp 1669390400
transform 1 0 50064 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_446
timestamp 1669390400
transform 1 0 51296 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_453
timestamp 1669390400
transform 1 0 52080 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_457
timestamp 1669390400
transform 1 0 52528 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_463
timestamp 1669390400
transform 1 0 53200 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_466
timestamp 1669390400
transform 1 0 53536 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_470
timestamp 1669390400
transform 1 0 53984 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_474
timestamp 1669390400
transform 1 0 54432 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_489
timestamp 1669390400
transform 1 0 56112 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_496
timestamp 1669390400
transform 1 0 56896 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_503
timestamp 1669390400
transform 1 0 57680 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_507
timestamp 1669390400
transform 1 0 58128 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_511
timestamp 1669390400
transform 1 0 58576 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_515
timestamp 1669390400
transform 1 0 59024 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_530
timestamp 1669390400
transform 1 0 60704 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_534
timestamp 1669390400
transform 1 0 61152 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_548
timestamp 1669390400
transform 1 0 62720 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_562
timestamp 1669390400
transform 1 0 64288 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_566
timestamp 1669390400
transform 1 0 64736 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_573
timestamp 1669390400
transform 1 0 65520 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_577
timestamp 1669390400
transform 1 0 65968 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_581
timestamp 1669390400
transform 1 0 66416 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_587
timestamp 1669390400
transform 1 0 67088 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_597
timestamp 1669390400
transform 1 0 68208 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_601
timestamp 1669390400
transform 1 0 68656 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_605
timestamp 1669390400
transform 1 0 69104 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_608
timestamp 1669390400
transform 1 0 69440 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_610
timestamp 1669390400
transform 1 0 69664 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_613
timestamp 1669390400
transform 1 0 70000 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_619
timestamp 1669390400
transform 1 0 70672 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_633
timestamp 1669390400
transform 1 0 72240 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_647
timestamp 1669390400
transform 1 0 73808 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_651
timestamp 1669390400
transform 1 0 74256 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_658
timestamp 1669390400
transform 1 0 75040 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_672
timestamp 1669390400
transform 1 0 76608 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_676
timestamp 1669390400
transform 1 0 77056 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_685
timestamp 1669390400
transform 1 0 78064 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_687
timestamp 1669390400
transform 1 0 78288 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_2
timestamp 1669390400
transform 1 0 1568 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_17
timestamp 1669390400
transform 1 0 3248 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_23
timestamp 1669390400
transform 1 0 3920 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_35
timestamp 1669390400
transform 1 0 5264 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_42
timestamp 1669390400
transform 1 0 6048 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_54
timestamp 1669390400
transform 1 0 7392 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_63
timestamp 1669390400
transform 1 0 8400 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_70
timestamp 1669390400
transform 1 0 9184 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_73
timestamp 1669390400
transform 1 0 9520 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_76
timestamp 1669390400
transform 1 0 9856 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_91
timestamp 1669390400
transform 1 0 11536 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_98
timestamp 1669390400
transform 1 0 12320 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_102
timestamp 1669390400
transform 1 0 12768 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_104
timestamp 1669390400
transform 1 0 12992 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_113
timestamp 1669390400
transform 1 0 14000 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_117
timestamp 1669390400
transform 1 0 14448 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_120
timestamp 1669390400
transform 1 0 14784 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_124
timestamp 1669390400
transform 1 0 15232 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_128
timestamp 1669390400
transform 1 0 15680 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_136
timestamp 1669390400
transform 1 0 16576 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_140
timestamp 1669390400
transform 1 0 17024 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_144
timestamp 1669390400
transform 1 0 17472 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_156
timestamp 1669390400
transform 1 0 18816 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_163
timestamp 1669390400
transform 1 0 19600 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_169
timestamp 1669390400
transform 1 0 20272 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_173
timestamp 1669390400
transform 1 0 20720 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_177
timestamp 1669390400
transform 1 0 21168 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_179
timestamp 1669390400
transform 1 0 21392 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_182
timestamp 1669390400
transform 1 0 21728 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_192
timestamp 1669390400
transform 1 0 22848 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_207
timestamp 1669390400
transform 1 0 24528 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_209
timestamp 1669390400
transform 1 0 24752 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_212
timestamp 1669390400
transform 1 0 25088 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_215
timestamp 1669390400
transform 1 0 25424 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_225
timestamp 1669390400
transform 1 0 26544 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_231
timestamp 1669390400
transform 1 0 27216 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_241
timestamp 1669390400
transform 1 0 28336 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_248
timestamp 1669390400
transform 1 0 29120 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_250
timestamp 1669390400
transform 1 0 29344 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_253
timestamp 1669390400
transform 1 0 29680 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_257
timestamp 1669390400
transform 1 0 30128 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_264
timestamp 1669390400
transform 1 0 30912 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_276
timestamp 1669390400
transform 1 0 32256 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_283
timestamp 1669390400
transform 1 0 33040 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_286
timestamp 1669390400
transform 1 0 33376 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_292
timestamp 1669390400
transform 1 0 34048 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_296
timestamp 1669390400
transform 1 0 34496 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_303
timestamp 1669390400
transform 1 0 35280 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_310
timestamp 1669390400
transform 1 0 36064 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_317
timestamp 1669390400
transform 1 0 36848 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_324
timestamp 1669390400
transform 1 0 37632 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_328
timestamp 1669390400
transform 1 0 38080 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_332
timestamp 1669390400
transform 1 0 38528 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_340
timestamp 1669390400
transform 1 0 39424 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_343
timestamp 1669390400
transform 1 0 39760 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_347
timestamp 1669390400
transform 1 0 40208 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_354
timestamp 1669390400
transform 1 0 40992 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_357
timestamp 1669390400
transform 1 0 41328 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_368
timestamp 1669390400
transform 1 0 42560 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_375
timestamp 1669390400
transform 1 0 43344 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_379
timestamp 1669390400
transform 1 0 43792 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_383
timestamp 1669390400
transform 1 0 44240 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_415
timestamp 1669390400
transform 1 0 47824 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_425
timestamp 1669390400
transform 1 0 48944 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_428
timestamp 1669390400
transform 1 0 49280 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_431
timestamp 1669390400
transform 1 0 49616 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_433
timestamp 1669390400
transform 1 0 49840 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_436
timestamp 1669390400
transform 1 0 50176 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_461
timestamp 1669390400
transform 1 0 52976 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_465
timestamp 1669390400
transform 1 0 53424 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_468
timestamp 1669390400
transform 1 0 53760 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_484
timestamp 1669390400
transform 1 0 55552 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_494
timestamp 1669390400
transform 1 0 56672 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_496
timestamp 1669390400
transform 1 0 56896 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_499
timestamp 1669390400
transform 1 0 57232 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_508
timestamp 1669390400
transform 1 0 58240 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_512
timestamp 1669390400
transform 1 0 58688 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_516
timestamp 1669390400
transform 1 0 59136 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_541
timestamp 1669390400
transform 1 0 61936 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_553
timestamp 1669390400
transform 1 0 63280 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_557
timestamp 1669390400
transform 1 0 63728 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_561
timestamp 1669390400
transform 1 0 64176 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_565
timestamp 1669390400
transform 1 0 64624 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_567
timestamp 1669390400
transform 1 0 64848 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_570
timestamp 1669390400
transform 1 0 65184 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_573
timestamp 1669390400
transform 1 0 65520 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_577
timestamp 1669390400
transform 1 0 65968 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_579
timestamp 1669390400
transform 1 0 66192 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_582
timestamp 1669390400
transform 1 0 66528 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_586
timestamp 1669390400
transform 1 0 66976 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_593
timestamp 1669390400
transform 1 0 67760 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_600
timestamp 1669390400
transform 1 0 68544 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_607
timestamp 1669390400
transform 1 0 69328 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_611
timestamp 1669390400
transform 1 0 69776 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_615
timestamp 1669390400
transform 1 0 70224 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_619
timestamp 1669390400
transform 1 0 70672 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_623
timestamp 1669390400
transform 1 0 71120 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_625
timestamp 1669390400
transform 1 0 71344 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_631
timestamp 1669390400
transform 1 0 72016 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_635
timestamp 1669390400
transform 1 0 72464 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_641
timestamp 1669390400
transform 1 0 73136 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_650
timestamp 1669390400
transform 1 0 74144 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_654
timestamp 1669390400
transform 1 0 74592 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_670
timestamp 1669390400
transform 1 0 76384 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_677
timestamp 1669390400
transform 1 0 77168 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_681
timestamp 1669390400
transform 1 0 77616 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_685
timestamp 1669390400
transform 1 0 78064 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_687
timestamp 1669390400
transform 1 0 78288 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_2
timestamp 1669390400
transform 1 0 1568 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_6
timestamp 1669390400
transform 1 0 2016 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_14
timestamp 1669390400
transform 1 0 2912 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_24
timestamp 1669390400
transform 1 0 4032 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_31
timestamp 1669390400
transform 1 0 4816 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_37
timestamp 1669390400
transform 1 0 5488 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_43
timestamp 1669390400
transform 1 0 6160 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_47
timestamp 1669390400
transform 1 0 6608 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_53
timestamp 1669390400
transform 1 0 7280 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_65
timestamp 1669390400
transform 1 0 8624 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_69
timestamp 1669390400
transform 1 0 9072 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_73
timestamp 1669390400
transform 1 0 9520 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_77
timestamp 1669390400
transform 1 0 9968 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_81
timestamp 1669390400
transform 1 0 10416 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_94
timestamp 1669390400
transform 1 0 11872 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_98
timestamp 1669390400
transform 1 0 12320 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_101
timestamp 1669390400
transform 1 0 12656 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_105
timestamp 1669390400
transform 1 0 13104 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_108
timestamp 1669390400
transform 1 0 13440 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_114
timestamp 1669390400
transform 1 0 14112 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_116
timestamp 1669390400
transform 1 0 14336 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_125
timestamp 1669390400
transform 1 0 15344 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_129
timestamp 1669390400
transform 1 0 15792 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_135
timestamp 1669390400
transform 1 0 16464 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_139
timestamp 1669390400
transform 1 0 16912 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_146
timestamp 1669390400
transform 1 0 17696 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_158
timestamp 1669390400
transform 1 0 19040 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_165
timestamp 1669390400
transform 1 0 19824 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_167
timestamp 1669390400
transform 1 0 20048 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_170
timestamp 1669390400
transform 1 0 20384 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_174
timestamp 1669390400
transform 1 0 20832 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_176
timestamp 1669390400
transform 1 0 21056 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_179
timestamp 1669390400
transform 1 0 21392 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_183
timestamp 1669390400
transform 1 0 21840 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_189
timestamp 1669390400
transform 1 0 22512 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_196
timestamp 1669390400
transform 1 0 23296 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_203
timestamp 1669390400
transform 1 0 24080 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_207
timestamp 1669390400
transform 1 0 24528 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_211
timestamp 1669390400
transform 1 0 24976 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_213
timestamp 1669390400
transform 1 0 25200 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_216
timestamp 1669390400
transform 1 0 25536 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_230
timestamp 1669390400
transform 1 0 27104 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_240
timestamp 1669390400
transform 1 0 28224 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_244
timestamp 1669390400
transform 1 0 28672 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_250
timestamp 1669390400
transform 1 0 29344 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_256
timestamp 1669390400
transform 1 0 30016 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_260
timestamp 1669390400
transform 1 0 30464 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_266
timestamp 1669390400
transform 1 0 31136 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_274
timestamp 1669390400
transform 1 0 32032 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_278
timestamp 1669390400
transform 1 0 32480 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_282
timestamp 1669390400
transform 1 0 32928 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_288
timestamp 1669390400
transform 1 0 33600 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_292
timestamp 1669390400
transform 1 0 34048 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_302
timestamp 1669390400
transform 1 0 35168 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_310
timestamp 1669390400
transform 1 0 36064 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_317
timestamp 1669390400
transform 1 0 36848 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_321
timestamp 1669390400
transform 1 0 37296 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_324
timestamp 1669390400
transform 1 0 37632 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_328
timestamp 1669390400
transform 1 0 38080 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_330
timestamp 1669390400
transform 1 0 38304 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_336
timestamp 1669390400
transform 1 0 38976 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_348
timestamp 1669390400
transform 1 0 40320 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_352
timestamp 1669390400
transform 1 0 40768 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_362
timestamp 1669390400
transform 1 0 41888 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_366
timestamp 1669390400
transform 1 0 42336 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_370
timestamp 1669390400
transform 1 0 42784 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_378
timestamp 1669390400
transform 1 0 43680 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_382
timestamp 1669390400
transform 1 0 44128 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_389
timestamp 1669390400
transform 1 0 44912 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_392
timestamp 1669390400
transform 1 0 45248 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_406
timestamp 1669390400
transform 1 0 46816 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_414
timestamp 1669390400
transform 1 0 47712 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_424
timestamp 1669390400
transform 1 0 48832 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_426
timestamp 1669390400
transform 1 0 49056 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_429
timestamp 1669390400
transform 1 0 49392 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_439
timestamp 1669390400
transform 1 0 50512 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_446
timestamp 1669390400
transform 1 0 51296 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_450
timestamp 1669390400
transform 1 0 51744 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_454
timestamp 1669390400
transform 1 0 52192 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_458
timestamp 1669390400
transform 1 0 52640 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_460
timestamp 1669390400
transform 1 0 52864 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_463
timestamp 1669390400
transform 1 0 53200 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_467
timestamp 1669390400
transform 1 0 53648 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_470
timestamp 1669390400
transform 1 0 53984 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_474
timestamp 1669390400
transform 1 0 54432 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_478
timestamp 1669390400
transform 1 0 54880 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_480
timestamp 1669390400
transform 1 0 55104 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_483
timestamp 1669390400
transform 1 0 55440 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_485
timestamp 1669390400
transform 1 0 55664 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_488
timestamp 1669390400
transform 1 0 56000 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_490
timestamp 1669390400
transform 1 0 56224 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_504
timestamp 1669390400
transform 1 0 57792 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_508
timestamp 1669390400
transform 1 0 58240 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_512
timestamp 1669390400
transform 1 0 58688 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_516
timestamp 1669390400
transform 1 0 59136 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_520
timestamp 1669390400
transform 1 0 59584 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_524
timestamp 1669390400
transform 1 0 60032 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_534
timestamp 1669390400
transform 1 0 61152 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_542
timestamp 1669390400
transform 1 0 62048 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_550
timestamp 1669390400
transform 1 0 62944 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_557
timestamp 1669390400
transform 1 0 63728 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_565
timestamp 1669390400
transform 1 0 64624 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_567
timestamp 1669390400
transform 1 0 64848 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_576
timestamp 1669390400
transform 1 0 65856 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_580
timestamp 1669390400
transform 1 0 66304 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_582
timestamp 1669390400
transform 1 0 66528 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_596
timestamp 1669390400
transform 1 0 68096 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_600
timestamp 1669390400
transform 1 0 68544 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_602
timestamp 1669390400
transform 1 0 68768 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_605
timestamp 1669390400
transform 1 0 69104 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_612
timestamp 1669390400
transform 1 0 69888 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_619
timestamp 1669390400
transform 1 0 70672 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_626
timestamp 1669390400
transform 1 0 71456 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_636
timestamp 1669390400
transform 1 0 72576 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_644
timestamp 1669390400
transform 1 0 73472 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_648
timestamp 1669390400
transform 1 0 73920 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_652
timestamp 1669390400
transform 1 0 74368 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_655
timestamp 1669390400
transform 1 0 74704 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_659
timestamp 1669390400
transform 1 0 75152 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_663
timestamp 1669390400
transform 1 0 75600 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_667
timestamp 1669390400
transform 1 0 76048 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_673
timestamp 1669390400
transform 1 0 76720 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_676
timestamp 1669390400
transform 1 0 77056 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_682
timestamp 1669390400
transform 1 0 77728 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_686
timestamp 1669390400
transform 1 0 78176 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_2
timestamp 1669390400
transform 1 0 1568 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_4
timestamp 1669390400
transform 1 0 1792 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_7
timestamp 1669390400
transform 1 0 2128 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_14
timestamp 1669390400
transform 1 0 2912 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_24
timestamp 1669390400
transform 1 0 4032 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_34
timestamp 1669390400
transform 1 0 5152 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_60
timestamp 1669390400
transform 1 0 8064 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_69
timestamp 1669390400
transform 1 0 9072 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_73
timestamp 1669390400
transform 1 0 9520 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_77
timestamp 1669390400
transform 1 0 9968 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_79
timestamp 1669390400
transform 1 0 10192 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_84
timestamp 1669390400
transform 1 0 10752 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_94
timestamp 1669390400
transform 1 0 11872 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_103
timestamp 1669390400
transform 1 0 12880 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_114
timestamp 1669390400
transform 1 0 14112 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_118
timestamp 1669390400
transform 1 0 14560 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_128
timestamp 1669390400
transform 1 0 15680 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_132
timestamp 1669390400
transform 1 0 16128 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_134
timestamp 1669390400
transform 1 0 16352 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_137
timestamp 1669390400
transform 1 0 16688 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_141
timestamp 1669390400
transform 1 0 17136 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_144
timestamp 1669390400
transform 1 0 17472 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_147
timestamp 1669390400
transform 1 0 17808 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_158
timestamp 1669390400
transform 1 0 19040 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_168
timestamp 1669390400
transform 1 0 20160 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_174
timestamp 1669390400
transform 1 0 20832 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_181
timestamp 1669390400
transform 1 0 21616 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_207
timestamp 1669390400
transform 1 0 24528 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_211
timestamp 1669390400
transform 1 0 24976 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_215
timestamp 1669390400
transform 1 0 25424 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_221
timestamp 1669390400
transform 1 0 26096 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_225
timestamp 1669390400
transform 1 0 26544 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_233
timestamp 1669390400
transform 1 0 27440 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_242
timestamp 1669390400
transform 1 0 28448 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_257
timestamp 1669390400
transform 1 0 30128 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_264
timestamp 1669390400
transform 1 0 30912 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_279
timestamp 1669390400
transform 1 0 32592 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_283
timestamp 1669390400
transform 1 0 33040 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_286
timestamp 1669390400
transform 1 0 33376 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_300
timestamp 1669390400
transform 1 0 34944 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_314
timestamp 1669390400
transform 1 0 36512 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_318
timestamp 1669390400
transform 1 0 36960 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_326
timestamp 1669390400
transform 1 0 37856 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_340
timestamp 1669390400
transform 1 0 39424 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_354
timestamp 1669390400
transform 1 0 40992 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_357
timestamp 1669390400
transform 1 0 41328 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_360
timestamp 1669390400
transform 1 0 41664 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_364
timestamp 1669390400
transform 1 0 42112 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_372
timestamp 1669390400
transform 1 0 43008 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_386
timestamp 1669390400
transform 1 0 44576 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_396
timestamp 1669390400
transform 1 0 45696 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_400
timestamp 1669390400
transform 1 0 46144 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_425
timestamp 1669390400
transform 1 0 48944 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_428
timestamp 1669390400
transform 1 0 49280 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_434
timestamp 1669390400
transform 1 0 49952 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_436
timestamp 1669390400
transform 1 0 50176 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_439
timestamp 1669390400
transform 1 0 50512 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_455
timestamp 1669390400
transform 1 0 52304 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_458
timestamp 1669390400
transform 1 0 52640 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_468
timestamp 1669390400
transform 1 0 53760 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_475
timestamp 1669390400
transform 1 0 54544 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_479
timestamp 1669390400
transform 1 0 54992 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_483
timestamp 1669390400
transform 1 0 55440 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_485
timestamp 1669390400
transform 1 0 55664 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_488
timestamp 1669390400
transform 1 0 56000 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_496
timestamp 1669390400
transform 1 0 56896 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_499
timestamp 1669390400
transform 1 0 57232 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_506
timestamp 1669390400
transform 1 0 58016 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_510
timestamp 1669390400
transform 1 0 58464 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_526
timestamp 1669390400
transform 1 0 60256 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_534
timestamp 1669390400
transform 1 0 61152 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_538
timestamp 1669390400
transform 1 0 61600 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_547
timestamp 1669390400
transform 1 0 62608 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_557
timestamp 1669390400
transform 1 0 63728 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_567
timestamp 1669390400
transform 1 0 64848 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_570
timestamp 1669390400
transform 1 0 65184 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_580
timestamp 1669390400
transform 1 0 66304 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_594
timestamp 1669390400
transform 1 0 67872 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_602
timestamp 1669390400
transform 1 0 68768 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_604
timestamp 1669390400
transform 1 0 68992 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_611
timestamp 1669390400
transform 1 0 69776 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_618
timestamp 1669390400
transform 1 0 70560 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_622
timestamp 1669390400
transform 1 0 71008 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_624
timestamp 1669390400
transform 1 0 71232 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_638
timestamp 1669390400
transform 1 0 72800 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_641
timestamp 1669390400
transform 1 0 73136 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_648
timestamp 1669390400
transform 1 0 73920 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_652
timestamp 1669390400
transform 1 0 74368 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_666
timestamp 1669390400
transform 1 0 75936 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_680
timestamp 1669390400
transform 1 0 77504 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_687
timestamp 1669390400
transform 1 0 78288 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_2
timestamp 1669390400
transform 1 0 1568 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_4
timestamp 1669390400
transform 1 0 1792 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_7
timestamp 1669390400
transform 1 0 2128 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_22
timestamp 1669390400
transform 1 0 3808 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_32
timestamp 1669390400
transform 1 0 4928 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_34
timestamp 1669390400
transform 1 0 5152 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_37
timestamp 1669390400
transform 1 0 5488 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_44
timestamp 1669390400
transform 1 0 6272 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_52
timestamp 1669390400
transform 1 0 7168 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_56
timestamp 1669390400
transform 1 0 7616 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_58
timestamp 1669390400
transform 1 0 7840 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_72
timestamp 1669390400
transform 1 0 9408 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_88
timestamp 1669390400
transform 1 0 11200 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_92
timestamp 1669390400
transform 1 0 11648 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_94
timestamp 1669390400
transform 1 0 11872 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_97
timestamp 1669390400
transform 1 0 12208 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_101
timestamp 1669390400
transform 1 0 12656 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_105
timestamp 1669390400
transform 1 0 13104 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_108
timestamp 1669390400
transform 1 0 13440 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_119
timestamp 1669390400
transform 1 0 14672 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_126
timestamp 1669390400
transform 1 0 15456 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_130
timestamp 1669390400
transform 1 0 15904 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_134
timestamp 1669390400
transform 1 0 16352 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_136
timestamp 1669390400
transform 1 0 16576 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_139
timestamp 1669390400
transform 1 0 16912 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_143
timestamp 1669390400
transform 1 0 17360 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_150
timestamp 1669390400
transform 1 0 18144 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_176
timestamp 1669390400
transform 1 0 21056 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_179
timestamp 1669390400
transform 1 0 21392 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_190
timestamp 1669390400
transform 1 0 22624 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_206
timestamp 1669390400
transform 1 0 24416 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_220
timestamp 1669390400
transform 1 0 25984 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_230
timestamp 1669390400
transform 1 0 27104 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_238
timestamp 1669390400
transform 1 0 28000 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_241
timestamp 1669390400
transform 1 0 28336 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_247
timestamp 1669390400
transform 1 0 29008 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_250
timestamp 1669390400
transform 1 0 29344 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_259
timestamp 1669390400
transform 1 0 30352 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_263
timestamp 1669390400
transform 1 0 30800 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_266
timestamp 1669390400
transform 1 0 31136 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_282
timestamp 1669390400
transform 1 0 32928 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_286
timestamp 1669390400
transform 1 0 33376 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_288
timestamp 1669390400
transform 1 0 33600 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_297
timestamp 1669390400
transform 1 0 34608 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_299
timestamp 1669390400
transform 1 0 34832 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_302
timestamp 1669390400
transform 1 0 35168 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_309
timestamp 1669390400
transform 1 0 35952 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_313
timestamp 1669390400
transform 1 0 36400 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_317
timestamp 1669390400
transform 1 0 36848 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_321
timestamp 1669390400
transform 1 0 37296 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_339
timestamp 1669390400
transform 1 0 39312 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_346
timestamp 1669390400
transform 1 0 40096 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_352
timestamp 1669390400
transform 1 0 40768 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_356
timestamp 1669390400
transform 1 0 41216 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_372
timestamp 1669390400
transform 1 0 43008 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_376
timestamp 1669390400
transform 1 0 43456 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_379
timestamp 1669390400
transform 1 0 43792 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_386
timestamp 1669390400
transform 1 0 44576 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_392
timestamp 1669390400
transform 1 0 45248 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_408
timestamp 1669390400
transform 1 0 47040 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_416
timestamp 1669390400
transform 1 0 47936 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_420
timestamp 1669390400
transform 1 0 48384 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_429
timestamp 1669390400
transform 1 0 49392 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_437
timestamp 1669390400
transform 1 0 50288 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_441
timestamp 1669390400
transform 1 0 50736 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_445
timestamp 1669390400
transform 1 0 51184 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_460
timestamp 1669390400
transform 1 0 52864 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_463
timestamp 1669390400
transform 1 0 53200 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_477
timestamp 1669390400
transform 1 0 54768 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_481
timestamp 1669390400
transform 1 0 55216 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_489
timestamp 1669390400
transform 1 0 56112 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_502
timestamp 1669390400
transform 1 0 57568 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_510
timestamp 1669390400
transform 1 0 58464 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_512
timestamp 1669390400
transform 1 0 58688 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_515
timestamp 1669390400
transform 1 0 59024 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_523
timestamp 1669390400
transform 1 0 59920 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_529
timestamp 1669390400
transform 1 0 60592 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_531
timestamp 1669390400
transform 1 0 60816 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_534
timestamp 1669390400
transform 1 0 61152 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_549
timestamp 1669390400
transform 1 0 62832 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_564
timestamp 1669390400
transform 1 0 64512 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_568
timestamp 1669390400
transform 1 0 64960 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_576
timestamp 1669390400
transform 1 0 65856 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_580
timestamp 1669390400
transform 1 0 66304 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_584
timestamp 1669390400
transform 1 0 66752 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_588
timestamp 1669390400
transform 1 0 67200 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_592
timestamp 1669390400
transform 1 0 67648 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_600
timestamp 1669390400
transform 1 0 68544 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_602
timestamp 1669390400
transform 1 0 68768 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_605
timestamp 1669390400
transform 1 0 69104 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_609
timestamp 1669390400
transform 1 0 69552 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_616
timestamp 1669390400
transform 1 0 70336 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_631
timestamp 1669390400
transform 1 0 72016 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_635
timestamp 1669390400
transform 1 0 72464 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_643
timestamp 1669390400
transform 1 0 73360 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_649
timestamp 1669390400
transform 1 0 74032 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_659
timestamp 1669390400
transform 1 0 75152 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_673
timestamp 1669390400
transform 1 0 76720 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_676
timestamp 1669390400
transform 1 0 77056 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_685
timestamp 1669390400
transform 1 0 78064 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_687
timestamp 1669390400
transform 1 0 78288 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_2
timestamp 1669390400
transform 1 0 1568 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_17
timestamp 1669390400
transform 1 0 3248 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_44
timestamp 1669390400
transform 1 0 6272 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_60
timestamp 1669390400
transform 1 0 8064 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_70
timestamp 1669390400
transform 1 0 9184 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_73
timestamp 1669390400
transform 1 0 9520 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_87
timestamp 1669390400
transform 1 0 11088 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_91
timestamp 1669390400
transform 1 0 11536 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_95
timestamp 1669390400
transform 1 0 11984 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_102
timestamp 1669390400
transform 1 0 12768 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_127
timestamp 1669390400
transform 1 0 15568 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_133
timestamp 1669390400
transform 1 0 16240 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_137
timestamp 1669390400
transform 1 0 16688 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_141
timestamp 1669390400
transform 1 0 17136 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_144
timestamp 1669390400
transform 1 0 17472 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_147
timestamp 1669390400
transform 1 0 17808 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_154
timestamp 1669390400
transform 1 0 18592 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_161
timestamp 1669390400
transform 1 0 19376 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_167
timestamp 1669390400
transform 1 0 20048 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_174
timestamp 1669390400
transform 1 0 20832 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_178
timestamp 1669390400
transform 1 0 21280 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_182
timestamp 1669390400
transform 1 0 21728 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_184
timestamp 1669390400
transform 1 0 21952 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_190
timestamp 1669390400
transform 1 0 22624 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_194
timestamp 1669390400
transform 1 0 23072 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_198
timestamp 1669390400
transform 1 0 23520 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_206
timestamp 1669390400
transform 1 0 24416 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_212
timestamp 1669390400
transform 1 0 25088 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_215
timestamp 1669390400
transform 1 0 25424 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_228
timestamp 1669390400
transform 1 0 26880 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_232
timestamp 1669390400
transform 1 0 27328 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_239
timestamp 1669390400
transform 1 0 28112 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_265
timestamp 1669390400
transform 1 0 31024 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_281
timestamp 1669390400
transform 1 0 32816 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_283
timestamp 1669390400
transform 1 0 33040 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_286
timestamp 1669390400
transform 1 0 33376 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_300
timestamp 1669390400
transform 1 0 34944 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_308
timestamp 1669390400
transform 1 0 35840 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_311
timestamp 1669390400
transform 1 0 36176 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_319
timestamp 1669390400
transform 1 0 37072 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_322
timestamp 1669390400
transform 1 0 37408 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_330
timestamp 1669390400
transform 1 0 38304 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_333
timestamp 1669390400
transform 1 0 38640 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_348
timestamp 1669390400
transform 1 0 40320 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_352
timestamp 1669390400
transform 1 0 40768 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_354
timestamp 1669390400
transform 1 0 40992 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_357
timestamp 1669390400
transform 1 0 41328 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_365
timestamp 1669390400
transform 1 0 42224 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_369
timestamp 1669390400
transform 1 0 42672 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_373
timestamp 1669390400
transform 1 0 43120 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_375
timestamp 1669390400
transform 1 0 43344 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_389
timestamp 1669390400
transform 1 0 44912 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_405
timestamp 1669390400
transform 1 0 46704 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_413
timestamp 1669390400
transform 1 0 47600 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_417
timestamp 1669390400
transform 1 0 48048 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_419
timestamp 1669390400
transform 1 0 48272 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_425
timestamp 1669390400
transform 1 0 48944 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_428
timestamp 1669390400
transform 1 0 49280 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_442
timestamp 1669390400
transform 1 0 50848 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_458
timestamp 1669390400
transform 1 0 52640 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_460
timestamp 1669390400
transform 1 0 52864 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_463
timestamp 1669390400
transform 1 0 53200 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_477
timestamp 1669390400
transform 1 0 54768 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_483
timestamp 1669390400
transform 1 0 55440 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_489
timestamp 1669390400
transform 1 0 56112 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_496
timestamp 1669390400
transform 1 0 56896 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_499
timestamp 1669390400
transform 1 0 57232 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_508
timestamp 1669390400
transform 1 0 58240 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_512
timestamp 1669390400
transform 1 0 58688 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_514
timestamp 1669390400
transform 1 0 58912 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_527
timestamp 1669390400
transform 1 0 60368 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_537
timestamp 1669390400
transform 1 0 61488 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_544
timestamp 1669390400
transform 1 0 62272 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_548
timestamp 1669390400
transform 1 0 62720 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_557
timestamp 1669390400
transform 1 0 63728 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_561
timestamp 1669390400
transform 1 0 64176 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_567
timestamp 1669390400
transform 1 0 64848 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_570
timestamp 1669390400
transform 1 0 65184 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_579
timestamp 1669390400
transform 1 0 66192 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_581
timestamp 1669390400
transform 1 0 66416 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_587
timestamp 1669390400
transform 1 0 67088 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_599
timestamp 1669390400
transform 1 0 68432 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_603
timestamp 1669390400
transform 1 0 68880 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_607
timestamp 1669390400
transform 1 0 69328 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_611
timestamp 1669390400
transform 1 0 69776 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_626
timestamp 1669390400
transform 1 0 71456 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_634
timestamp 1669390400
transform 1 0 72352 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_638
timestamp 1669390400
transform 1 0 72800 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_641
timestamp 1669390400
transform 1 0 73136 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_647
timestamp 1669390400
transform 1 0 73808 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_651
timestamp 1669390400
transform 1 0 74256 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_655
timestamp 1669390400
transform 1 0 74704 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_670
timestamp 1669390400
transform 1 0 76384 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_684
timestamp 1669390400
transform 1 0 77952 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_2
timestamp 1669390400
transform 1 0 1568 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_4
timestamp 1669390400
transform 1 0 1792 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_7
timestamp 1669390400
transform 1 0 2128 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_11
timestamp 1669390400
transform 1 0 2576 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_15
timestamp 1669390400
transform 1 0 3024 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_27
timestamp 1669390400
transform 1 0 4368 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_34
timestamp 1669390400
transform 1 0 5152 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_37
timestamp 1669390400
transform 1 0 5488 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_53
timestamp 1669390400
transform 1 0 7280 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_59
timestamp 1669390400
transform 1 0 7952 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_66
timestamp 1669390400
transform 1 0 8736 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_70
timestamp 1669390400
transform 1 0 9184 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_86
timestamp 1669390400
transform 1 0 10976 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_90
timestamp 1669390400
transform 1 0 11424 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_94
timestamp 1669390400
transform 1 0 11872 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_104
timestamp 1669390400
transform 1 0 12992 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_108
timestamp 1669390400
transform 1 0 13440 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_114
timestamp 1669390400
transform 1 0 14112 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_118
timestamp 1669390400
transform 1 0 14560 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_122
timestamp 1669390400
transform 1 0 15008 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_126
timestamp 1669390400
transform 1 0 15456 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_130
timestamp 1669390400
transform 1 0 15904 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_134
timestamp 1669390400
transform 1 0 16352 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_144
timestamp 1669390400
transform 1 0 17472 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_146
timestamp 1669390400
transform 1 0 17696 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_149
timestamp 1669390400
transform 1 0 18032 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_156
timestamp 1669390400
transform 1 0 18816 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_163
timestamp 1669390400
transform 1 0 19600 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_175
timestamp 1669390400
transform 1 0 20944 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_179
timestamp 1669390400
transform 1 0 21392 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_182
timestamp 1669390400
transform 1 0 21728 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_186
timestamp 1669390400
transform 1 0 22176 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_202
timestamp 1669390400
transform 1 0 23968 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_206
timestamp 1669390400
transform 1 0 24416 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_221
timestamp 1669390400
transform 1 0 26096 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_229
timestamp 1669390400
transform 1 0 26992 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_233
timestamp 1669390400
transform 1 0 27440 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_239
timestamp 1669390400
transform 1 0 28112 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_247
timestamp 1669390400
transform 1 0 29008 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_250
timestamp 1669390400
transform 1 0 29344 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_256
timestamp 1669390400
transform 1 0 30016 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_260
timestamp 1669390400
transform 1 0 30464 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_268
timestamp 1669390400
transform 1 0 31360 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_271
timestamp 1669390400
transform 1 0 31696 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_297
timestamp 1669390400
transform 1 0 34608 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_307
timestamp 1669390400
transform 1 0 35728 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_311
timestamp 1669390400
transform 1 0 36176 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_318
timestamp 1669390400
transform 1 0 36960 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_321
timestamp 1669390400
transform 1 0 37296 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_335
timestamp 1669390400
transform 1 0 38864 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_339
timestamp 1669390400
transform 1 0 39312 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_341
timestamp 1669390400
transform 1 0 39536 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_354
timestamp 1669390400
transform 1 0 40992 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_364
timestamp 1669390400
transform 1 0 42112 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_371
timestamp 1669390400
transform 1 0 42896 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_386
timestamp 1669390400
transform 1 0 44576 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_392
timestamp 1669390400
transform 1 0 45248 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_401
timestamp 1669390400
transform 1 0 46256 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_417
timestamp 1669390400
transform 1 0 48048 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_421
timestamp 1669390400
transform 1 0 48496 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_423
timestamp 1669390400
transform 1 0 48720 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_436
timestamp 1669390400
transform 1 0 50176 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_446
timestamp 1669390400
transform 1 0 51296 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_454
timestamp 1669390400
transform 1 0 52192 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_460
timestamp 1669390400
transform 1 0 52864 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_463
timestamp 1669390400
transform 1 0 53200 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_477
timestamp 1669390400
transform 1 0 54768 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_487
timestamp 1669390400
transform 1 0 55888 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_491
timestamp 1669390400
transform 1 0 56336 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_495
timestamp 1669390400
transform 1 0 56784 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_498
timestamp 1669390400
transform 1 0 57120 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_514
timestamp 1669390400
transform 1 0 58912 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_528
timestamp 1669390400
transform 1 0 60480 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_534
timestamp 1669390400
transform 1 0 61152 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_543
timestamp 1669390400
transform 1 0 62160 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_547
timestamp 1669390400
transform 1 0 62608 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_551
timestamp 1669390400
transform 1 0 63056 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_555
timestamp 1669390400
transform 1 0 63504 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_565
timestamp 1669390400
transform 1 0 64624 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_575
timestamp 1669390400
transform 1 0 65744 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_591
timestamp 1669390400
transform 1 0 67536 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_601
timestamp 1669390400
transform 1 0 68656 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_605
timestamp 1669390400
transform 1 0 69104 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_608
timestamp 1669390400
transform 1 0 69440 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_612
timestamp 1669390400
transform 1 0 69888 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_618
timestamp 1669390400
transform 1 0 70560 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_632
timestamp 1669390400
transform 1 0 72128 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_636
timestamp 1669390400
transform 1 0 72576 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_652
timestamp 1669390400
transform 1 0 74368 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_673
timestamp 1669390400
transform 1 0 76720 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_676
timestamp 1669390400
transform 1 0 77056 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_681
timestamp 1669390400
transform 1 0 77616 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_685
timestamp 1669390400
transform 1 0 78064 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_687
timestamp 1669390400
transform 1 0 78288 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_2
timestamp 1669390400
transform 1 0 1568 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_5
timestamp 1669390400
transform 1 0 1904 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_12
timestamp 1669390400
transform 1 0 2688 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_26
timestamp 1669390400
transform 1 0 4256 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_33
timestamp 1669390400
transform 1 0 5040 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_37
timestamp 1669390400
transform 1 0 5488 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_41
timestamp 1669390400
transform 1 0 5936 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_49
timestamp 1669390400
transform 1 0 6832 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_53
timestamp 1669390400
transform 1 0 7280 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_67
timestamp 1669390400
transform 1 0 8848 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_73
timestamp 1669390400
transform 1 0 9520 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_79
timestamp 1669390400
transform 1 0 10192 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_87
timestamp 1669390400
transform 1 0 11088 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_97
timestamp 1669390400
transform 1 0 12208 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_122
timestamp 1669390400
transform 1 0 15008 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_126
timestamp 1669390400
transform 1 0 15456 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_130
timestamp 1669390400
transform 1 0 15904 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_134
timestamp 1669390400
transform 1 0 16352 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_141
timestamp 1669390400
transform 1 0 17136 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_144
timestamp 1669390400
transform 1 0 17472 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_146
timestamp 1669390400
transform 1 0 17696 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_149
timestamp 1669390400
transform 1 0 18032 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_161
timestamp 1669390400
transform 1 0 19376 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_167
timestamp 1669390400
transform 1 0 20048 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_171
timestamp 1669390400
transform 1 0 20496 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_196
timestamp 1669390400
transform 1 0 23296 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_204
timestamp 1669390400
transform 1 0 24192 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_206
timestamp 1669390400
transform 1 0 24416 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_212
timestamp 1669390400
transform 1 0 25088 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_215
timestamp 1669390400
transform 1 0 25424 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_224
timestamp 1669390400
transform 1 0 26432 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_228
timestamp 1669390400
transform 1 0 26880 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_234
timestamp 1669390400
transform 1 0 27552 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_260
timestamp 1669390400
transform 1 0 30464 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_276
timestamp 1669390400
transform 1 0 32256 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_286
timestamp 1669390400
transform 1 0 33376 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_290
timestamp 1669390400
transform 1 0 33824 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_294
timestamp 1669390400
transform 1 0 34272 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_304
timestamp 1669390400
transform 1 0 35392 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_314
timestamp 1669390400
transform 1 0 36512 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_318
timestamp 1669390400
transform 1 0 36960 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_322
timestamp 1669390400
transform 1 0 37408 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_329
timestamp 1669390400
transform 1 0 38192 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_344
timestamp 1669390400
transform 1 0 39872 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_354
timestamp 1669390400
transform 1 0 40992 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_357
timestamp 1669390400
transform 1 0 41328 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_365
timestamp 1669390400
transform 1 0 42224 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_369
timestamp 1669390400
transform 1 0 42672 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_371
timestamp 1669390400
transform 1 0 42896 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_380
timestamp 1669390400
transform 1 0 43904 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_382
timestamp 1669390400
transform 1 0 44128 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_395
timestamp 1669390400
transform 1 0 45584 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_404
timestamp 1669390400
transform 1 0 46592 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_425
timestamp 1669390400
transform 1 0 48944 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_428
timestamp 1669390400
transform 1 0 49280 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_441
timestamp 1669390400
transform 1 0 50736 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_457
timestamp 1669390400
transform 1 0 52528 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_465
timestamp 1669390400
transform 1 0 53424 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_475
timestamp 1669390400
transform 1 0 54544 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_485
timestamp 1669390400
transform 1 0 55664 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_493
timestamp 1669390400
transform 1 0 56560 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_499
timestamp 1669390400
transform 1 0 57232 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_515
timestamp 1669390400
transform 1 0 59024 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_529
timestamp 1669390400
transform 1 0 60592 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_537
timestamp 1669390400
transform 1 0 61488 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_543
timestamp 1669390400
transform 1 0 62160 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_558
timestamp 1669390400
transform 1 0 63840 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_562
timestamp 1669390400
transform 1 0 64288 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_564
timestamp 1669390400
transform 1 0 64512 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_567
timestamp 1669390400
transform 1 0 64848 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_570
timestamp 1669390400
transform 1 0 65184 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_576
timestamp 1669390400
transform 1 0 65856 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_580
timestamp 1669390400
transform 1 0 66304 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_584
timestamp 1669390400
transform 1 0 66752 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_591
timestamp 1669390400
transform 1 0 67536 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_595
timestamp 1669390400
transform 1 0 67984 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_599
timestamp 1669390400
transform 1 0 68432 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_607
timestamp 1669390400
transform 1 0 69328 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_613
timestamp 1669390400
transform 1 0 70000 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_615
timestamp 1669390400
transform 1 0 70224 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_618
timestamp 1669390400
transform 1 0 70560 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_622
timestamp 1669390400
transform 1 0 71008 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_628
timestamp 1669390400
transform 1 0 71680 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_638
timestamp 1669390400
transform 1 0 72800 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_641
timestamp 1669390400
transform 1 0 73136 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_647
timestamp 1669390400
transform 1 0 73808 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_655
timestamp 1669390400
transform 1 0 74704 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_664
timestamp 1669390400
transform 1 0 75712 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_679
timestamp 1669390400
transform 1 0 77392 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_687
timestamp 1669390400
transform 1 0 78288 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_2
timestamp 1669390400
transform 1 0 1568 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_17
timestamp 1669390400
transform 1 0 3248 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_24
timestamp 1669390400
transform 1 0 4032 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_31
timestamp 1669390400
transform 1 0 4816 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_37
timestamp 1669390400
transform 1 0 5488 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_40
timestamp 1669390400
transform 1 0 5824 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_44
timestamp 1669390400
transform 1 0 6272 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_48
timestamp 1669390400
transform 1 0 6720 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_54
timestamp 1669390400
transform 1 0 7392 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_68
timestamp 1669390400
transform 1 0 8960 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_78
timestamp 1669390400
transform 1 0 10080 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_94
timestamp 1669390400
transform 1 0 11872 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_105
timestamp 1669390400
transform 1 0 13104 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_108
timestamp 1669390400
transform 1 0 13440 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_114
timestamp 1669390400
transform 1 0 14112 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_121
timestamp 1669390400
transform 1 0 14896 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_125
timestamp 1669390400
transform 1 0 15344 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_129
timestamp 1669390400
transform 1 0 15792 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_133
timestamp 1669390400
transform 1 0 16240 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_137
timestamp 1669390400
transform 1 0 16688 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_141
timestamp 1669390400
transform 1 0 17136 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_167
timestamp 1669390400
transform 1 0 20048 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_171
timestamp 1669390400
transform 1 0 20496 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_175
timestamp 1669390400
transform 1 0 20944 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_179
timestamp 1669390400
transform 1 0 21392 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_182
timestamp 1669390400
transform 1 0 21728 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_186
timestamp 1669390400
transform 1 0 22176 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_190
timestamp 1669390400
transform 1 0 22624 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_198
timestamp 1669390400
transform 1 0 23520 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_205
timestamp 1669390400
transform 1 0 24304 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_209
timestamp 1669390400
transform 1 0 24752 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_223
timestamp 1669390400
transform 1 0 26320 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_231
timestamp 1669390400
transform 1 0 27216 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_233
timestamp 1669390400
transform 1 0 27440 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_240
timestamp 1669390400
transform 1 0 28224 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_247
timestamp 1669390400
transform 1 0 29008 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_250
timestamp 1669390400
transform 1 0 29344 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_266
timestamp 1669390400
transform 1 0 31136 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_270
timestamp 1669390400
transform 1 0 31584 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_295
timestamp 1669390400
transform 1 0 34384 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_305
timestamp 1669390400
transform 1 0 35504 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_309
timestamp 1669390400
transform 1 0 35952 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_313
timestamp 1669390400
transform 1 0 36400 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_317
timestamp 1669390400
transform 1 0 36848 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_321
timestamp 1669390400
transform 1 0 37296 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_325
timestamp 1669390400
transform 1 0 37744 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_339
timestamp 1669390400
transform 1 0 39312 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_346
timestamp 1669390400
transform 1 0 40096 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_353
timestamp 1669390400
transform 1 0 40880 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_357
timestamp 1669390400
transform 1 0 41328 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_361
timestamp 1669390400
transform 1 0 41776 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_386
timestamp 1669390400
transform 1 0 44576 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_392
timestamp 1669390400
transform 1 0 45248 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_394
timestamp 1669390400
transform 1 0 45472 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_408
timestamp 1669390400
transform 1 0 47040 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_416
timestamp 1669390400
transform 1 0 47936 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_418
timestamp 1669390400
transform 1 0 48160 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_431
timestamp 1669390400
transform 1 0 49616 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_438
timestamp 1669390400
transform 1 0 50400 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_445
timestamp 1669390400
transform 1 0 51184 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_449
timestamp 1669390400
transform 1 0 51632 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_453
timestamp 1669390400
transform 1 0 52080 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_463
timestamp 1669390400
transform 1 0 53200 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_476
timestamp 1669390400
transform 1 0 54656 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_480
timestamp 1669390400
transform 1 0 55104 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_488
timestamp 1669390400
transform 1 0 56000 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_502
timestamp 1669390400
transform 1 0 57568 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_509
timestamp 1669390400
transform 1 0 58352 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_517
timestamp 1669390400
transform 1 0 59248 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_531
timestamp 1669390400
transform 1 0 60816 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_534
timestamp 1669390400
transform 1 0 61152 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_543
timestamp 1669390400
transform 1 0 62160 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_550
timestamp 1669390400
transform 1 0 62944 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_554
timestamp 1669390400
transform 1 0 63392 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_563
timestamp 1669390400
transform 1 0 64400 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_571
timestamp 1669390400
transform 1 0 65296 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_575
timestamp 1669390400
transform 1 0 65744 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_590
timestamp 1669390400
transform 1 0 67424 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_600
timestamp 1669390400
transform 1 0 68544 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_602
timestamp 1669390400
transform 1 0 68768 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_605
timestamp 1669390400
transform 1 0 69104 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_619
timestamp 1669390400
transform 1 0 70672 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_623
timestamp 1669390400
transform 1 0 71120 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_636
timestamp 1669390400
transform 1 0 72576 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_650
timestamp 1669390400
transform 1 0 74144 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_654
timestamp 1669390400
transform 1 0 74592 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_670
timestamp 1669390400
transform 1 0 76384 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_676
timestamp 1669390400
transform 1 0 77056 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_682
timestamp 1669390400
transform 1 0 77728 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_686
timestamp 1669390400
transform 1 0 78176 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_2
timestamp 1669390400
transform 1 0 1568 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_6
timestamp 1669390400
transform 1 0 2016 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_10
timestamp 1669390400
transform 1 0 2464 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_18
timestamp 1669390400
transform 1 0 3360 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_30
timestamp 1669390400
transform 1 0 4704 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_34
timestamp 1669390400
transform 1 0 5152 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_38
timestamp 1669390400
transform 1 0 5600 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_42
timestamp 1669390400
transform 1 0 6048 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_58
timestamp 1669390400
transform 1 0 7840 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_70
timestamp 1669390400
transform 1 0 9184 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_73
timestamp 1669390400
transform 1 0 9520 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_76
timestamp 1669390400
transform 1 0 9856 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_84
timestamp 1669390400
transform 1 0 10752 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_93
timestamp 1669390400
transform 1 0 11760 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_120
timestamp 1669390400
transform 1 0 14784 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_126
timestamp 1669390400
transform 1 0 15456 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_130
timestamp 1669390400
transform 1 0 15904 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_134
timestamp 1669390400
transform 1 0 16352 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_141
timestamp 1669390400
transform 1 0 17136 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_144
timestamp 1669390400
transform 1 0 17472 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_157
timestamp 1669390400
transform 1 0 18928 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_164
timestamp 1669390400
transform 1 0 19712 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_168
timestamp 1669390400
transform 1 0 20160 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_170
timestamp 1669390400
transform 1 0 20384 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_173
timestamp 1669390400
transform 1 0 20720 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_184
timestamp 1669390400
transform 1 0 21952 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_190
timestamp 1669390400
transform 1 0 22624 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_194
timestamp 1669390400
transform 1 0 23072 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_209
timestamp 1669390400
transform 1 0 24752 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_215
timestamp 1669390400
transform 1 0 25424 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_231
timestamp 1669390400
transform 1 0 27216 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_235
timestamp 1669390400
transform 1 0 27664 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_245
timestamp 1669390400
transform 1 0 28784 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_253
timestamp 1669390400
transform 1 0 29680 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_255
timestamp 1669390400
transform 1 0 29904 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_258
timestamp 1669390400
transform 1 0 30240 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_262
timestamp 1669390400
transform 1 0 30688 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_266
timestamp 1669390400
transform 1 0 31136 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_268
timestamp 1669390400
transform 1 0 31360 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_279
timestamp 1669390400
transform 1 0 32592 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_283
timestamp 1669390400
transform 1 0 33040 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_286
timestamp 1669390400
transform 1 0 33376 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_290
timestamp 1669390400
transform 1 0 33824 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_300
timestamp 1669390400
transform 1 0 34944 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_304
timestamp 1669390400
transform 1 0 35392 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_308
timestamp 1669390400
transform 1 0 35840 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_324
timestamp 1669390400
transform 1 0 37632 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_340
timestamp 1669390400
transform 1 0 39424 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_344
timestamp 1669390400
transform 1 0 39872 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_352
timestamp 1669390400
transform 1 0 40768 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_354
timestamp 1669390400
transform 1 0 40992 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_357
timestamp 1669390400
transform 1 0 41328 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_365
timestamp 1669390400
transform 1 0 42224 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_369
timestamp 1669390400
transform 1 0 42672 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_377
timestamp 1669390400
transform 1 0 43568 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_384
timestamp 1669390400
transform 1 0 44352 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_388
timestamp 1669390400
transform 1 0 44800 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_392
timestamp 1669390400
transform 1 0 45248 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_395
timestamp 1669390400
transform 1 0 45584 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_403
timestamp 1669390400
transform 1 0 46480 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_405
timestamp 1669390400
transform 1 0 46704 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_408
timestamp 1669390400
transform 1 0 47040 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_412
timestamp 1669390400
transform 1 0 47488 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_414
timestamp 1669390400
transform 1 0 47712 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_423
timestamp 1669390400
transform 1 0 48720 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_425
timestamp 1669390400
transform 1 0 48944 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_428
timestamp 1669390400
transform 1 0 49280 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_436
timestamp 1669390400
transform 1 0 50176 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_443
timestamp 1669390400
transform 1 0 50960 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_447
timestamp 1669390400
transform 1 0 51408 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_451
timestamp 1669390400
transform 1 0 51856 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_477
timestamp 1669390400
transform 1 0 54768 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_493
timestamp 1669390400
transform 1 0 56560 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_499
timestamp 1669390400
transform 1 0 57232 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_502
timestamp 1669390400
transform 1 0 57568 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_518
timestamp 1669390400
transform 1 0 59360 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_522
timestamp 1669390400
transform 1 0 59808 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_532
timestamp 1669390400
transform 1 0 60928 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_536
timestamp 1669390400
transform 1 0 61376 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_542
timestamp 1669390400
transform 1 0 62048 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_546
timestamp 1669390400
transform 1 0 62496 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_560
timestamp 1669390400
transform 1 0 64064 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_564
timestamp 1669390400
transform 1 0 64512 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_570
timestamp 1669390400
transform 1 0 65184 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_573
timestamp 1669390400
transform 1 0 65520 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_577
timestamp 1669390400
transform 1 0 65968 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_593
timestamp 1669390400
transform 1 0 67760 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_601
timestamp 1669390400
transform 1 0 68656 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_610
timestamp 1669390400
transform 1 0 69664 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_618
timestamp 1669390400
transform 1 0 70560 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_625
timestamp 1669390400
transform 1 0 71344 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_629
timestamp 1669390400
transform 1 0 71792 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_633
timestamp 1669390400
transform 1 0 72240 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_638
timestamp 1669390400
transform 1 0 72800 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_641
timestamp 1669390400
transform 1 0 73136 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_647
timestamp 1669390400
transform 1 0 73808 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_651
timestamp 1669390400
transform 1 0 74256 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_655
timestamp 1669390400
transform 1 0 74704 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_659
timestamp 1669390400
transform 1 0 75152 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_662
timestamp 1669390400
transform 1 0 75488 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_676
timestamp 1669390400
transform 1 0 77056 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_683
timestamp 1669390400
transform 1 0 77840 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_687
timestamp 1669390400
transform 1 0 78288 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_2
timestamp 1669390400
transform 1 0 1568 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_6
timestamp 1669390400
transform 1 0 2016 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_9
timestamp 1669390400
transform 1 0 2352 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_24
timestamp 1669390400
transform 1 0 4032 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_32
timestamp 1669390400
transform 1 0 4928 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_34
timestamp 1669390400
transform 1 0 5152 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_37
timestamp 1669390400
transform 1 0 5488 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_39
timestamp 1669390400
transform 1 0 5712 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_53
timestamp 1669390400
transform 1 0 7280 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_60
timestamp 1669390400
transform 1 0 8064 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_68
timestamp 1669390400
transform 1 0 8960 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_72
timestamp 1669390400
transform 1 0 9408 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_79
timestamp 1669390400
transform 1 0 10192 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_83
timestamp 1669390400
transform 1 0 10640 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_85
timestamp 1669390400
transform 1 0 10864 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_96
timestamp 1669390400
transform 1 0 12096 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_103
timestamp 1669390400
transform 1 0 12880 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_105
timestamp 1669390400
transform 1 0 13104 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_108
timestamp 1669390400
transform 1 0 13440 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_114
timestamp 1669390400
transform 1 0 14112 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_118
timestamp 1669390400
transform 1 0 14560 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_122
timestamp 1669390400
transform 1 0 15008 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_126
timestamp 1669390400
transform 1 0 15456 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_128
timestamp 1669390400
transform 1 0 15680 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_131
timestamp 1669390400
transform 1 0 16016 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_135
timestamp 1669390400
transform 1 0 16464 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_139
timestamp 1669390400
transform 1 0 16912 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_143
timestamp 1669390400
transform 1 0 17360 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_154
timestamp 1669390400
transform 1 0 18592 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_158
timestamp 1669390400
transform 1 0 19040 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_161
timestamp 1669390400
transform 1 0 19376 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_165
timestamp 1669390400
transform 1 0 19824 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_176
timestamp 1669390400
transform 1 0 21056 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_179
timestamp 1669390400
transform 1 0 21392 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_188
timestamp 1669390400
transform 1 0 22400 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_192
timestamp 1669390400
transform 1 0 22848 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_198
timestamp 1669390400
transform 1 0 23520 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_212
timestamp 1669390400
transform 1 0 25088 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_216
timestamp 1669390400
transform 1 0 25536 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_226
timestamp 1669390400
transform 1 0 26656 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_233
timestamp 1669390400
transform 1 0 27440 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_241
timestamp 1669390400
transform 1 0 28336 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_247
timestamp 1669390400
transform 1 0 29008 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_250
timestamp 1669390400
transform 1 0 29344 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_256
timestamp 1669390400
transform 1 0 30016 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_260
timestamp 1669390400
transform 1 0 30464 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_267
timestamp 1669390400
transform 1 0 31248 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_281
timestamp 1669390400
transform 1 0 32816 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_285
timestamp 1669390400
transform 1 0 33264 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_292
timestamp 1669390400
transform 1 0 34048 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_299
timestamp 1669390400
transform 1 0 34832 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_306
timestamp 1669390400
transform 1 0 35616 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_310
timestamp 1669390400
transform 1 0 36064 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_318
timestamp 1669390400
transform 1 0 36960 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_321
timestamp 1669390400
transform 1 0 37296 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_325
timestamp 1669390400
transform 1 0 37744 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_339
timestamp 1669390400
transform 1 0 39312 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_350
timestamp 1669390400
transform 1 0 40544 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_352
timestamp 1669390400
transform 1 0 40768 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_355
timestamp 1669390400
transform 1 0 41104 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_362
timestamp 1669390400
transform 1 0 41888 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_366
timestamp 1669390400
transform 1 0 42336 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_370
timestamp 1669390400
transform 1 0 42784 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_386
timestamp 1669390400
transform 1 0 44576 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_392
timestamp 1669390400
transform 1 0 45248 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_396
timestamp 1669390400
transform 1 0 45696 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_398
timestamp 1669390400
transform 1 0 45920 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_407
timestamp 1669390400
transform 1 0 46928 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_411
timestamp 1669390400
transform 1 0 47376 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_417
timestamp 1669390400
transform 1 0 48048 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_427
timestamp 1669390400
transform 1 0 49168 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_431
timestamp 1669390400
transform 1 0 49616 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_435
timestamp 1669390400
transform 1 0 50064 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_439
timestamp 1669390400
transform 1 0 50512 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_442
timestamp 1669390400
transform 1 0 50848 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_444
timestamp 1669390400
transform 1 0 51072 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_453
timestamp 1669390400
transform 1 0 52080 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_463
timestamp 1669390400
transform 1 0 53200 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_471
timestamp 1669390400
transform 1 0 54096 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_477
timestamp 1669390400
transform 1 0 54768 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_481
timestamp 1669390400
transform 1 0 55216 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_488
timestamp 1669390400
transform 1 0 56000 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_498
timestamp 1669390400
transform 1 0 57120 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_506
timestamp 1669390400
transform 1 0 58016 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_527
timestamp 1669390400
transform 1 0 60368 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_531
timestamp 1669390400
transform 1 0 60816 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_534
timestamp 1669390400
transform 1 0 61152 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_544
timestamp 1669390400
transform 1 0 62272 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_554
timestamp 1669390400
transform 1 0 63392 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_558
timestamp 1669390400
transform 1 0 63840 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_569
timestamp 1669390400
transform 1 0 65072 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_573
timestamp 1669390400
transform 1 0 65520 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_587
timestamp 1669390400
transform 1 0 67088 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_605
timestamp 1669390400
transform 1 0 69104 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_618
timestamp 1669390400
transform 1 0 70560 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_622
timestamp 1669390400
transform 1 0 71008 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_626
timestamp 1669390400
transform 1 0 71456 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_630
timestamp 1669390400
transform 1 0 71904 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_644
timestamp 1669390400
transform 1 0 73472 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_658
timestamp 1669390400
transform 1 0 75040 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_660
timestamp 1669390400
transform 1 0 75264 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_663
timestamp 1669390400
transform 1 0 75600 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_670
timestamp 1669390400
transform 1 0 76384 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_676
timestamp 1669390400
transform 1 0 77056 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_682
timestamp 1669390400
transform 1 0 77728 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_686
timestamp 1669390400
transform 1 0 78176 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_2
timestamp 1669390400
transform 1 0 1568 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_17
timestamp 1669390400
transform 1 0 3248 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_25
timestamp 1669390400
transform 1 0 4144 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_33
timestamp 1669390400
transform 1 0 5040 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_17_37
timestamp 1669390400
transform 1 0 5488 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_45
timestamp 1669390400
transform 1 0 6384 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_17_60
timestamp 1669390400
transform 1 0 8064 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_70
timestamp 1669390400
transform 1 0 9184 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_73
timestamp 1669390400
transform 1 0 9520 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_17_82
timestamp 1669390400
transform 1 0 10528 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_90
timestamp 1669390400
transform 1 0 11424 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_96
timestamp 1669390400
transform 1 0 12096 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_100
timestamp 1669390400
transform 1 0 12544 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_104
timestamp 1669390400
transform 1 0 12992 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_111
timestamp 1669390400
transform 1 0 13776 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_113
timestamp 1669390400
transform 1 0 14000 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_116
timestamp 1669390400
transform 1 0 14336 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_17_120
timestamp 1669390400
transform 1 0 14784 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_130
timestamp 1669390400
transform 1 0 15904 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_134
timestamp 1669390400
transform 1 0 16352 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_141
timestamp 1669390400
transform 1 0 17136 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_144
timestamp 1669390400
transform 1 0 17472 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_155
timestamp 1669390400
transform 1 0 18704 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_161
timestamp 1669390400
transform 1 0 19376 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_165
timestamp 1669390400
transform 1 0 19824 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_175
timestamp 1669390400
transform 1 0 20944 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_190
timestamp 1669390400
transform 1 0 22624 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_194
timestamp 1669390400
transform 1 0 23072 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_198
timestamp 1669390400
transform 1 0 23520 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_202
timestamp 1669390400
transform 1 0 23968 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_212
timestamp 1669390400
transform 1 0 25088 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_215
timestamp 1669390400
transform 1 0 25424 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_17_240
timestamp 1669390400
transform 1 0 28224 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_250
timestamp 1669390400
transform 1 0 29344 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_254
timestamp 1669390400
transform 1 0 29792 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_261
timestamp 1669390400
transform 1 0 30576 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_276
timestamp 1669390400
transform 1 0 32256 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_283
timestamp 1669390400
transform 1 0 33040 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_286
timestamp 1669390400
transform 1 0 33376 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_17_289
timestamp 1669390400
transform 1 0 33712 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_310
timestamp 1669390400
transform 1 0 36064 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_331
timestamp 1669390400
transform 1 0 38416 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_335
timestamp 1669390400
transform 1 0 38864 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_339
timestamp 1669390400
transform 1 0 39312 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_343
timestamp 1669390400
transform 1 0 39760 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_347
timestamp 1669390400
transform 1 0 40208 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_354
timestamp 1669390400
transform 1 0 40992 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_357
timestamp 1669390400
transform 1 0 41328 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_359
timestamp 1669390400
transform 1 0 41552 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_17_383
timestamp 1669390400
transform 1 0 44240 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_391
timestamp 1669390400
transform 1 0 45136 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_397
timestamp 1669390400
transform 1 0 45808 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_404
timestamp 1669390400
transform 1 0 46592 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_410
timestamp 1669390400
transform 1 0 47264 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_420
timestamp 1669390400
transform 1 0 48384 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_424
timestamp 1669390400
transform 1 0 48832 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_428
timestamp 1669390400
transform 1 0 49280 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_440
timestamp 1669390400
transform 1 0 50624 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_455
timestamp 1669390400
transform 1 0 52304 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_463
timestamp 1669390400
transform 1 0 53200 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_469
timestamp 1669390400
transform 1 0 53872 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_479
timestamp 1669390400
transform 1 0 54992 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_481
timestamp 1669390400
transform 1 0 55216 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_494
timestamp 1669390400
transform 1 0 56672 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_496
timestamp 1669390400
transform 1 0 56896 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_499
timestamp 1669390400
transform 1 0 57232 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_17_508
timestamp 1669390400
transform 1 0 58240 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_524
timestamp 1669390400
transform 1 0 60032 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_528
timestamp 1669390400
transform 1 0 60480 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_532
timestamp 1669390400
transform 1 0 60928 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_545
timestamp 1669390400
transform 1 0 62384 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_549
timestamp 1669390400
transform 1 0 62832 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_553
timestamp 1669390400
transform 1 0 63280 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_557
timestamp 1669390400
transform 1 0 63728 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_567
timestamp 1669390400
transform 1 0 64848 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_570
timestamp 1669390400
transform 1 0 65184 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_583
timestamp 1669390400
transform 1 0 66640 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_17_593
timestamp 1669390400
transform 1 0 67760 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_601
timestamp 1669390400
transform 1 0 68656 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_605
timestamp 1669390400
transform 1 0 69104 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_17_615
timestamp 1669390400
transform 1 0 70224 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_17_631
timestamp 1669390400
transform 1 0 72016 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_641
timestamp 1669390400
transform 1 0 73136 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_643
timestamp 1669390400
transform 1 0 73360 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_652
timestamp 1669390400
transform 1 0 74368 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_670
timestamp 1669390400
transform 1 0 76384 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_684
timestamp 1669390400
transform 1 0 77952 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_2
timestamp 1669390400
transform 1 0 1568 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_4
timestamp 1669390400
transform 1 0 1792 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_11
timestamp 1669390400
transform 1 0 2576 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_26
timestamp 1669390400
transform 1 0 4256 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_30
timestamp 1669390400
transform 1 0 4704 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_34
timestamp 1669390400
transform 1 0 5152 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_37
timestamp 1669390400
transform 1 0 5488 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_42
timestamp 1669390400
transform 1 0 6048 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_46
timestamp 1669390400
transform 1 0 6496 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_56
timestamp 1669390400
transform 1 0 7616 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_58
timestamp 1669390400
transform 1 0 7840 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_61
timestamp 1669390400
transform 1 0 8176 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_68
timestamp 1669390400
transform 1 0 8960 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_80
timestamp 1669390400
transform 1 0 10304 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_18_84
timestamp 1669390400
transform 1 0 10752 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_92
timestamp 1669390400
transform 1 0 11648 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_95
timestamp 1669390400
transform 1 0 11984 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_102
timestamp 1669390400
transform 1 0 12768 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_108
timestamp 1669390400
transform 1 0 13440 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_114
timestamp 1669390400
transform 1 0 14112 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_118
timestamp 1669390400
transform 1 0 14560 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_18_122
timestamp 1669390400
transform 1 0 15008 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_130
timestamp 1669390400
transform 1 0 15904 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_155
timestamp 1669390400
transform 1 0 18704 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_162
timestamp 1669390400
transform 1 0 19488 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_166
timestamp 1669390400
transform 1 0 19936 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_172
timestamp 1669390400
transform 1 0 20608 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_176
timestamp 1669390400
transform 1 0 21056 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_179
timestamp 1669390400
transform 1 0 21392 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_181
timestamp 1669390400
transform 1 0 21616 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_187
timestamp 1669390400
transform 1 0 22288 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_189
timestamp 1669390400
transform 1 0 22512 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_18_192
timestamp 1669390400
transform 1 0 22848 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_18_208
timestamp 1669390400
transform 1 0 24640 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_216
timestamp 1669390400
transform 1 0 25536 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_219
timestamp 1669390400
transform 1 0 25872 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_18_229
timestamp 1669390400
transform 1 0 26992 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_237
timestamp 1669390400
transform 1 0 27888 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_241
timestamp 1669390400
transform 1 0 28336 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_247
timestamp 1669390400
transform 1 0 29008 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_250
timestamp 1669390400
transform 1 0 29344 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_254
timestamp 1669390400
transform 1 0 29792 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_261
timestamp 1669390400
transform 1 0 30576 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_282
timestamp 1669390400
transform 1 0 32928 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_286
timestamp 1669390400
transform 1 0 33376 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_290
timestamp 1669390400
transform 1 0 33824 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_294
timestamp 1669390400
transform 1 0 34272 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_298
timestamp 1669390400
transform 1 0 34720 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_305
timestamp 1669390400
transform 1 0 35504 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_307
timestamp 1669390400
transform 1 0 35728 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_310
timestamp 1669390400
transform 1 0 36064 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_317
timestamp 1669390400
transform 1 0 36848 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_321
timestamp 1669390400
transform 1 0 37296 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_334
timestamp 1669390400
transform 1 0 38752 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_344
timestamp 1669390400
transform 1 0 39872 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_351
timestamp 1669390400
transform 1 0 40656 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_355
timestamp 1669390400
transform 1 0 41104 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_18_365
timestamp 1669390400
transform 1 0 42224 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_381
timestamp 1669390400
transform 1 0 44016 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_385
timestamp 1669390400
transform 1 0 44464 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_389
timestamp 1669390400
transform 1 0 44912 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_392
timestamp 1669390400
transform 1 0 45248 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_406
timestamp 1669390400
transform 1 0 46816 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_18_416
timestamp 1669390400
transform 1 0 47936 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_424
timestamp 1669390400
transform 1 0 48832 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_427
timestamp 1669390400
transform 1 0 49168 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_431
timestamp 1669390400
transform 1 0 49616 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_435
timestamp 1669390400
transform 1 0 50064 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_439
timestamp 1669390400
transform 1 0 50512 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_443
timestamp 1669390400
transform 1 0 50960 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_450
timestamp 1669390400
transform 1 0 51744 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_458
timestamp 1669390400
transform 1 0 52640 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_460
timestamp 1669390400
transform 1 0 52864 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_463
timestamp 1669390400
transform 1 0 53200 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_18_466
timestamp 1669390400
transform 1 0 53536 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_498
timestamp 1669390400
transform 1 0 57120 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_502
timestamp 1669390400
transform 1 0 57568 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_504
timestamp 1669390400
transform 1 0 57792 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_18_513
timestamp 1669390400
transform 1 0 58800 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_529
timestamp 1669390400
transform 1 0 60592 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_531
timestamp 1669390400
transform 1 0 60816 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_534
timestamp 1669390400
transform 1 0 61152 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_544
timestamp 1669390400
transform 1 0 62272 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_548
timestamp 1669390400
transform 1 0 62720 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_552
timestamp 1669390400
transform 1 0 63168 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_556
timestamp 1669390400
transform 1 0 63616 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_560
timestamp 1669390400
transform 1 0 64064 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_564
timestamp 1669390400
transform 1 0 64512 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_566
timestamp 1669390400
transform 1 0 64736 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_569
timestamp 1669390400
transform 1 0 65072 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_573
timestamp 1669390400
transform 1 0 65520 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_18_577
timestamp 1669390400
transform 1 0 65968 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_18_593
timestamp 1669390400
transform 1 0 67760 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_601
timestamp 1669390400
transform 1 0 68656 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_605
timestamp 1669390400
transform 1 0 69104 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_619
timestamp 1669390400
transform 1 0 70672 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_18_629
timestamp 1669390400
transform 1 0 71792 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_637
timestamp 1669390400
transform 1 0 72688 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_641
timestamp 1669390400
transform 1 0 73136 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_645
timestamp 1669390400
transform 1 0 73584 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_649
timestamp 1669390400
transform 1 0 74032 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_656
timestamp 1669390400
transform 1 0 74816 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_670
timestamp 1669390400
transform 1 0 76384 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_676
timestamp 1669390400
transform 1 0 77056 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_682
timestamp 1669390400
transform 1 0 77728 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_686
timestamp 1669390400
transform 1 0 78176 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_2
timestamp 1669390400
transform 1 0 1568 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_6
timestamp 1669390400
transform 1 0 2016 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_10
timestamp 1669390400
transform 1 0 2464 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_18
timestamp 1669390400
transform 1 0 3360 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_25
timestamp 1669390400
transform 1 0 4144 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_29
timestamp 1669390400
transform 1 0 4592 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_42
timestamp 1669390400
transform 1 0 6048 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_19_49
timestamp 1669390400
transform 1 0 6832 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_59
timestamp 1669390400
transform 1 0 7952 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_63
timestamp 1669390400
transform 1 0 8400 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_70
timestamp 1669390400
transform 1 0 9184 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_73
timestamp 1669390400
transform 1 0 9520 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_79
timestamp 1669390400
transform 1 0 10192 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_83
timestamp 1669390400
transform 1 0 10640 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_110
timestamp 1669390400
transform 1 0 13664 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_120
timestamp 1669390400
transform 1 0 14784 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_126
timestamp 1669390400
transform 1 0 15456 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_130
timestamp 1669390400
transform 1 0 15904 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_134
timestamp 1669390400
transform 1 0 16352 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_141
timestamp 1669390400
transform 1 0 17136 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_144
timestamp 1669390400
transform 1 0 17472 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_150
timestamp 1669390400
transform 1 0 18144 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_157
timestamp 1669390400
transform 1 0 18928 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_163
timestamp 1669390400
transform 1 0 19600 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_170
timestamp 1669390400
transform 1 0 20384 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_174
timestamp 1669390400
transform 1 0 20832 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_190
timestamp 1669390400
transform 1 0 22624 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_200
timestamp 1669390400
transform 1 0 23744 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_208
timestamp 1669390400
transform 1 0 24640 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_212
timestamp 1669390400
transform 1 0 25088 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_215
timestamp 1669390400
transform 1 0 25424 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_224
timestamp 1669390400
transform 1 0 26432 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_228
timestamp 1669390400
transform 1 0 26880 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_232
timestamp 1669390400
transform 1 0 27328 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_239
timestamp 1669390400
transform 1 0 28112 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_245
timestamp 1669390400
transform 1 0 28784 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_247
timestamp 1669390400
transform 1 0 29008 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_271
timestamp 1669390400
transform 1 0 31696 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_281
timestamp 1669390400
transform 1 0 32816 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_283
timestamp 1669390400
transform 1 0 33040 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_19_286
timestamp 1669390400
transform 1 0 33376 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_294
timestamp 1669390400
transform 1 0 34272 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_300
timestamp 1669390400
transform 1 0 34944 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_310
timestamp 1669390400
transform 1 0 36064 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_312
timestamp 1669390400
transform 1 0 36288 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_318
timestamp 1669390400
transform 1 0 36960 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_324
timestamp 1669390400
transform 1 0 37632 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_328
timestamp 1669390400
transform 1 0 38080 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_339
timestamp 1669390400
transform 1 0 39312 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_354
timestamp 1669390400
transform 1 0 40992 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_357
timestamp 1669390400
transform 1 0 41328 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_359
timestamp 1669390400
transform 1 0 41552 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_373
timestamp 1669390400
transform 1 0 43120 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_19_381
timestamp 1669390400
transform 1 0 44016 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_391
timestamp 1669390400
transform 1 0 45136 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_398
timestamp 1669390400
transform 1 0 45920 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_402
timestamp 1669390400
transform 1 0 46368 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_19_415
timestamp 1669390400
transform 1 0 47824 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_423
timestamp 1669390400
transform 1 0 48720 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_425
timestamp 1669390400
transform 1 0 48944 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_428
timestamp 1669390400
transform 1 0 49280 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_437
timestamp 1669390400
transform 1 0 50288 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_439
timestamp 1669390400
transform 1 0 50512 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_442
timestamp 1669390400
transform 1 0 50848 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_453
timestamp 1669390400
transform 1 0 52080 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_457
timestamp 1669390400
transform 1 0 52528 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_461
timestamp 1669390400
transform 1 0 52976 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_474
timestamp 1669390400
transform 1 0 54432 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_19_484
timestamp 1669390400
transform 1 0 55552 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_492
timestamp 1669390400
transform 1 0 56448 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_496
timestamp 1669390400
transform 1 0 56896 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_499
timestamp 1669390400
transform 1 0 57232 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_511
timestamp 1669390400
transform 1 0 58576 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_19_523
timestamp 1669390400
transform 1 0 59920 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_531
timestamp 1669390400
transform 1 0 60816 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_533
timestamp 1669390400
transform 1 0 61040 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_19_547
timestamp 1669390400
transform 1 0 62608 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_555
timestamp 1669390400
transform 1 0 63504 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_567
timestamp 1669390400
transform 1 0 64848 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_570
timestamp 1669390400
transform 1 0 65184 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_581
timestamp 1669390400
transform 1 0 66416 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_585
timestamp 1669390400
transform 1 0 66864 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_19_589
timestamp 1669390400
transform 1 0 67312 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_597
timestamp 1669390400
transform 1 0 68208 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_600
timestamp 1669390400
transform 1 0 68544 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_610
timestamp 1669390400
transform 1 0 69664 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_624
timestamp 1669390400
transform 1 0 71232 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_634
timestamp 1669390400
transform 1 0 72352 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_638
timestamp 1669390400
transform 1 0 72800 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_641
timestamp 1669390400
transform 1 0 73136 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_651
timestamp 1669390400
transform 1 0 74256 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_677
timestamp 1669390400
transform 1 0 77168 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_687
timestamp 1669390400
transform 1 0 78288 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_2
timestamp 1669390400
transform 1 0 1568 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_17
timestamp 1669390400
transform 1 0 3248 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_25
timestamp 1669390400
transform 1 0 4144 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_29
timestamp 1669390400
transform 1 0 4592 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_34
timestamp 1669390400
transform 1 0 5152 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_37
timestamp 1669390400
transform 1 0 5488 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_20_50
timestamp 1669390400
transform 1 0 6944 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_58
timestamp 1669390400
transform 1 0 7840 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_60
timestamp 1669390400
transform 1 0 8064 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_69
timestamp 1669390400
transform 1 0 9072 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_20_81
timestamp 1669390400
transform 1 0 10416 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_20_97
timestamp 1669390400
transform 1 0 12208 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_105
timestamp 1669390400
transform 1 0 13104 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_108
timestamp 1669390400
transform 1 0 13440 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_117
timestamp 1669390400
transform 1 0 14448 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_20_121
timestamp 1669390400
transform 1 0 14896 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_129
timestamp 1669390400
transform 1 0 15792 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_131
timestamp 1669390400
transform 1 0 16016 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_134
timestamp 1669390400
transform 1 0 16352 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_146
timestamp 1669390400
transform 1 0 17696 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_157
timestamp 1669390400
transform 1 0 18928 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_170
timestamp 1669390400
transform 1 0 20384 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_176
timestamp 1669390400
transform 1 0 21056 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_179
timestamp 1669390400
transform 1 0 21392 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_182
timestamp 1669390400
transform 1 0 21728 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_188
timestamp 1669390400
transform 1 0 22400 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_192
timestamp 1669390400
transform 1 0 22848 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_218
timestamp 1669390400
transform 1 0 25760 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_225
timestamp 1669390400
transform 1 0 26544 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_227
timestamp 1669390400
transform 1 0 26768 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_230
timestamp 1669390400
transform 1 0 27104 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_237
timestamp 1669390400
transform 1 0 27888 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_239
timestamp 1669390400
transform 1 0 28112 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_242
timestamp 1669390400
transform 1 0 28448 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_244
timestamp 1669390400
transform 1 0 28672 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_247
timestamp 1669390400
transform 1 0 29008 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_250
timestamp 1669390400
transform 1 0 29344 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_252
timestamp 1669390400
transform 1 0 29568 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_255
timestamp 1669390400
transform 1 0 29904 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_265
timestamp 1669390400
transform 1 0 31024 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_272
timestamp 1669390400
transform 1 0 31808 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_20_276
timestamp 1669390400
transform 1 0 32256 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_284
timestamp 1669390400
transform 1 0 33152 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_300
timestamp 1669390400
transform 1 0 34944 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_314
timestamp 1669390400
transform 1 0 36512 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_318
timestamp 1669390400
transform 1 0 36960 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_321
timestamp 1669390400
transform 1 0 37296 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_323
timestamp 1669390400
transform 1 0 37520 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_326
timestamp 1669390400
transform 1 0 37856 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_330
timestamp 1669390400
transform 1 0 38304 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_334
timestamp 1669390400
transform 1 0 38752 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_338
timestamp 1669390400
transform 1 0 39200 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_345
timestamp 1669390400
transform 1 0 39984 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_352
timestamp 1669390400
transform 1 0 40768 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_356
timestamp 1669390400
transform 1 0 41216 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_360
timestamp 1669390400
transform 1 0 41664 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_364
timestamp 1669390400
transform 1 0 42112 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_371
timestamp 1669390400
transform 1 0 42896 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_375
timestamp 1669390400
transform 1 0 43344 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_382
timestamp 1669390400
transform 1 0 44128 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_384
timestamp 1669390400
transform 1 0 44352 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_387
timestamp 1669390400
transform 1 0 44688 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_389
timestamp 1669390400
transform 1 0 44912 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_392
timestamp 1669390400
transform 1 0 45248 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_20_395
timestamp 1669390400
transform 1 0 45584 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_411
timestamp 1669390400
transform 1 0 47376 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_439
timestamp 1669390400
transform 1 0 50512 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_446
timestamp 1669390400
transform 1 0 51296 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_450
timestamp 1669390400
transform 1 0 51744 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_454
timestamp 1669390400
transform 1 0 52192 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_457
timestamp 1669390400
transform 1 0 52528 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_463
timestamp 1669390400
transform 1 0 53200 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_20_477
timestamp 1669390400
transform 1 0 54768 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_498
timestamp 1669390400
transform 1 0 57120 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_508
timestamp 1669390400
transform 1 0 58240 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_512
timestamp 1669390400
transform 1 0 58688 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_514
timestamp 1669390400
transform 1 0 58912 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_528
timestamp 1669390400
transform 1 0 60480 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_534
timestamp 1669390400
transform 1 0 61152 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_20_542
timestamp 1669390400
transform 1 0 62048 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_550
timestamp 1669390400
transform 1 0 62944 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_553
timestamp 1669390400
transform 1 0 63280 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_557
timestamp 1669390400
transform 1 0 63728 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_567
timestamp 1669390400
transform 1 0 64848 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_593
timestamp 1669390400
transform 1 0 67760 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_597
timestamp 1669390400
transform 1 0 68208 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_599
timestamp 1669390400
transform 1 0 68432 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_602
timestamp 1669390400
transform 1 0 68768 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_605
timestamp 1669390400
transform 1 0 69104 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_611
timestamp 1669390400
transform 1 0 69776 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_626
timestamp 1669390400
transform 1 0 71456 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_20_630
timestamp 1669390400
transform 1 0 71904 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_646
timestamp 1669390400
transform 1 0 73696 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_650
timestamp 1669390400
transform 1 0 74144 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_654
timestamp 1669390400
transform 1 0 74592 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_670
timestamp 1669390400
transform 1 0 76384 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_676
timestamp 1669390400
transform 1 0 77056 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_20_679
timestamp 1669390400
transform 1 0 77392 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_687
timestamp 1669390400
transform 1 0 78288 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_2
timestamp 1669390400
transform 1 0 1568 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_5
timestamp 1669390400
transform 1 0 1904 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_15
timestamp 1669390400
transform 1 0 3024 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_27
timestamp 1669390400
transform 1 0 4368 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_31
timestamp 1669390400
transform 1 0 4816 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_35
timestamp 1669390400
transform 1 0 5264 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_37
timestamp 1669390400
transform 1 0 5488 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_21_46
timestamp 1669390400
transform 1 0 6496 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_21_62
timestamp 1669390400
transform 1 0 8288 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_70
timestamp 1669390400
transform 1 0 9184 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_73
timestamp 1669390400
transform 1 0 9520 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_21_97
timestamp 1669390400
transform 1 0 12208 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_118
timestamp 1669390400
transform 1 0 14560 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_21_125
timestamp 1669390400
transform 1 0 15344 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_133
timestamp 1669390400
transform 1 0 16240 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_137
timestamp 1669390400
transform 1 0 16688 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_141
timestamp 1669390400
transform 1 0 17136 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_144
timestamp 1669390400
transform 1 0 17472 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_169
timestamp 1669390400
transform 1 0 20272 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_173
timestamp 1669390400
transform 1 0 20720 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_176
timestamp 1669390400
transform 1 0 21056 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_180
timestamp 1669390400
transform 1 0 21504 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_184
timestamp 1669390400
transform 1 0 21952 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_193
timestamp 1669390400
transform 1 0 22960 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_197
timestamp 1669390400
transform 1 0 23408 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_200
timestamp 1669390400
transform 1 0 23744 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_210
timestamp 1669390400
transform 1 0 24864 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_212
timestamp 1669390400
transform 1 0 25088 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_215
timestamp 1669390400
transform 1 0 25424 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_221
timestamp 1669390400
transform 1 0 26096 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_225
timestamp 1669390400
transform 1 0 26544 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_229
timestamp 1669390400
transform 1 0 26992 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_236
timestamp 1669390400
transform 1 0 27776 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_243
timestamp 1669390400
transform 1 0 28560 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_249
timestamp 1669390400
transform 1 0 29232 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_256
timestamp 1669390400
transform 1 0 30016 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_21_268
timestamp 1669390400
transform 1 0 31360 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_286
timestamp 1669390400
transform 1 0 33376 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_288
timestamp 1669390400
transform 1 0 33600 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_291
timestamp 1669390400
transform 1 0 33936 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_297
timestamp 1669390400
transform 1 0 34608 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_311
timestamp 1669390400
transform 1 0 36176 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_315
timestamp 1669390400
transform 1 0 36624 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_317
timestamp 1669390400
transform 1 0 36848 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_21_320
timestamp 1669390400
transform 1 0 37184 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_328
timestamp 1669390400
transform 1 0 38080 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_332
timestamp 1669390400
transform 1 0 38528 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_335
timestamp 1669390400
transform 1 0 38864 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_339
timestamp 1669390400
transform 1 0 39312 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_346
timestamp 1669390400
transform 1 0 40096 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_354
timestamp 1669390400
transform 1 0 40992 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_357
timestamp 1669390400
transform 1 0 41328 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_21_364
timestamp 1669390400
transform 1 0 42112 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_372
timestamp 1669390400
transform 1 0 43008 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_374
timestamp 1669390400
transform 1 0 43232 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_377
timestamp 1669390400
transform 1 0 43568 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_387
timestamp 1669390400
transform 1 0 44688 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_397
timestamp 1669390400
transform 1 0 45808 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_404
timestamp 1669390400
transform 1 0 46592 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_21_408
timestamp 1669390400
transform 1 0 47040 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_416
timestamp 1669390400
transform 1 0 47936 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_418
timestamp 1669390400
transform 1 0 48160 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_425
timestamp 1669390400
transform 1 0 48944 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_428
timestamp 1669390400
transform 1 0 49280 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_21_435
timestamp 1669390400
transform 1 0 50064 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_21_451
timestamp 1669390400
transform 1 0 51856 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_459
timestamp 1669390400
transform 1 0 52752 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_468
timestamp 1669390400
transform 1 0 53760 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_21_476
timestamp 1669390400
transform 1 0 54656 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_484
timestamp 1669390400
transform 1 0 55552 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_493
timestamp 1669390400
transform 1 0 56560 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_21_499
timestamp 1669390400
transform 1 0 57232 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_515
timestamp 1669390400
transform 1 0 59024 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_519
timestamp 1669390400
transform 1 0 59472 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_21_528
timestamp 1669390400
transform 1 0 60480 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_549
timestamp 1669390400
transform 1 0 62832 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_21_553
timestamp 1669390400
transform 1 0 63280 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_563
timestamp 1669390400
transform 1 0 64400 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_567
timestamp 1669390400
transform 1 0 64848 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_570
timestamp 1669390400
transform 1 0 65184 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_573
timestamp 1669390400
transform 1 0 65520 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_577
timestamp 1669390400
transform 1 0 65968 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_581
timestamp 1669390400
transform 1 0 66416 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_592
timestamp 1669390400
transform 1 0 67648 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_596
timestamp 1669390400
transform 1 0 68096 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_602
timestamp 1669390400
transform 1 0 68768 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_606
timestamp 1669390400
transform 1 0 69216 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_612
timestamp 1669390400
transform 1 0 69888 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_618
timestamp 1669390400
transform 1 0 70560 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_632
timestamp 1669390400
transform 1 0 72128 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_636
timestamp 1669390400
transform 1 0 72576 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_638
timestamp 1669390400
transform 1 0 72800 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_641
timestamp 1669390400
transform 1 0 73136 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_644
timestamp 1669390400
transform 1 0 73472 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_646
timestamp 1669390400
transform 1 0 73696 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_655
timestamp 1669390400
transform 1 0 74704 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_670
timestamp 1669390400
transform 1 0 76384 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_682
timestamp 1669390400
transform 1 0 77728 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_686
timestamp 1669390400
transform 1 0 78176 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_2
timestamp 1669390400
transform 1 0 1568 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_17
timestamp 1669390400
transform 1 0 3248 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_27
timestamp 1669390400
transform 1 0 4368 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_34
timestamp 1669390400
transform 1 0 5152 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_37
timestamp 1669390400
transform 1 0 5488 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_40
timestamp 1669390400
transform 1 0 5824 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_44
timestamp 1669390400
transform 1 0 6272 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_48
timestamp 1669390400
transform 1 0 6720 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_58
timestamp 1669390400
transform 1 0 7840 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_62
timestamp 1669390400
transform 1 0 8288 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_64
timestamp 1669390400
transform 1 0 8512 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_67
timestamp 1669390400
transform 1 0 8848 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_74
timestamp 1669390400
transform 1 0 9632 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_78
timestamp 1669390400
transform 1 0 10080 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_85
timestamp 1669390400
transform 1 0 10864 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_89
timestamp 1669390400
transform 1 0 11312 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_22_93
timestamp 1669390400
transform 1 0 11760 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_101
timestamp 1669390400
transform 1 0 12656 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_105
timestamp 1669390400
transform 1 0 13104 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_108
timestamp 1669390400
transform 1 0 13440 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_22_117
timestamp 1669390400
transform 1 0 14448 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_125
timestamp 1669390400
transform 1 0 15344 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_127
timestamp 1669390400
transform 1 0 15568 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_152
timestamp 1669390400
transform 1 0 18368 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_156
timestamp 1669390400
transform 1 0 18816 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_158
timestamp 1669390400
transform 1 0 19040 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_161
timestamp 1669390400
transform 1 0 19376 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_165
timestamp 1669390400
transform 1 0 19824 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_169
timestamp 1669390400
transform 1 0 20272 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_176
timestamp 1669390400
transform 1 0 21056 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_179
timestamp 1669390400
transform 1 0 21392 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_189
timestamp 1669390400
transform 1 0 22512 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_195
timestamp 1669390400
transform 1 0 23184 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_205
timestamp 1669390400
transform 1 0 24304 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_209
timestamp 1669390400
transform 1 0 24752 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_213
timestamp 1669390400
transform 1 0 25200 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_217
timestamp 1669390400
transform 1 0 25648 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_221
timestamp 1669390400
transform 1 0 26096 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_228
timestamp 1669390400
transform 1 0 26880 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_240
timestamp 1669390400
transform 1 0 28224 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_247
timestamp 1669390400
transform 1 0 29008 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_250
timestamp 1669390400
transform 1 0 29344 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_253
timestamp 1669390400
transform 1 0 29680 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_22_278
timestamp 1669390400
transform 1 0 32480 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_286
timestamp 1669390400
transform 1 0 33376 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_292
timestamp 1669390400
transform 1 0 34048 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_302
timestamp 1669390400
transform 1 0 35168 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_317
timestamp 1669390400
transform 1 0 36848 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_321
timestamp 1669390400
transform 1 0 37296 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_323
timestamp 1669390400
transform 1 0 37520 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_326
timestamp 1669390400
transform 1 0 37856 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_330
timestamp 1669390400
transform 1 0 38304 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_341
timestamp 1669390400
transform 1 0 39536 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_356
timestamp 1669390400
transform 1 0 41216 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_22_366
timestamp 1669390400
transform 1 0 42336 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_382
timestamp 1669390400
transform 1 0 44128 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_389
timestamp 1669390400
transform 1 0 44912 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_392
timestamp 1669390400
transform 1 0 45248 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_22_405
timestamp 1669390400
transform 1 0 46704 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_413
timestamp 1669390400
transform 1 0 47600 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_415
timestamp 1669390400
transform 1 0 47824 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_22_440
timestamp 1669390400
transform 1 0 50624 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_448
timestamp 1669390400
transform 1 0 51520 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_452
timestamp 1669390400
transform 1 0 51968 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_460
timestamp 1669390400
transform 1 0 52864 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_463
timestamp 1669390400
transform 1 0 53200 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_476
timestamp 1669390400
transform 1 0 54656 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_480
timestamp 1669390400
transform 1 0 55104 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_22_493
timestamp 1669390400
transform 1 0 56560 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_501
timestamp 1669390400
transform 1 0 57456 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_503
timestamp 1669390400
transform 1 0 57680 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_516
timestamp 1669390400
transform 1 0 59136 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_531
timestamp 1669390400
transform 1 0 60816 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_534
timestamp 1669390400
transform 1 0 61152 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_536
timestamp 1669390400
transform 1 0 61376 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_556
timestamp 1669390400
transform 1 0 63616 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_560
timestamp 1669390400
transform 1 0 64064 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_566
timestamp 1669390400
transform 1 0 64736 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_568
timestamp 1669390400
transform 1 0 64960 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_574
timestamp 1669390400
transform 1 0 65632 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_599
timestamp 1669390400
transform 1 0 68432 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_605
timestamp 1669390400
transform 1 0 69104 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_613
timestamp 1669390400
transform 1 0 70000 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_625
timestamp 1669390400
transform 1 0 71344 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_635
timestamp 1669390400
transform 1 0 72464 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_639
timestamp 1669390400
transform 1 0 72912 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_643
timestamp 1669390400
transform 1 0 73360 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_652
timestamp 1669390400
transform 1 0 74368 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_22_666
timestamp 1669390400
transform 1 0 75936 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_676
timestamp 1669390400
transform 1 0 77056 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_685
timestamp 1669390400
transform 1 0 78064 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_687
timestamp 1669390400
transform 1 0 78288 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_2
timestamp 1669390400
transform 1 0 1568 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_8
timestamp 1669390400
transform 1 0 2240 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_15
timestamp 1669390400
transform 1 0 3024 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_40
timestamp 1669390400
transform 1 0 5824 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_44
timestamp 1669390400
transform 1 0 6272 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_48
timestamp 1669390400
transform 1 0 6720 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_55
timestamp 1669390400
transform 1 0 7504 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_59
timestamp 1669390400
transform 1 0 7952 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_63
timestamp 1669390400
transform 1 0 8400 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_65
timestamp 1669390400
transform 1 0 8624 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_70
timestamp 1669390400
transform 1 0 9184 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_73
timestamp 1669390400
transform 1 0 9520 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_23_82
timestamp 1669390400
transform 1 0 10528 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_98
timestamp 1669390400
transform 1 0 12320 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_23_111
timestamp 1669390400
transform 1 0 13776 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_119
timestamp 1669390400
transform 1 0 14672 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_123
timestamp 1669390400
transform 1 0 15120 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_126
timestamp 1669390400
transform 1 0 15456 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_130
timestamp 1669390400
transform 1 0 15904 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_134
timestamp 1669390400
transform 1 0 16352 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_141
timestamp 1669390400
transform 1 0 17136 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_144
timestamp 1669390400
transform 1 0 17472 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_155
timestamp 1669390400
transform 1 0 18704 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_159
timestamp 1669390400
transform 1 0 19152 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_161
timestamp 1669390400
transform 1 0 19376 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_164
timestamp 1669390400
transform 1 0 19712 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_168
timestamp 1669390400
transform 1 0 20160 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_175
timestamp 1669390400
transform 1 0 20944 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_182
timestamp 1669390400
transform 1 0 21728 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_192
timestamp 1669390400
transform 1 0 22848 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_196
timestamp 1669390400
transform 1 0 23296 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_200
timestamp 1669390400
transform 1 0 23744 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_204
timestamp 1669390400
transform 1 0 24192 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_208
timestamp 1669390400
transform 1 0 24640 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_212
timestamp 1669390400
transform 1 0 25088 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_215
timestamp 1669390400
transform 1 0 25424 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_225
timestamp 1669390400
transform 1 0 26544 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_229
timestamp 1669390400
transform 1 0 26992 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_23_255
timestamp 1669390400
transform 1 0 29904 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_271
timestamp 1669390400
transform 1 0 31696 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_276
timestamp 1669390400
transform 1 0 32256 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_283
timestamp 1669390400
transform 1 0 33040 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_23_286
timestamp 1669390400
transform 1 0 33376 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_302
timestamp 1669390400
transform 1 0 35168 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_319
timestamp 1669390400
transform 1 0 37072 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_329
timestamp 1669390400
transform 1 0 38192 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_333
timestamp 1669390400
transform 1 0 38640 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_335
timestamp 1669390400
transform 1 0 38864 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_338
timestamp 1669390400
transform 1 0 39200 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_342
timestamp 1669390400
transform 1 0 39648 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_349
timestamp 1669390400
transform 1 0 40432 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_353
timestamp 1669390400
transform 1 0 40880 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_357
timestamp 1669390400
transform 1 0 41328 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_23_369
timestamp 1669390400
transform 1 0 42672 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_377
timestamp 1669390400
transform 1 0 43568 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_386
timestamp 1669390400
transform 1 0 44576 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_390
timestamp 1669390400
transform 1 0 45024 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_394
timestamp 1669390400
transform 1 0 45472 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_23_398
timestamp 1669390400
transform 1 0 45920 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_406
timestamp 1669390400
transform 1 0 46816 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_410
timestamp 1669390400
transform 1 0 47264 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_412
timestamp 1669390400
transform 1 0 47488 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_418
timestamp 1669390400
transform 1 0 48160 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_425
timestamp 1669390400
transform 1 0 48944 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_428
timestamp 1669390400
transform 1 0 49280 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_23_437
timestamp 1669390400
transform 1 0 50288 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_23_453
timestamp 1669390400
transform 1 0 52080 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_461
timestamp 1669390400
transform 1 0 52976 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_463
timestamp 1669390400
transform 1 0 53200 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_470
timestamp 1669390400
transform 1 0 53984 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_23_474
timestamp 1669390400
transform 1 0 54432 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_492
timestamp 1669390400
transform 1 0 56448 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_496
timestamp 1669390400
transform 1 0 56896 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_499
timestamp 1669390400
transform 1 0 57232 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_509
timestamp 1669390400
transform 1 0 58352 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_513
timestamp 1669390400
transform 1 0 58800 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_517
timestamp 1669390400
transform 1 0 59248 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_521
timestamp 1669390400
transform 1 0 59696 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_525
timestamp 1669390400
transform 1 0 60144 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_533
timestamp 1669390400
transform 1 0 61040 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_23_540
timestamp 1669390400
transform 1 0 61824 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_548
timestamp 1669390400
transform 1 0 62720 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_554
timestamp 1669390400
transform 1 0 63392 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_564
timestamp 1669390400
transform 1 0 64512 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_570
timestamp 1669390400
transform 1 0 65184 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_576
timestamp 1669390400
transform 1 0 65856 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_578
timestamp 1669390400
transform 1 0 66080 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_587
timestamp 1669390400
transform 1 0 67088 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_591
timestamp 1669390400
transform 1 0 67536 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_23_595
timestamp 1669390400
transform 1 0 67984 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_603
timestamp 1669390400
transform 1 0 68880 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_609
timestamp 1669390400
transform 1 0 69552 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_613
timestamp 1669390400
transform 1 0 70000 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_617
timestamp 1669390400
transform 1 0 70448 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_23_630
timestamp 1669390400
transform 1 0 71904 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_638
timestamp 1669390400
transform 1 0 72800 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_23_641
timestamp 1669390400
transform 1 0 73136 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_649
timestamp 1669390400
transform 1 0 74032 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_651
timestamp 1669390400
transform 1 0 74256 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_654
timestamp 1669390400
transform 1 0 74592 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_670
timestamp 1669390400
transform 1 0 76384 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_23_677
timestamp 1669390400
transform 1 0 77168 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_685
timestamp 1669390400
transform 1 0 78064 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_687
timestamp 1669390400
transform 1 0 78288 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_2
timestamp 1669390400
transform 1 0 1568 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_8
timestamp 1669390400
transform 1 0 2240 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_12
timestamp 1669390400
transform 1 0 2688 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_16
timestamp 1669390400
transform 1 0 3136 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_24
timestamp 1669390400
transform 1 0 4032 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_31
timestamp 1669390400
transform 1 0 4816 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_37
timestamp 1669390400
transform 1 0 5488 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_40
timestamp 1669390400
transform 1 0 5824 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_44
timestamp 1669390400
transform 1 0 6272 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_51
timestamp 1669390400
transform 1 0 7056 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_53
timestamp 1669390400
transform 1 0 7280 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_66
timestamp 1669390400
transform 1 0 8736 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_24_81
timestamp 1669390400
transform 1 0 10416 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_89
timestamp 1669390400
transform 1 0 11312 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_93
timestamp 1669390400
transform 1 0 11760 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_97
timestamp 1669390400
transform 1 0 12208 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_105
timestamp 1669390400
transform 1 0 13104 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_108
timestamp 1669390400
transform 1 0 13440 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_117
timestamp 1669390400
transform 1 0 14448 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_124
timestamp 1669390400
transform 1 0 15232 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_128
timestamp 1669390400
transform 1 0 15680 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_132
timestamp 1669390400
transform 1 0 16128 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_138
timestamp 1669390400
transform 1 0 16800 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_140
timestamp 1669390400
transform 1 0 17024 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_24_143
timestamp 1669390400
transform 1 0 17360 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_159
timestamp 1669390400
transform 1 0 19152 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_163
timestamp 1669390400
transform 1 0 19600 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_174
timestamp 1669390400
transform 1 0 20832 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_176
timestamp 1669390400
transform 1 0 21056 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_179
timestamp 1669390400
transform 1 0 21392 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_181
timestamp 1669390400
transform 1 0 21616 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_184
timestamp 1669390400
transform 1 0 21952 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_24_188
timestamp 1669390400
transform 1 0 22400 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_206
timestamp 1669390400
transform 1 0 24416 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_210
timestamp 1669390400
transform 1 0 24864 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_220
timestamp 1669390400
transform 1 0 25984 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_227
timestamp 1669390400
transform 1 0 26768 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_231
timestamp 1669390400
transform 1 0 27216 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_237
timestamp 1669390400
transform 1 0 27888 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_241
timestamp 1669390400
transform 1 0 28336 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_245
timestamp 1669390400
transform 1 0 28784 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_247
timestamp 1669390400
transform 1 0 29008 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_24_250
timestamp 1669390400
transform 1 0 29344 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_266
timestamp 1669390400
transform 1 0 31136 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_270
timestamp 1669390400
transform 1 0 31584 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_284
timestamp 1669390400
transform 1 0 33152 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_24_294
timestamp 1669390400
transform 1 0 34272 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_310
timestamp 1669390400
transform 1 0 36064 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_314
timestamp 1669390400
transform 1 0 36512 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_318
timestamp 1669390400
transform 1 0 36960 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_321
timestamp 1669390400
transform 1 0 37296 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_24_334
timestamp 1669390400
transform 1 0 38752 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_342
timestamp 1669390400
transform 1 0 39648 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_357
timestamp 1669390400
transform 1 0 41328 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_24_361
timestamp 1669390400
transform 1 0 41776 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_369
timestamp 1669390400
transform 1 0 42672 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_371
timestamp 1669390400
transform 1 0 42896 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_374
timestamp 1669390400
transform 1 0 43232 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_389
timestamp 1669390400
transform 1 0 44912 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_392
timestamp 1669390400
transform 1 0 45248 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_406
timestamp 1669390400
transform 1 0 46816 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_412
timestamp 1669390400
transform 1 0 47488 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_24_433
timestamp 1669390400
transform 1 0 49840 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_441
timestamp 1669390400
transform 1 0 50736 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_445
timestamp 1669390400
transform 1 0 51184 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_452
timestamp 1669390400
transform 1 0 51968 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_459
timestamp 1669390400
transform 1 0 52752 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_463
timestamp 1669390400
transform 1 0 53200 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_476
timestamp 1669390400
transform 1 0 54656 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_480
timestamp 1669390400
transform 1 0 55104 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_484
timestamp 1669390400
transform 1 0 55552 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_494
timestamp 1669390400
transform 1 0 56672 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_498
timestamp 1669390400
transform 1 0 57120 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_505
timestamp 1669390400
transform 1 0 57904 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_512
timestamp 1669390400
transform 1 0 58688 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_519
timestamp 1669390400
transform 1 0 59472 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_523
timestamp 1669390400
transform 1 0 59920 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_527
timestamp 1669390400
transform 1 0 60368 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_531
timestamp 1669390400
transform 1 0 60816 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_534
timestamp 1669390400
transform 1 0 61152 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_24_537
timestamp 1669390400
transform 1 0 61488 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_553
timestamp 1669390400
transform 1 0 63280 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_559
timestamp 1669390400
transform 1 0 63952 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_563
timestamp 1669390400
transform 1 0 64400 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_570
timestamp 1669390400
transform 1 0 65184 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_577
timestamp 1669390400
transform 1 0 65968 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_581
timestamp 1669390400
transform 1 0 66416 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_592
timestamp 1669390400
transform 1 0 67648 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_596
timestamp 1669390400
transform 1 0 68096 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_600
timestamp 1669390400
transform 1 0 68544 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_602
timestamp 1669390400
transform 1 0 68768 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_24_605
timestamp 1669390400
transform 1 0 69104 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_613
timestamp 1669390400
transform 1 0 70000 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_617
timestamp 1669390400
transform 1 0 70448 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_620
timestamp 1669390400
transform 1 0 70784 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_627
timestamp 1669390400
transform 1 0 71568 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_641
timestamp 1669390400
transform 1 0 73136 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_645
timestamp 1669390400
transform 1 0 73584 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_658
timestamp 1669390400
transform 1 0 75040 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_673
timestamp 1669390400
transform 1 0 76720 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_676
timestamp 1669390400
transform 1 0 77056 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_685
timestamp 1669390400
transform 1 0 78064 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_687
timestamp 1669390400
transform 1 0 78288 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_25_2
timestamp 1669390400
transform 1 0 1568 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_23
timestamp 1669390400
transform 1 0 3920 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_31
timestamp 1669390400
transform 1 0 4816 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_35
timestamp 1669390400
transform 1 0 5264 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_39
timestamp 1669390400
transform 1 0 5712 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_54
timestamp 1669390400
transform 1 0 7392 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_58
timestamp 1669390400
transform 1 0 7840 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_25_62
timestamp 1669390400
transform 1 0 8288 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_70
timestamp 1669390400
transform 1 0 9184 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_73
timestamp 1669390400
transform 1 0 9520 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_25_79
timestamp 1669390400
transform 1 0 10192 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_87
timestamp 1669390400
transform 1 0 11088 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_25_91
timestamp 1669390400
transform 1 0 11536 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_99
timestamp 1669390400
transform 1 0 12432 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_101
timestamp 1669390400
transform 1 0 12656 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_126
timestamp 1669390400
transform 1 0 15456 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_141
timestamp 1669390400
transform 1 0 17136 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_144
timestamp 1669390400
transform 1 0 17472 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_148
timestamp 1669390400
transform 1 0 17920 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_151
timestamp 1669390400
transform 1 0 18256 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_155
timestamp 1669390400
transform 1 0 18704 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_162
timestamp 1669390400
transform 1 0 19488 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_25_188
timestamp 1669390400
transform 1 0 22400 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_196
timestamp 1669390400
transform 1 0 23296 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_200
timestamp 1669390400
transform 1 0 23744 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_210
timestamp 1669390400
transform 1 0 24864 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_212
timestamp 1669390400
transform 1 0 25088 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_215
timestamp 1669390400
transform 1 0 25424 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_221
timestamp 1669390400
transform 1 0 26096 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_228
timestamp 1669390400
transform 1 0 26880 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_232
timestamp 1669390400
transform 1 0 27328 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_25_256
timestamp 1669390400
transform 1 0 30016 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_25_272
timestamp 1669390400
transform 1 0 31808 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_280
timestamp 1669390400
transform 1 0 32704 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_286
timestamp 1669390400
transform 1 0 33376 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_299
timestamp 1669390400
transform 1 0 34832 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_25_303
timestamp 1669390400
transform 1 0 35280 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_313
timestamp 1669390400
transform 1 0 36400 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_323
timestamp 1669390400
transform 1 0 37520 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_327
timestamp 1669390400
transform 1 0 37968 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_330
timestamp 1669390400
transform 1 0 38304 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_345
timestamp 1669390400
transform 1 0 39984 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_352
timestamp 1669390400
transform 1 0 40768 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_354
timestamp 1669390400
transform 1 0 40992 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_357
timestamp 1669390400
transform 1 0 41328 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_25_364
timestamp 1669390400
transform 1 0 42112 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_380
timestamp 1669390400
transform 1 0 43904 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_384
timestamp 1669390400
transform 1 0 44352 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_386
timestamp 1669390400
transform 1 0 44576 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_402
timestamp 1669390400
transform 1 0 46368 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_412
timestamp 1669390400
transform 1 0 47488 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_420
timestamp 1669390400
transform 1 0 48384 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_424
timestamp 1669390400
transform 1 0 48832 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_428
timestamp 1669390400
transform 1 0 49280 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_441
timestamp 1669390400
transform 1 0 50736 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_445
timestamp 1669390400
transform 1 0 51184 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_449
timestamp 1669390400
transform 1 0 51632 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_462
timestamp 1669390400
transform 1 0 53088 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_25_474
timestamp 1669390400
transform 1 0 54432 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_482
timestamp 1669390400
transform 1 0 55328 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_486
timestamp 1669390400
transform 1 0 55776 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_496
timestamp 1669390400
transform 1 0 56896 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_499
timestamp 1669390400
transform 1 0 57232 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_505
timestamp 1669390400
transform 1 0 57904 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_509
timestamp 1669390400
transform 1 0 58352 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_519
timestamp 1669390400
transform 1 0 59472 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_531
timestamp 1669390400
transform 1 0 60816 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_557
timestamp 1669390400
transform 1 0 63728 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_567
timestamp 1669390400
transform 1 0 64848 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_570
timestamp 1669390400
transform 1 0 65184 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_573
timestamp 1669390400
transform 1 0 65520 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_583
timestamp 1669390400
transform 1 0 66640 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_25_608
timestamp 1669390400
transform 1 0 69440 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_616
timestamp 1669390400
transform 1 0 70336 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_619
timestamp 1669390400
transform 1 0 70672 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_634
timestamp 1669390400
transform 1 0 72352 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_638
timestamp 1669390400
transform 1 0 72800 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_641
timestamp 1669390400
transform 1 0 73136 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_650
timestamp 1669390400
transform 1 0 74144 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_658
timestamp 1669390400
transform 1 0 75040 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_672
timestamp 1669390400
transform 1 0 76608 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_25_676
timestamp 1669390400
transform 1 0 77056 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_684
timestamp 1669390400
transform 1 0 77952 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_2
timestamp 1669390400
transform 1 0 1568 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_17
timestamp 1669390400
transform 1 0 3248 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_25
timestamp 1669390400
transform 1 0 4144 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_29
timestamp 1669390400
transform 1 0 4592 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_33
timestamp 1669390400
transform 1 0 5040 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_26_37
timestamp 1669390400
transform 1 0 5488 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_45
timestamp 1669390400
transform 1 0 6384 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_49
timestamp 1669390400
transform 1 0 6832 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_51
timestamp 1669390400
transform 1 0 7056 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_60
timestamp 1669390400
transform 1 0 8064 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_64
timestamp 1669390400
transform 1 0 8512 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_68
timestamp 1669390400
transform 1 0 8960 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_72
timestamp 1669390400
transform 1 0 9408 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_76
timestamp 1669390400
transform 1 0 9856 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_89
timestamp 1669390400
transform 1 0 11312 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_95
timestamp 1669390400
transform 1 0 11984 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_99
timestamp 1669390400
transform 1 0 12432 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_105
timestamp 1669390400
transform 1 0 13104 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_108
timestamp 1669390400
transform 1 0 13440 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_115
timestamp 1669390400
transform 1 0 14224 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_26_119
timestamp 1669390400
transform 1 0 14672 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_135
timestamp 1669390400
transform 1 0 16464 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_139
timestamp 1669390400
transform 1 0 16912 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_141
timestamp 1669390400
transform 1 0 17136 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_144
timestamp 1669390400
transform 1 0 17472 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_148
timestamp 1669390400
transform 1 0 17920 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_155
timestamp 1669390400
transform 1 0 18704 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_169
timestamp 1669390400
transform 1 0 20272 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_173
timestamp 1669390400
transform 1 0 20720 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_176
timestamp 1669390400
transform 1 0 21056 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_179
timestamp 1669390400
transform 1 0 21392 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_185
timestamp 1669390400
transform 1 0 22064 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_189
timestamp 1669390400
transform 1 0 22512 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_200
timestamp 1669390400
transform 1 0 23744 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_204
timestamp 1669390400
transform 1 0 24192 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_208
timestamp 1669390400
transform 1 0 24640 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_212
timestamp 1669390400
transform 1 0 25088 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_223
timestamp 1669390400
transform 1 0 26320 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_235
timestamp 1669390400
transform 1 0 27664 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_26_239
timestamp 1669390400
transform 1 0 28112 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_247
timestamp 1669390400
transform 1 0 29008 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_250
timestamp 1669390400
transform 1 0 29344 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_254
timestamp 1669390400
transform 1 0 29792 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_256
timestamp 1669390400
transform 1 0 30016 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_26_262
timestamp 1669390400
transform 1 0 30688 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_280
timestamp 1669390400
transform 1 0 32704 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_294
timestamp 1669390400
transform 1 0 34272 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_301
timestamp 1669390400
transform 1 0 35056 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_26_308
timestamp 1669390400
transform 1 0 35840 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_318
timestamp 1669390400
transform 1 0 36960 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_321
timestamp 1669390400
transform 1 0 37296 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_331
timestamp 1669390400
transform 1 0 38416 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_338
timestamp 1669390400
transform 1 0 39200 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_340
timestamp 1669390400
transform 1 0 39424 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_343
timestamp 1669390400
transform 1 0 39760 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_351
timestamp 1669390400
transform 1 0 40656 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_359
timestamp 1669390400
transform 1 0 41552 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_26_369
timestamp 1669390400
transform 1 0 42672 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_389
timestamp 1669390400
transform 1 0 44912 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_26_392
timestamp 1669390400
transform 1 0 45248 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_408
timestamp 1669390400
transform 1 0 47040 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_422
timestamp 1669390400
transform 1 0 48608 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_426
timestamp 1669390400
transform 1 0 49056 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_430
timestamp 1669390400
transform 1 0 49504 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_26_434
timestamp 1669390400
transform 1 0 49952 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_442
timestamp 1669390400
transform 1 0 50848 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_26_445
timestamp 1669390400
transform 1 0 51184 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_453
timestamp 1669390400
transform 1 0 52080 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_460
timestamp 1669390400
transform 1 0 52864 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_463
timestamp 1669390400
transform 1 0 53200 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_26_472
timestamp 1669390400
transform 1 0 54208 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_488
timestamp 1669390400
transform 1 0 56000 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_492
timestamp 1669390400
transform 1 0 56448 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_494
timestamp 1669390400
transform 1 0 56672 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_497
timestamp 1669390400
transform 1 0 57008 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_511
timestamp 1669390400
transform 1 0 58576 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_518
timestamp 1669390400
transform 1 0 59360 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_525
timestamp 1669390400
transform 1 0 60144 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_529
timestamp 1669390400
transform 1 0 60592 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_531
timestamp 1669390400
transform 1 0 60816 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_534
timestamp 1669390400
transform 1 0 61152 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_26_543
timestamp 1669390400
transform 1 0 62160 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_559
timestamp 1669390400
transform 1 0 63952 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_563
timestamp 1669390400
transform 1 0 64400 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_565
timestamp 1669390400
transform 1 0 64624 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_568
timestamp 1669390400
transform 1 0 64960 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_575
timestamp 1669390400
transform 1 0 65744 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_584
timestamp 1669390400
transform 1 0 66752 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_588
timestamp 1669390400
transform 1 0 67200 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_592
timestamp 1669390400
transform 1 0 67648 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_596
timestamp 1669390400
transform 1 0 68096 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_600
timestamp 1669390400
transform 1 0 68544 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_602
timestamp 1669390400
transform 1 0 68768 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_26_605
timestamp 1669390400
transform 1 0 69104 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_621
timestamp 1669390400
transform 1 0 70896 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_625
timestamp 1669390400
transform 1 0 71344 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_26_638
timestamp 1669390400
transform 1 0 72800 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_654
timestamp 1669390400
transform 1 0 74592 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_670
timestamp 1669390400
transform 1 0 76384 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_676
timestamp 1669390400
transform 1 0 77056 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_26_679
timestamp 1669390400
transform 1 0 77392 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_687
timestamp 1669390400
transform 1 0 78288 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_2
timestamp 1669390400
transform 1 0 1568 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_6
timestamp 1669390400
transform 1 0 2016 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_8
timestamp 1669390400
transform 1 0 2240 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_22
timestamp 1669390400
transform 1 0 3808 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_29
timestamp 1669390400
transform 1 0 4592 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_27_33
timestamp 1669390400
transform 1 0 5040 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_41
timestamp 1669390400
transform 1 0 5936 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_43
timestamp 1669390400
transform 1 0 6160 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_56
timestamp 1669390400
transform 1 0 7616 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_64
timestamp 1669390400
transform 1 0 8512 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_70
timestamp 1669390400
transform 1 0 9184 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_73
timestamp 1669390400
transform 1 0 9520 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_79
timestamp 1669390400
transform 1 0 10192 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_86
timestamp 1669390400
transform 1 0 10976 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_93
timestamp 1669390400
transform 1 0 11760 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_97
timestamp 1669390400
transform 1 0 12208 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_99
timestamp 1669390400
transform 1 0 12432 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_112
timestamp 1669390400
transform 1 0 13888 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_126
timestamp 1669390400
transform 1 0 15456 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_136
timestamp 1669390400
transform 1 0 16576 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_140
timestamp 1669390400
transform 1 0 17024 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_144
timestamp 1669390400
transform 1 0 17472 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_148
timestamp 1669390400
transform 1 0 17920 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_150
timestamp 1669390400
transform 1 0 18144 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_175
timestamp 1669390400
transform 1 0 20944 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_179
timestamp 1669390400
transform 1 0 21392 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_182
timestamp 1669390400
transform 1 0 21728 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_186
timestamp 1669390400
transform 1 0 22176 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_197
timestamp 1669390400
transform 1 0 23408 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_201
timestamp 1669390400
transform 1 0 23856 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_204
timestamp 1669390400
transform 1 0 24192 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_208
timestamp 1669390400
transform 1 0 24640 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_212
timestamp 1669390400
transform 1 0 25088 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_215
timestamp 1669390400
transform 1 0 25424 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_218
timestamp 1669390400
transform 1 0 25760 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_229
timestamp 1669390400
transform 1 0 26992 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_231
timestamp 1669390400
transform 1 0 27216 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_238
timestamp 1669390400
transform 1 0 28000 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_27_242
timestamp 1669390400
transform 1 0 28448 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_250
timestamp 1669390400
transform 1 0 29344 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_27_266
timestamp 1669390400
transform 1 0 31136 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_274
timestamp 1669390400
transform 1 0 32032 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_283
timestamp 1669390400
transform 1 0 33040 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_286
timestamp 1669390400
transform 1 0 33376 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_300
timestamp 1669390400
transform 1 0 34944 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_27_307
timestamp 1669390400
transform 1 0 35728 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_327
timestamp 1669390400
transform 1 0 37968 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_27_342
timestamp 1669390400
transform 1 0 39648 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_350
timestamp 1669390400
transform 1 0 40544 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_354
timestamp 1669390400
transform 1 0 40992 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_27_357
timestamp 1669390400
transform 1 0 41328 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_378
timestamp 1669390400
transform 1 0 43680 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_387
timestamp 1669390400
transform 1 0 44688 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_391
timestamp 1669390400
transform 1 0 45136 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_395
timestamp 1669390400
transform 1 0 45584 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_399
timestamp 1669390400
transform 1 0 46032 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_401
timestamp 1669390400
transform 1 0 46256 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_425
timestamp 1669390400
transform 1 0 48944 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_27_428
timestamp 1669390400
transform 1 0 49280 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_27_444
timestamp 1669390400
transform 1 0 51072 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_452
timestamp 1669390400
transform 1 0 51968 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_466
timestamp 1669390400
transform 1 0 53536 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_27_480
timestamp 1669390400
transform 1 0 55104 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_496
timestamp 1669390400
transform 1 0 56896 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_499
timestamp 1669390400
transform 1 0 57232 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_513
timestamp 1669390400
transform 1 0 58800 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_520
timestamp 1669390400
transform 1 0 59584 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_524
timestamp 1669390400
transform 1 0 60032 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_528
timestamp 1669390400
transform 1 0 60480 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_532
timestamp 1669390400
transform 1 0 60928 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_547
timestamp 1669390400
transform 1 0 62608 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_551
timestamp 1669390400
transform 1 0 63056 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_553
timestamp 1669390400
transform 1 0 63280 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_556
timestamp 1669390400
transform 1 0 63616 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_560
timestamp 1669390400
transform 1 0 64064 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_567
timestamp 1669390400
transform 1 0 64848 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_570
timestamp 1669390400
transform 1 0 65184 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_576
timestamp 1669390400
transform 1 0 65856 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_580
timestamp 1669390400
transform 1 0 66304 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_587
timestamp 1669390400
transform 1 0 67088 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_591
timestamp 1669390400
transform 1 0 67536 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_27_595
timestamp 1669390400
transform 1 0 67984 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_603
timestamp 1669390400
transform 1 0 68880 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_606
timestamp 1669390400
transform 1 0 69216 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_610
timestamp 1669390400
transform 1 0 69664 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_613
timestamp 1669390400
transform 1 0 70000 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_627
timestamp 1669390400
transform 1 0 71568 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_634
timestamp 1669390400
transform 1 0 72352 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_638
timestamp 1669390400
transform 1 0 72800 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_641
timestamp 1669390400
transform 1 0 73136 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_647
timestamp 1669390400
transform 1 0 73808 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_651
timestamp 1669390400
transform 1 0 74256 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_655
timestamp 1669390400
transform 1 0 74704 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_662
timestamp 1669390400
transform 1 0 75488 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_676
timestamp 1669390400
transform 1 0 77056 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_683
timestamp 1669390400
transform 1 0 77840 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_687
timestamp 1669390400
transform 1 0 78288 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_28_2
timestamp 1669390400
transform 1 0 1568 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_23
timestamp 1669390400
transform 1 0 3920 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_31
timestamp 1669390400
transform 1 0 4816 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_37
timestamp 1669390400
transform 1 0 5488 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_53
timestamp 1669390400
transform 1 0 7280 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_61
timestamp 1669390400
transform 1 0 8176 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_63
timestamp 1669390400
transform 1 0 8400 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_66
timestamp 1669390400
transform 1 0 8736 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_72
timestamp 1669390400
transform 1 0 9408 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_76
timestamp 1669390400
transform 1 0 9856 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_90
timestamp 1669390400
transform 1 0 11424 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_94
timestamp 1669390400
transform 1 0 11872 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_98
timestamp 1669390400
transform 1 0 12320 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_102
timestamp 1669390400
transform 1 0 12768 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_28_108
timestamp 1669390400
transform 1 0 13440 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_116
timestamp 1669390400
transform 1 0 14336 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_120
timestamp 1669390400
transform 1 0 14784 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_28_124
timestamp 1669390400
transform 1 0 15232 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_140
timestamp 1669390400
transform 1 0 17024 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_142
timestamp 1669390400
transform 1 0 17248 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_145
timestamp 1669390400
transform 1 0 17584 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_166
timestamp 1669390400
transform 1 0 19936 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_173
timestamp 1669390400
transform 1 0 20720 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_179
timestamp 1669390400
transform 1 0 21392 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_189
timestamp 1669390400
transform 1 0 22512 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_191
timestamp 1669390400
transform 1 0 22736 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_194
timestamp 1669390400
transform 1 0 23072 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_204
timestamp 1669390400
transform 1 0 24192 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_212
timestamp 1669390400
transform 1 0 25088 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_216
timestamp 1669390400
transform 1 0 25536 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_219
timestamp 1669390400
transform 1 0 25872 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_223
timestamp 1669390400
transform 1 0 26320 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_230
timestamp 1669390400
transform 1 0 27104 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_242
timestamp 1669390400
transform 1 0 28448 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_246
timestamp 1669390400
transform 1 0 28896 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_28_250
timestamp 1669390400
transform 1 0 29344 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_28_266
timestamp 1669390400
transform 1 0 31136 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_274
timestamp 1669390400
transform 1 0 32032 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_278
timestamp 1669390400
transform 1 0 32480 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_280
timestamp 1669390400
transform 1 0 32704 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_286
timestamp 1669390400
transform 1 0 33376 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_28_300
timestamp 1669390400
transform 1 0 34944 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_316
timestamp 1669390400
transform 1 0 36736 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_318
timestamp 1669390400
transform 1 0 36960 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_321
timestamp 1669390400
transform 1 0 37296 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_325
timestamp 1669390400
transform 1 0 37744 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_329
timestamp 1669390400
transform 1 0 38192 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_335
timestamp 1669390400
transform 1 0 38864 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_339
timestamp 1669390400
transform 1 0 39312 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_350
timestamp 1669390400
transform 1 0 40544 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_354
timestamp 1669390400
transform 1 0 40992 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_28_358
timestamp 1669390400
transform 1 0 41440 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_386
timestamp 1669390400
transform 1 0 44576 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_392
timestamp 1669390400
transform 1 0 45248 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_28_398
timestamp 1669390400
transform 1 0 45920 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_28_430
timestamp 1669390400
transform 1 0 49504 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_28_446
timestamp 1669390400
transform 1 0 51296 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_454
timestamp 1669390400
transform 1 0 52192 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_458
timestamp 1669390400
transform 1 0 52640 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_460
timestamp 1669390400
transform 1 0 52864 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_463
timestamp 1669390400
transform 1 0 53200 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_28_476
timestamp 1669390400
transform 1 0 54656 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_494
timestamp 1669390400
transform 1 0 56672 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_501
timestamp 1669390400
transform 1 0 57456 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_513
timestamp 1669390400
transform 1 0 58800 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_517
timestamp 1669390400
transform 1 0 59248 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_521
timestamp 1669390400
transform 1 0 59696 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_525
timestamp 1669390400
transform 1 0 60144 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_529
timestamp 1669390400
transform 1 0 60592 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_531
timestamp 1669390400
transform 1 0 60816 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_534
timestamp 1669390400
transform 1 0 61152 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_537
timestamp 1669390400
transform 1 0 61488 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_541
timestamp 1669390400
transform 1 0 61936 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_551
timestamp 1669390400
transform 1 0 63056 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_555
timestamp 1669390400
transform 1 0 63504 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_559
timestamp 1669390400
transform 1 0 63952 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_563
timestamp 1669390400
transform 1 0 64400 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_567
timestamp 1669390400
transform 1 0 64848 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_571
timestamp 1669390400
transform 1 0 65296 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_573
timestamp 1669390400
transform 1 0 65520 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_587
timestamp 1669390400
transform 1 0 67088 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_602
timestamp 1669390400
transform 1 0 68768 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_605
timestamp 1669390400
transform 1 0 69104 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_28_614
timestamp 1669390400
transform 1 0 70112 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_630
timestamp 1669390400
transform 1 0 71904 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_28_637
timestamp 1669390400
transform 1 0 72688 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_28_653
timestamp 1669390400
transform 1 0 74480 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_673
timestamp 1669390400
transform 1 0 76720 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_676
timestamp 1669390400
transform 1 0 77056 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_681
timestamp 1669390400
transform 1 0 77616 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_685
timestamp 1669390400
transform 1 0 78064 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_687
timestamp 1669390400
transform 1 0 78288 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_2
timestamp 1669390400
transform 1 0 1568 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_17
timestamp 1669390400
transform 1 0 3248 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_29
timestamp 1669390400
transform 1 0 4592 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_39
timestamp 1669390400
transform 1 0 5712 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_49
timestamp 1669390400
transform 1 0 6832 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_51
timestamp 1669390400
transform 1 0 7056 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_57
timestamp 1669390400
transform 1 0 7728 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_61
timestamp 1669390400
transform 1 0 8176 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_70
timestamp 1669390400
transform 1 0 9184 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_73
timestamp 1669390400
transform 1 0 9520 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_76
timestamp 1669390400
transform 1 0 9856 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_78
timestamp 1669390400
transform 1 0 10080 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_87
timestamp 1669390400
transform 1 0 11088 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_89
timestamp 1669390400
transform 1 0 11312 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_97
timestamp 1669390400
transform 1 0 12208 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_101
timestamp 1669390400
transform 1 0 12656 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_105
timestamp 1669390400
transform 1 0 13104 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_116
timestamp 1669390400
transform 1 0 14336 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_126
timestamp 1669390400
transform 1 0 15456 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_130
timestamp 1669390400
transform 1 0 15904 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_134
timestamp 1669390400
transform 1 0 16352 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_141
timestamp 1669390400
transform 1 0 17136 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_144
timestamp 1669390400
transform 1 0 17472 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_168
timestamp 1669390400
transform 1 0 20160 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_175
timestamp 1669390400
transform 1 0 20944 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_179
timestamp 1669390400
transform 1 0 21392 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_182
timestamp 1669390400
transform 1 0 21728 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_186
timestamp 1669390400
transform 1 0 22176 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_190
timestamp 1669390400
transform 1 0 22624 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_200
timestamp 1669390400
transform 1 0 23744 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_202
timestamp 1669390400
transform 1 0 23968 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_205
timestamp 1669390400
transform 1 0 24304 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_209
timestamp 1669390400
transform 1 0 24752 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_215
timestamp 1669390400
transform 1 0 25424 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_29_218
timestamp 1669390400
transform 1 0 25760 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_226
timestamp 1669390400
transform 1 0 26656 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_230
timestamp 1669390400
transform 1 0 27104 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_29_243
timestamp 1669390400
transform 1 0 28560 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_251
timestamp 1669390400
transform 1 0 29456 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_256
timestamp 1669390400
transform 1 0 30016 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_270
timestamp 1669390400
transform 1 0 31584 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_280
timestamp 1669390400
transform 1 0 32704 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_286
timestamp 1669390400
transform 1 0 33376 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_292
timestamp 1669390400
transform 1 0 34048 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_306
timestamp 1669390400
transform 1 0 35616 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_29_316
timestamp 1669390400
transform 1 0 36736 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_324
timestamp 1669390400
transform 1 0 37632 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_328
timestamp 1669390400
transform 1 0 38080 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_335
timestamp 1669390400
transform 1 0 38864 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_350
timestamp 1669390400
transform 1 0 40544 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_354
timestamp 1669390400
transform 1 0 40992 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_357
timestamp 1669390400
transform 1 0 41328 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_366
timestamp 1669390400
transform 1 0 42336 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_370
timestamp 1669390400
transform 1 0 42784 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_372
timestamp 1669390400
transform 1 0 43008 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_375
timestamp 1669390400
transform 1 0 43344 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_382
timestamp 1669390400
transform 1 0 44128 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_392
timestamp 1669390400
transform 1 0 45248 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_29_396
timestamp 1669390400
transform 1 0 45696 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_412
timestamp 1669390400
transform 1 0 47488 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_416
timestamp 1669390400
transform 1 0 47936 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_425
timestamp 1669390400
transform 1 0 48944 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_428
timestamp 1669390400
transform 1 0 49280 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_435
timestamp 1669390400
transform 1 0 50064 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_29_443
timestamp 1669390400
transform 1 0 50960 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_451
timestamp 1669390400
transform 1 0 51856 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_455
timestamp 1669390400
transform 1 0 52304 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_29_469
timestamp 1669390400
transform 1 0 53872 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_485
timestamp 1669390400
transform 1 0 55664 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_489
timestamp 1669390400
transform 1 0 56112 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_492
timestamp 1669390400
transform 1 0 56448 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_496
timestamp 1669390400
transform 1 0 56896 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_499
timestamp 1669390400
transform 1 0 57232 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_509
timestamp 1669390400
transform 1 0 58352 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_513
timestamp 1669390400
transform 1 0 58800 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_517
timestamp 1669390400
transform 1 0 59248 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_521
timestamp 1669390400
transform 1 0 59696 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_531
timestamp 1669390400
transform 1 0 60816 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_545
timestamp 1669390400
transform 1 0 62384 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_559
timestamp 1669390400
transform 1 0 63952 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_563
timestamp 1669390400
transform 1 0 64400 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_567
timestamp 1669390400
transform 1 0 64848 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_570
timestamp 1669390400
transform 1 0 65184 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_575
timestamp 1669390400
transform 1 0 65744 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_579
timestamp 1669390400
transform 1 0 66192 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_589
timestamp 1669390400
transform 1 0 67312 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_29_597
timestamp 1669390400
transform 1 0 68208 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_613
timestamp 1669390400
transform 1 0 70000 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_619
timestamp 1669390400
transform 1 0 70672 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_623
timestamp 1669390400
transform 1 0 71120 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_638
timestamp 1669390400
transform 1 0 72800 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_641
timestamp 1669390400
transform 1 0 73136 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_645
timestamp 1669390400
transform 1 0 73584 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_654
timestamp 1669390400
transform 1 0 74592 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_670
timestamp 1669390400
transform 1 0 76384 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_685
timestamp 1669390400
transform 1 0 78064 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_687
timestamp 1669390400
transform 1 0 78288 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_30_2
timestamp 1669390400
transform 1 0 1568 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_10
timestamp 1669390400
transform 1 0 2464 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_14
timestamp 1669390400
transform 1 0 2912 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_27
timestamp 1669390400
transform 1 0 4368 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_31
timestamp 1669390400
transform 1 0 4816 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_34
timestamp 1669390400
transform 1 0 5152 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_37
timestamp 1669390400
transform 1 0 5488 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_44
timestamp 1669390400
transform 1 0 6272 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_48
timestamp 1669390400
transform 1 0 6720 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_30_52
timestamp 1669390400
transform 1 0 7168 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_62
timestamp 1669390400
transform 1 0 8288 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_71
timestamp 1669390400
transform 1 0 9296 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_75
timestamp 1669390400
transform 1 0 9744 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_87
timestamp 1669390400
transform 1 0 11088 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_94
timestamp 1669390400
transform 1 0 11872 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_98
timestamp 1669390400
transform 1 0 12320 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_101
timestamp 1669390400
transform 1 0 12656 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_105
timestamp 1669390400
transform 1 0 13104 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_108
timestamp 1669390400
transform 1 0 13440 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_111
timestamp 1669390400
transform 1 0 13776 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_118
timestamp 1669390400
transform 1 0 14560 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_125
timestamp 1669390400
transform 1 0 15344 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_129
timestamp 1669390400
transform 1 0 15792 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_133
timestamp 1669390400
transform 1 0 16240 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_135
timestamp 1669390400
transform 1 0 16464 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_138
timestamp 1669390400
transform 1 0 16800 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_142
timestamp 1669390400
transform 1 0 17248 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_146
timestamp 1669390400
transform 1 0 17696 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_153
timestamp 1669390400
transform 1 0 18480 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_160
timestamp 1669390400
transform 1 0 19264 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_162
timestamp 1669390400
transform 1 0 19488 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_168
timestamp 1669390400
transform 1 0 20160 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_172
timestamp 1669390400
transform 1 0 20608 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_175
timestamp 1669390400
transform 1 0 20944 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_179
timestamp 1669390400
transform 1 0 21392 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_182
timestamp 1669390400
transform 1 0 21728 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_186
timestamp 1669390400
transform 1 0 22176 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_197
timestamp 1669390400
transform 1 0 23408 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_207
timestamp 1669390400
transform 1 0 24528 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_211
timestamp 1669390400
transform 1 0 24976 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_215
timestamp 1669390400
transform 1 0 25424 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_219
timestamp 1669390400
transform 1 0 25872 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_222
timestamp 1669390400
transform 1 0 26208 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_229
timestamp 1669390400
transform 1 0 26992 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_237
timestamp 1669390400
transform 1 0 27888 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_243
timestamp 1669390400
transform 1 0 28560 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_247
timestamp 1669390400
transform 1 0 29008 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_30_250
timestamp 1669390400
transform 1 0 29344 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_258
timestamp 1669390400
transform 1 0 30240 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_262
timestamp 1669390400
transform 1 0 30688 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_266
timestamp 1669390400
transform 1 0 31136 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_275
timestamp 1669390400
transform 1 0 32144 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_30_279
timestamp 1669390400
transform 1 0 32592 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_287
timestamp 1669390400
transform 1 0 33488 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_290
timestamp 1669390400
transform 1 0 33824 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_300
timestamp 1669390400
transform 1 0 34944 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_315
timestamp 1669390400
transform 1 0 36624 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_30_321
timestamp 1669390400
transform 1 0 37296 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_329
timestamp 1669390400
transform 1 0 38192 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_331
timestamp 1669390400
transform 1 0 38416 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_334
timestamp 1669390400
transform 1 0 38752 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_340
timestamp 1669390400
transform 1 0 39424 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_358
timestamp 1669390400
transform 1 0 41440 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_362
timestamp 1669390400
transform 1 0 41888 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_30_366
timestamp 1669390400
transform 1 0 42336 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_374
timestamp 1669390400
transform 1 0 43232 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_376
timestamp 1669390400
transform 1 0 43456 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_389
timestamp 1669390400
transform 1 0 44912 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_392
timestamp 1669390400
transform 1 0 45248 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_30_403
timestamp 1669390400
transform 1 0 46480 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_411
timestamp 1669390400
transform 1 0 47376 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_415
timestamp 1669390400
transform 1 0 47824 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_30_431
timestamp 1669390400
transform 1 0 49616 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_447
timestamp 1669390400
transform 1 0 51408 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_451
timestamp 1669390400
transform 1 0 51856 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_453
timestamp 1669390400
transform 1 0 52080 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_460
timestamp 1669390400
transform 1 0 52864 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_463
timestamp 1669390400
transform 1 0 53200 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_472
timestamp 1669390400
transform 1 0 54208 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_30_480
timestamp 1669390400
transform 1 0 55104 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_494
timestamp 1669390400
transform 1 0 56672 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_504
timestamp 1669390400
transform 1 0 57792 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_30_518
timestamp 1669390400
transform 1 0 59360 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_526
timestamp 1669390400
transform 1 0 60256 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_530
timestamp 1669390400
transform 1 0 60704 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_534
timestamp 1669390400
transform 1 0 61152 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_536
timestamp 1669390400
transform 1 0 61376 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_542
timestamp 1669390400
transform 1 0 62048 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_546
timestamp 1669390400
transform 1 0 62496 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_548
timestamp 1669390400
transform 1 0 62720 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_555
timestamp 1669390400
transform 1 0 63504 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_562
timestamp 1669390400
transform 1 0 64288 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_566
timestamp 1669390400
transform 1 0 64736 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_572
timestamp 1669390400
transform 1 0 65408 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_30_582
timestamp 1669390400
transform 1 0 66528 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_590
timestamp 1669390400
transform 1 0 67424 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_594
timestamp 1669390400
transform 1 0 67872 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_596
timestamp 1669390400
transform 1 0 68096 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_602
timestamp 1669390400
transform 1 0 68768 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_605
timestamp 1669390400
transform 1 0 69104 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_618
timestamp 1669390400
transform 1 0 70560 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_632
timestamp 1669390400
transform 1 0 72128 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_30_642
timestamp 1669390400
transform 1 0 73248 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_652
timestamp 1669390400
transform 1 0 74368 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_660
timestamp 1669390400
transform 1 0 75264 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_672
timestamp 1669390400
transform 1 0 76608 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_676
timestamp 1669390400
transform 1 0 77056 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_683
timestamp 1669390400
transform 1 0 77840 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_687
timestamp 1669390400
transform 1 0 78288 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_2
timestamp 1669390400
transform 1 0 1568 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_6
timestamp 1669390400
transform 1 0 2016 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_8
timestamp 1669390400
transform 1 0 2240 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_32
timestamp 1669390400
transform 1 0 4928 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_42
timestamp 1669390400
transform 1 0 6048 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_49
timestamp 1669390400
transform 1 0 6832 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_53
timestamp 1669390400
transform 1 0 7280 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_55
timestamp 1669390400
transform 1 0 7504 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_68
timestamp 1669390400
transform 1 0 8960 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_70
timestamp 1669390400
transform 1 0 9184 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_73
timestamp 1669390400
transform 1 0 9520 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_77
timestamp 1669390400
transform 1 0 9968 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_92
timestamp 1669390400
transform 1 0 11648 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_96
timestamp 1669390400
transform 1 0 12096 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_100
timestamp 1669390400
transform 1 0 12544 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_103
timestamp 1669390400
transform 1 0 12880 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_110
timestamp 1669390400
transform 1 0 13664 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_117
timestamp 1669390400
transform 1 0 14448 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_124
timestamp 1669390400
transform 1 0 15232 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_128
timestamp 1669390400
transform 1 0 15680 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_132
timestamp 1669390400
transform 1 0 16128 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_134
timestamp 1669390400
transform 1 0 16352 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_137
timestamp 1669390400
transform 1 0 16688 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_141
timestamp 1669390400
transform 1 0 17136 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_144
timestamp 1669390400
transform 1 0 17472 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_153
timestamp 1669390400
transform 1 0 18480 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_161
timestamp 1669390400
transform 1 0 19376 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_165
timestamp 1669390400
transform 1 0 19824 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_169
timestamp 1669390400
transform 1 0 20272 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_173
timestamp 1669390400
transform 1 0 20720 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_177
timestamp 1669390400
transform 1 0 21168 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_181
timestamp 1669390400
transform 1 0 21616 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_185
timestamp 1669390400
transform 1 0 22064 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_194
timestamp 1669390400
transform 1 0 23072 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_202
timestamp 1669390400
transform 1 0 23968 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_206
timestamp 1669390400
transform 1 0 24416 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_212
timestamp 1669390400
transform 1 0 25088 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_215
timestamp 1669390400
transform 1 0 25424 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_218
timestamp 1669390400
transform 1 0 25760 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_222
timestamp 1669390400
transform 1 0 26208 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_240
timestamp 1669390400
transform 1 0 28224 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_250
timestamp 1669390400
transform 1 0 29344 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_254
timestamp 1669390400
transform 1 0 29792 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_258
timestamp 1669390400
transform 1 0 30240 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_265
timestamp 1669390400
transform 1 0 31024 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_280
timestamp 1669390400
transform 1 0 32704 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_31_286
timestamp 1669390400
transform 1 0 33376 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_294
timestamp 1669390400
transform 1 0 34272 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_298
timestamp 1669390400
transform 1 0 34720 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_300
timestamp 1669390400
transform 1 0 34944 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_303
timestamp 1669390400
transform 1 0 35280 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_307
timestamp 1669390400
transform 1 0 35728 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_31_322
timestamp 1669390400
transform 1 0 37408 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_340
timestamp 1669390400
transform 1 0 39424 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_354
timestamp 1669390400
transform 1 0 40992 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_357
timestamp 1669390400
transform 1 0 41328 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_31_366
timestamp 1669390400
transform 1 0 42336 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_382
timestamp 1669390400
transform 1 0 44128 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_396
timestamp 1669390400
transform 1 0 45696 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_31_406
timestamp 1669390400
transform 1 0 46816 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_422
timestamp 1669390400
transform 1 0 48608 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_428
timestamp 1669390400
transform 1 0 49280 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_31_442
timestamp 1669390400
transform 1 0 50848 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_450
timestamp 1669390400
transform 1 0 51744 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_470
timestamp 1669390400
transform 1 0 53984 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_482
timestamp 1669390400
transform 1 0 55328 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_486
timestamp 1669390400
transform 1 0 55776 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_489
timestamp 1669390400
transform 1 0 56112 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_496
timestamp 1669390400
transform 1 0 56896 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_499
timestamp 1669390400
transform 1 0 57232 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_502
timestamp 1669390400
transform 1 0 57568 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_512
timestamp 1669390400
transform 1 0 58688 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_520
timestamp 1669390400
transform 1 0 59584 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_524
timestamp 1669390400
transform 1 0 60032 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_526
timestamp 1669390400
transform 1 0 60256 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_529
timestamp 1669390400
transform 1 0 60592 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_533
timestamp 1669390400
transform 1 0 61040 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_542
timestamp 1669390400
transform 1 0 62048 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_546
timestamp 1669390400
transform 1 0 62496 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_31_552
timestamp 1669390400
transform 1 0 63168 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_570
timestamp 1669390400
transform 1 0 65184 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_31_579
timestamp 1669390400
transform 1 0 66192 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_31_595
timestamp 1669390400
transform 1 0 67984 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_31_615
timestamp 1669390400
transform 1 0 70224 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_629
timestamp 1669390400
transform 1 0 71792 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_633
timestamp 1669390400
transform 1 0 72240 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_637
timestamp 1669390400
transform 1 0 72688 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_31_641
timestamp 1669390400
transform 1 0 73136 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_651
timestamp 1669390400
transform 1 0 74256 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_655
timestamp 1669390400
transform 1 0 74704 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_667
timestamp 1669390400
transform 1 0 76048 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_677
timestamp 1669390400
transform 1 0 77168 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_685
timestamp 1669390400
transform 1 0 78064 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_687
timestamp 1669390400
transform 1 0 78288 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_32_2
timestamp 1669390400
transform 1 0 1568 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_10
timestamp 1669390400
transform 1 0 2464 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_18
timestamp 1669390400
transform 1 0 3360 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_22
timestamp 1669390400
transform 1 0 3808 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_26
timestamp 1669390400
transform 1 0 4256 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_34
timestamp 1669390400
transform 1 0 5152 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_37
timestamp 1669390400
transform 1 0 5488 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_40
timestamp 1669390400
transform 1 0 5824 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_44
timestamp 1669390400
transform 1 0 6272 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_46
timestamp 1669390400
transform 1 0 6496 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_55
timestamp 1669390400
transform 1 0 7504 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_32_59
timestamp 1669390400
transform 1 0 7952 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_75
timestamp 1669390400
transform 1 0 9744 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_90
timestamp 1669390400
transform 1 0 11424 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_94
timestamp 1669390400
transform 1 0 11872 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_98
timestamp 1669390400
transform 1 0 12320 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_102
timestamp 1669390400
transform 1 0 12768 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_108
timestamp 1669390400
transform 1 0 13440 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_112
timestamp 1669390400
transform 1 0 13888 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_122
timestamp 1669390400
transform 1 0 15008 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_32_126
timestamp 1669390400
transform 1 0 15456 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_134
timestamp 1669390400
transform 1 0 16352 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_140
timestamp 1669390400
transform 1 0 17024 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_150
timestamp 1669390400
transform 1 0 18144 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_176
timestamp 1669390400
transform 1 0 21056 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_32_179
timestamp 1669390400
transform 1 0 21392 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_189
timestamp 1669390400
transform 1 0 22512 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_195
timestamp 1669390400
transform 1 0 23184 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_199
timestamp 1669390400
transform 1 0 23632 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_214
timestamp 1669390400
transform 1 0 25312 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_221
timestamp 1669390400
transform 1 0 26096 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_223
timestamp 1669390400
transform 1 0 26320 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_231
timestamp 1669390400
transform 1 0 27216 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_238
timestamp 1669390400
transform 1 0 28000 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_240
timestamp 1669390400
transform 1 0 28224 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_247
timestamp 1669390400
transform 1 0 29008 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_250
timestamp 1669390400
transform 1 0 29344 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_263
timestamp 1669390400
transform 1 0 30800 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_267
timestamp 1669390400
transform 1 0 31248 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_271
timestamp 1669390400
transform 1 0 31696 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_285
timestamp 1669390400
transform 1 0 33264 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_292
timestamp 1669390400
transform 1 0 34048 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_32_296
timestamp 1669390400
transform 1 0 34496 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_304
timestamp 1669390400
transform 1 0 35392 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_307
timestamp 1669390400
transform 1 0 35728 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_311
timestamp 1669390400
transform 1 0 36176 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_318
timestamp 1669390400
transform 1 0 36960 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_321
timestamp 1669390400
transform 1 0 37296 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_32_330
timestamp 1669390400
transform 1 0 38304 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_338
timestamp 1669390400
transform 1 0 39200 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_342
timestamp 1669390400
transform 1 0 39648 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_344
timestamp 1669390400
transform 1 0 39872 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_347
timestamp 1669390400
transform 1 0 40208 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_32_357
timestamp 1669390400
transform 1 0 41328 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_389
timestamp 1669390400
transform 1 0 44912 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_32_392
timestamp 1669390400
transform 1 0 45248 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_412
timestamp 1669390400
transform 1 0 47488 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_416
timestamp 1669390400
transform 1 0 47936 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_32_423
timestamp 1669390400
transform 1 0 48720 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_431
timestamp 1669390400
transform 1 0 49616 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_32_441
timestamp 1669390400
transform 1 0 50736 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_449
timestamp 1669390400
transform 1 0 51632 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_453
timestamp 1669390400
transform 1 0 52080 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_458
timestamp 1669390400
transform 1 0 52640 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_460
timestamp 1669390400
transform 1 0 52864 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_463
timestamp 1669390400
transform 1 0 53200 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_471
timestamp 1669390400
transform 1 0 54096 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_479
timestamp 1669390400
transform 1 0 54992 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_486
timestamp 1669390400
transform 1 0 55776 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_32_490
timestamp 1669390400
transform 1 0 56224 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_511
timestamp 1669390400
transform 1 0 58576 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_515
timestamp 1669390400
transform 1 0 59024 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_531
timestamp 1669390400
transform 1 0 60816 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_534
timestamp 1669390400
transform 1 0 61152 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_32_543
timestamp 1669390400
transform 1 0 62160 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_571
timestamp 1669390400
transform 1 0 65296 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_585
timestamp 1669390400
transform 1 0 66864 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_599
timestamp 1669390400
transform 1 0 68432 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_605
timestamp 1669390400
transform 1 0 69104 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_32_611
timestamp 1669390400
transform 1 0 69776 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_32_632
timestamp 1669390400
transform 1 0 72128 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_640
timestamp 1669390400
transform 1 0 73024 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_644
timestamp 1669390400
transform 1 0 73472 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_658
timestamp 1669390400
transform 1 0 75040 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_673
timestamp 1669390400
transform 1 0 76720 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_676
timestamp 1669390400
transform 1 0 77056 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_685
timestamp 1669390400
transform 1 0 78064 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_687
timestamp 1669390400
transform 1 0 78288 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_2
timestamp 1669390400
transform 1 0 1568 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_17
timestamp 1669390400
transform 1 0 3248 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_31
timestamp 1669390400
transform 1 0 4816 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_33_35
timestamp 1669390400
transform 1 0 5264 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_43
timestamp 1669390400
transform 1 0 6160 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_57
timestamp 1669390400
transform 1 0 7728 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_33_61
timestamp 1669390400
transform 1 0 8176 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_69
timestamp 1669390400
transform 1 0 9072 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_73
timestamp 1669390400
transform 1 0 9520 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_75
timestamp 1669390400
transform 1 0 9744 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_78
timestamp 1669390400
transform 1 0 10080 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_80
timestamp 1669390400
transform 1 0 10304 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_94
timestamp 1669390400
transform 1 0 11872 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_101
timestamp 1669390400
transform 1 0 12656 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_105
timestamp 1669390400
transform 1 0 13104 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_109
timestamp 1669390400
transform 1 0 13552 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_111
timestamp 1669390400
transform 1 0 13776 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_114
timestamp 1669390400
transform 1 0 14112 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_128
timestamp 1669390400
transform 1 0 15680 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_132
timestamp 1669390400
transform 1 0 16128 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_136
timestamp 1669390400
transform 1 0 16576 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_140
timestamp 1669390400
transform 1 0 17024 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_144
timestamp 1669390400
transform 1 0 17472 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_148
timestamp 1669390400
transform 1 0 17920 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_154
timestamp 1669390400
transform 1 0 18592 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_33_164
timestamp 1669390400
transform 1 0 19712 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_172
timestamp 1669390400
transform 1 0 20608 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_182
timestamp 1669390400
transform 1 0 21728 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_196
timestamp 1669390400
transform 1 0 23296 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_204
timestamp 1669390400
transform 1 0 24192 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_208
timestamp 1669390400
transform 1 0 24640 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_212
timestamp 1669390400
transform 1 0 25088 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_215
timestamp 1669390400
transform 1 0 25424 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_217
timestamp 1669390400
transform 1 0 25648 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_220
timestamp 1669390400
transform 1 0 25984 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_224
timestamp 1669390400
transform 1 0 26432 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_226
timestamp 1669390400
transform 1 0 26656 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_239
timestamp 1669390400
transform 1 0 28112 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_246
timestamp 1669390400
transform 1 0 28896 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_252
timestamp 1669390400
transform 1 0 29568 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_33_256
timestamp 1669390400
transform 1 0 30016 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_264
timestamp 1669390400
transform 1 0 30912 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_268
timestamp 1669390400
transform 1 0 31360 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_283
timestamp 1669390400
transform 1 0 33040 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_286
timestamp 1669390400
transform 1 0 33376 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_33_292
timestamp 1669390400
transform 1 0 34048 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_308
timestamp 1669390400
transform 1 0 35840 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_312
timestamp 1669390400
transform 1 0 36288 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_328
timestamp 1669390400
transform 1 0 38080 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_334
timestamp 1669390400
transform 1 0 38752 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_344
timestamp 1669390400
transform 1 0 39872 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_354
timestamp 1669390400
transform 1 0 40992 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_357
timestamp 1669390400
transform 1 0 41328 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_382
timestamp 1669390400
transform 1 0 44128 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_386
timestamp 1669390400
transform 1 0 44576 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_400
timestamp 1669390400
transform 1 0 46144 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_33_408
timestamp 1669390400
transform 1 0 47040 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_416
timestamp 1669390400
transform 1 0 47936 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_425
timestamp 1669390400
transform 1 0 48944 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_428
timestamp 1669390400
transform 1 0 49280 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_442
timestamp 1669390400
transform 1 0 50848 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_33_449
timestamp 1669390400
transform 1 0 51632 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_457
timestamp 1669390400
transform 1 0 52528 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_33_464
timestamp 1669390400
transform 1 0 53312 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_472
timestamp 1669390400
transform 1 0 54208 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_481
timestamp 1669390400
transform 1 0 55216 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_496
timestamp 1669390400
transform 1 0 56896 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_499
timestamp 1669390400
transform 1 0 57232 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_503
timestamp 1669390400
transform 1 0 57680 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_517
timestamp 1669390400
transform 1 0 59248 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_524
timestamp 1669390400
transform 1 0 60032 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_528
timestamp 1669390400
transform 1 0 60480 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_33_532
timestamp 1669390400
transform 1 0 60928 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_33_548
timestamp 1669390400
transform 1 0 62720 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_561
timestamp 1669390400
transform 1 0 64176 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_567
timestamp 1669390400
transform 1 0 64848 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_33_570
timestamp 1669390400
transform 1 0 65184 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_586
timestamp 1669390400
transform 1 0 66976 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_588
timestamp 1669390400
transform 1 0 67200 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_591
timestamp 1669390400
transform 1 0 67536 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_595
timestamp 1669390400
transform 1 0 67984 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_599
timestamp 1669390400
transform 1 0 68432 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_601
timestamp 1669390400
transform 1 0 68656 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_33_604
timestamp 1669390400
transform 1 0 68992 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_612
timestamp 1669390400
transform 1 0 69888 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_615
timestamp 1669390400
transform 1 0 70224 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_622
timestamp 1669390400
transform 1 0 71008 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_629
timestamp 1669390400
transform 1 0 71792 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_633
timestamp 1669390400
transform 1 0 72240 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_637
timestamp 1669390400
transform 1 0 72688 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_33_641
timestamp 1669390400
transform 1 0 73136 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_649
timestamp 1669390400
transform 1 0 74032 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_653
timestamp 1669390400
transform 1 0 74480 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_655
timestamp 1669390400
transform 1 0 74704 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_670
timestamp 1669390400
transform 1 0 76384 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_674
timestamp 1669390400
transform 1 0 76832 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_678
timestamp 1669390400
transform 1 0 77280 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_682
timestamp 1669390400
transform 1 0 77728 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_686
timestamp 1669390400
transform 1 0 78176 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_2
timestamp 1669390400
transform 1 0 1568 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_6
timestamp 1669390400
transform 1 0 2016 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_10
timestamp 1669390400
transform 1 0 2464 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_18
timestamp 1669390400
transform 1 0 3360 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_22
timestamp 1669390400
transform 1 0 3808 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_28
timestamp 1669390400
transform 1 0 4480 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_32
timestamp 1669390400
transform 1 0 4928 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_34
timestamp 1669390400
transform 1 0 5152 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_34_37
timestamp 1669390400
transform 1 0 5488 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_45
timestamp 1669390400
transform 1 0 6384 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_34_58
timestamp 1669390400
transform 1 0 7840 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_66
timestamp 1669390400
transform 1 0 8736 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_70
timestamp 1669390400
transform 1 0 9184 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_76
timestamp 1669390400
transform 1 0 9856 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_78
timestamp 1669390400
transform 1 0 10080 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_87
timestamp 1669390400
transform 1 0 11088 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_101
timestamp 1669390400
transform 1 0 12656 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_105
timestamp 1669390400
transform 1 0 13104 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_108
timestamp 1669390400
transform 1 0 13440 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_117
timestamp 1669390400
transform 1 0 14448 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_127
timestamp 1669390400
transform 1 0 15568 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_134
timestamp 1669390400
transform 1 0 16352 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_138
timestamp 1669390400
transform 1 0 16800 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_140
timestamp 1669390400
transform 1 0 17024 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_34_143
timestamp 1669390400
transform 1 0 17360 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_151
timestamp 1669390400
transform 1 0 18256 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_34_166
timestamp 1669390400
transform 1 0 19936 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_174
timestamp 1669390400
transform 1 0 20832 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_176
timestamp 1669390400
transform 1 0 21056 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_34_179
timestamp 1669390400
transform 1 0 21392 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_187
timestamp 1669390400
transform 1 0 22288 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_191
timestamp 1669390400
transform 1 0 22736 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_195
timestamp 1669390400
transform 1 0 23184 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_205
timestamp 1669390400
transform 1 0 24304 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_211
timestamp 1669390400
transform 1 0 24976 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_215
timestamp 1669390400
transform 1 0 25424 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_225
timestamp 1669390400
transform 1 0 26544 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_229
timestamp 1669390400
transform 1 0 26992 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_233
timestamp 1669390400
transform 1 0 27440 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_237
timestamp 1669390400
transform 1 0 27888 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_240
timestamp 1669390400
transform 1 0 28224 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_244
timestamp 1669390400
transform 1 0 28672 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_247
timestamp 1669390400
transform 1 0 29008 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_250
timestamp 1669390400
transform 1 0 29344 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_266
timestamp 1669390400
transform 1 0 31136 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_273
timestamp 1669390400
transform 1 0 31920 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_277
timestamp 1669390400
transform 1 0 32368 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_284
timestamp 1669390400
transform 1 0 33152 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_288
timestamp 1669390400
transform 1 0 33600 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_292
timestamp 1669390400
transform 1 0 34048 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_300
timestamp 1669390400
transform 1 0 34944 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_310
timestamp 1669390400
transform 1 0 36064 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_317
timestamp 1669390400
transform 1 0 36848 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_321
timestamp 1669390400
transform 1 0 37296 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_34_324
timestamp 1669390400
transform 1 0 37632 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_358
timestamp 1669390400
transform 1 0 41440 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_34_362
timestamp 1669390400
transform 1 0 41888 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_378
timestamp 1669390400
transform 1 0 43680 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_381
timestamp 1669390400
transform 1 0 44016 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_389
timestamp 1669390400
transform 1 0 44912 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_392
timestamp 1669390400
transform 1 0 45248 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_396
timestamp 1669390400
transform 1 0 45696 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_411
timestamp 1669390400
transform 1 0 47376 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_417
timestamp 1669390400
transform 1 0 48048 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_34_421
timestamp 1669390400
transform 1 0 48496 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_429
timestamp 1669390400
transform 1 0 49392 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_34_443
timestamp 1669390400
transform 1 0 50960 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_459
timestamp 1669390400
transform 1 0 52752 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_463
timestamp 1669390400
transform 1 0 53200 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_466
timestamp 1669390400
transform 1 0 53536 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_473
timestamp 1669390400
transform 1 0 54320 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_480
timestamp 1669390400
transform 1 0 55104 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_487
timestamp 1669390400
transform 1 0 55888 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_491
timestamp 1669390400
transform 1 0 56336 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_495
timestamp 1669390400
transform 1 0 56784 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_503
timestamp 1669390400
transform 1 0 57680 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_505
timestamp 1669390400
transform 1 0 57904 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_34_512
timestamp 1669390400
transform 1 0 58688 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_528
timestamp 1669390400
transform 1 0 60480 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_531
timestamp 1669390400
transform 1 0 60816 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_534
timestamp 1669390400
transform 1 0 61152 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_34_547
timestamp 1669390400
transform 1 0 62608 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_34_563
timestamp 1669390400
transform 1 0 64400 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_571
timestamp 1669390400
transform 1 0 65296 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_575
timestamp 1669390400
transform 1 0 65744 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_589
timestamp 1669390400
transform 1 0 67312 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_596
timestamp 1669390400
transform 1 0 68096 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_602
timestamp 1669390400
transform 1 0 68768 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_605
timestamp 1669390400
transform 1 0 69104 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_616
timestamp 1669390400
transform 1 0 70336 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_624
timestamp 1669390400
transform 1 0 71232 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_626
timestamp 1669390400
transform 1 0 71456 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_635
timestamp 1669390400
transform 1 0 72464 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_34_639
timestamp 1669390400
transform 1 0 72912 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_647
timestamp 1669390400
transform 1 0 73808 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_655
timestamp 1669390400
transform 1 0 74704 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_669
timestamp 1669390400
transform 1 0 76272 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_673
timestamp 1669390400
transform 1 0 76720 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_676
timestamp 1669390400
transform 1 0 77056 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_685
timestamp 1669390400
transform 1 0 78064 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_687
timestamp 1669390400
transform 1 0 78288 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_35_2
timestamp 1669390400
transform 1 0 1568 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_10
timestamp 1669390400
transform 1 0 2464 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_17
timestamp 1669390400
transform 1 0 3248 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_43
timestamp 1669390400
transform 1 0 6160 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_53
timestamp 1669390400
transform 1 0 7280 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_57
timestamp 1669390400
transform 1 0 7728 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_59
timestamp 1669390400
transform 1 0 7952 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_62
timestamp 1669390400
transform 1 0 8288 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_70
timestamp 1669390400
transform 1 0 9184 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_73
timestamp 1669390400
transform 1 0 9520 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_35_89
timestamp 1669390400
transform 1 0 11312 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_105
timestamp 1669390400
transform 1 0 13104 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_107
timestamp 1669390400
transform 1 0 13328 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_113
timestamp 1669390400
transform 1 0 14000 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_117
timestamp 1669390400
transform 1 0 14448 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_126
timestamp 1669390400
transform 1 0 15456 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_141
timestamp 1669390400
transform 1 0 17136 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_144
timestamp 1669390400
transform 1 0 17472 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_147
timestamp 1669390400
transform 1 0 17808 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_151
timestamp 1669390400
transform 1 0 18256 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_160
timestamp 1669390400
transform 1 0 19264 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_35_174
timestamp 1669390400
transform 1 0 20832 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_190
timestamp 1669390400
transform 1 0 22624 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_193
timestamp 1669390400
transform 1 0 22960 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_207
timestamp 1669390400
transform 1 0 24528 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_209
timestamp 1669390400
transform 1 0 24752 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_212
timestamp 1669390400
transform 1 0 25088 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_215
timestamp 1669390400
transform 1 0 25424 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_228
timestamp 1669390400
transform 1 0 26880 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_35_238
timestamp 1669390400
transform 1 0 28000 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_246
timestamp 1669390400
transform 1 0 28896 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_250
timestamp 1669390400
transform 1 0 29344 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_254
timestamp 1669390400
transform 1 0 29792 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_268
timestamp 1669390400
transform 1 0 31360 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_278
timestamp 1669390400
transform 1 0 32480 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_282
timestamp 1669390400
transform 1 0 32928 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_286
timestamp 1669390400
transform 1 0 33376 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_292
timestamp 1669390400
transform 1 0 34048 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_296
timestamp 1669390400
transform 1 0 34496 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_35_321
timestamp 1669390400
transform 1 0 37296 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_329
timestamp 1669390400
transform 1 0 38192 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_333
timestamp 1669390400
transform 1 0 38640 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_335
timestamp 1669390400
transform 1 0 38864 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_344
timestamp 1669390400
transform 1 0 39872 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_354
timestamp 1669390400
transform 1 0 40992 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_357
timestamp 1669390400
transform 1 0 41328 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_35_366
timestamp 1669390400
transform 1 0 42336 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_374
timestamp 1669390400
transform 1 0 43232 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_35_384
timestamp 1669390400
transform 1 0 44352 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_392
timestamp 1669390400
transform 1 0 45248 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_395
timestamp 1669390400
transform 1 0 45584 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_35_405
timestamp 1669390400
transform 1 0 46704 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_413
timestamp 1669390400
transform 1 0 47600 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_417
timestamp 1669390400
transform 1 0 48048 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_425
timestamp 1669390400
transform 1 0 48944 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_35_428
timestamp 1669390400
transform 1 0 49280 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_453
timestamp 1669390400
transform 1 0 52080 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_35_457
timestamp 1669390400
transform 1 0 52528 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_465
timestamp 1669390400
transform 1 0 53424 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_468
timestamp 1669390400
transform 1 0 53760 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_480
timestamp 1669390400
transform 1 0 55104 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_484
timestamp 1669390400
transform 1 0 55552 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_488
timestamp 1669390400
transform 1 0 56000 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_492
timestamp 1669390400
transform 1 0 56448 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_496
timestamp 1669390400
transform 1 0 56896 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_35_499
timestamp 1669390400
transform 1 0 57232 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_507
timestamp 1669390400
transform 1 0 58128 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_514
timestamp 1669390400
transform 1 0 58912 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_518
timestamp 1669390400
transform 1 0 59360 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_520
timestamp 1669390400
transform 1 0 59584 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_523
timestamp 1669390400
transform 1 0 59920 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_527
timestamp 1669390400
transform 1 0 60368 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_535
timestamp 1669390400
transform 1 0 61264 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_556
timestamp 1669390400
transform 1 0 63616 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_35_560
timestamp 1669390400
transform 1 0 64064 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_570
timestamp 1669390400
transform 1 0 65184 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_582
timestamp 1669390400
transform 1 0 66528 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_592
timestamp 1669390400
transform 1 0 67648 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_596
timestamp 1669390400
transform 1 0 68096 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_602
timestamp 1669390400
transform 1 0 68768 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_612
timestamp 1669390400
transform 1 0 69888 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_626
timestamp 1669390400
transform 1 0 71456 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_636
timestamp 1669390400
transform 1 0 72576 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_638
timestamp 1669390400
transform 1 0 72800 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_35_641
timestamp 1669390400
transform 1 0 73136 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_649
timestamp 1669390400
transform 1 0 74032 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_653
timestamp 1669390400
transform 1 0 74480 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_659
timestamp 1669390400
transform 1 0 75152 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_671
timestamp 1669390400
transform 1 0 76496 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_679
timestamp 1669390400
transform 1 0 77392 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_683
timestamp 1669390400
transform 1 0 77840 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_687
timestamp 1669390400
transform 1 0 78288 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_2
timestamp 1669390400
transform 1 0 1568 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_17
timestamp 1669390400
transform 1 0 3248 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_21
timestamp 1669390400
transform 1 0 3696 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_25
timestamp 1669390400
transform 1 0 4144 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_34
timestamp 1669390400
transform 1 0 5152 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_37
timestamp 1669390400
transform 1 0 5488 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_36_46
timestamp 1669390400
transform 1 0 6496 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_62
timestamp 1669390400
transform 1 0 8288 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_66
timestamp 1669390400
transform 1 0 8736 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_92
timestamp 1669390400
transform 1 0 11648 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_36_96
timestamp 1669390400
transform 1 0 12096 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_104
timestamp 1669390400
transform 1 0 12992 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_108
timestamp 1669390400
transform 1 0 13440 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_122
timestamp 1669390400
transform 1 0 15008 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_130
timestamp 1669390400
transform 1 0 15904 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_134
timestamp 1669390400
transform 1 0 16352 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_36_148
timestamp 1669390400
transform 1 0 17920 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_164
timestamp 1669390400
transform 1 0 19712 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_176
timestamp 1669390400
transform 1 0 21056 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_179
timestamp 1669390400
transform 1 0 21392 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_36_192
timestamp 1669390400
transform 1 0 22848 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_200
timestamp 1669390400
transform 1 0 23744 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_204
timestamp 1669390400
transform 1 0 24192 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_211
timestamp 1669390400
transform 1 0 24976 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_36_215
timestamp 1669390400
transform 1 0 25424 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_223
timestamp 1669390400
transform 1 0 26320 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_36_237
timestamp 1669390400
transform 1 0 27888 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_245
timestamp 1669390400
transform 1 0 28784 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_247
timestamp 1669390400
transform 1 0 29008 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_36_250
timestamp 1669390400
transform 1 0 29344 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_258
timestamp 1669390400
transform 1 0 30240 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_262
timestamp 1669390400
transform 1 0 30688 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_277
timestamp 1669390400
transform 1 0 32368 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_281
timestamp 1669390400
transform 1 0 32816 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_36_291
timestamp 1669390400
transform 1 0 33936 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_36_307
timestamp 1669390400
transform 1 0 35728 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_315
timestamp 1669390400
transform 1 0 36624 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_321
timestamp 1669390400
transform 1 0 37296 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_330
timestamp 1669390400
transform 1 0 38304 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_334
timestamp 1669390400
transform 1 0 38752 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_337
timestamp 1669390400
transform 1 0 39088 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_36_363
timestamp 1669390400
transform 1 0 42000 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_383
timestamp 1669390400
transform 1 0 44240 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_387
timestamp 1669390400
transform 1 0 44688 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_389
timestamp 1669390400
transform 1 0 44912 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_392
timestamp 1669390400
transform 1 0 45248 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_396
timestamp 1669390400
transform 1 0 45696 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_398
timestamp 1669390400
transform 1 0 45920 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_408
timestamp 1669390400
transform 1 0 47040 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_415
timestamp 1669390400
transform 1 0 47824 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_36_419
timestamp 1669390400
transform 1 0 48272 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_427
timestamp 1669390400
transform 1 0 49168 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_439
timestamp 1669390400
transform 1 0 50512 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_448
timestamp 1669390400
transform 1 0 51520 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_452
timestamp 1669390400
transform 1 0 51968 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_456
timestamp 1669390400
transform 1 0 52416 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_460
timestamp 1669390400
transform 1 0 52864 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_463
timestamp 1669390400
transform 1 0 53200 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_472
timestamp 1669390400
transform 1 0 54208 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_497
timestamp 1669390400
transform 1 0 57008 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_501
timestamp 1669390400
transform 1 0 57456 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_505
timestamp 1669390400
transform 1 0 57904 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_507
timestamp 1669390400
transform 1 0 58128 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_510
timestamp 1669390400
transform 1 0 58464 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_514
timestamp 1669390400
transform 1 0 58912 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_523
timestamp 1669390400
transform 1 0 59920 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_530
timestamp 1669390400
transform 1 0 60704 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_534
timestamp 1669390400
transform 1 0 61152 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_543
timestamp 1669390400
transform 1 0 62160 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_549
timestamp 1669390400
transform 1 0 62832 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_560
timestamp 1669390400
transform 1 0 64064 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_36_564
timestamp 1669390400
transform 1 0 64512 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_572
timestamp 1669390400
transform 1 0 65408 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_579
timestamp 1669390400
transform 1 0 66192 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_581
timestamp 1669390400
transform 1 0 66416 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_586
timestamp 1669390400
transform 1 0 66976 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_36_590
timestamp 1669390400
transform 1 0 67424 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_598
timestamp 1669390400
transform 1 0 68320 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_602
timestamp 1669390400
transform 1 0 68768 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_605
timestamp 1669390400
transform 1 0 69104 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_607
timestamp 1669390400
transform 1 0 69328 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_626
timestamp 1669390400
transform 1 0 71456 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_628
timestamp 1669390400
transform 1 0 71680 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_36_633
timestamp 1669390400
transform 1 0 72240 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_646
timestamp 1669390400
transform 1 0 73696 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_654
timestamp 1669390400
transform 1 0 74592 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_670
timestamp 1669390400
transform 1 0 76384 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_676
timestamp 1669390400
transform 1 0 77056 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_683
timestamp 1669390400
transform 1 0 77840 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_687
timestamp 1669390400
transform 1 0 78288 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_37_2
timestamp 1669390400
transform 1 0 1568 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_10
timestamp 1669390400
transform 1 0 2464 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_18
timestamp 1669390400
transform 1 0 3360 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_22
timestamp 1669390400
transform 1 0 3808 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_37_32
timestamp 1669390400
transform 1 0 4928 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_48
timestamp 1669390400
transform 1 0 6720 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_57
timestamp 1669390400
transform 1 0 7728 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_65
timestamp 1669390400
transform 1 0 8624 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_67
timestamp 1669390400
transform 1 0 8848 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_70
timestamp 1669390400
transform 1 0 9184 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_37_73
timestamp 1669390400
transform 1 0 9520 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_37_89
timestamp 1669390400
transform 1 0 11312 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_97
timestamp 1669390400
transform 1 0 12208 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_99
timestamp 1669390400
transform 1 0 12432 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_108
timestamp 1669390400
transform 1 0 13440 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_123
timestamp 1669390400
transform 1 0 15120 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_127
timestamp 1669390400
transform 1 0 15568 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_129
timestamp 1669390400
transform 1 0 15792 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_37_132
timestamp 1669390400
transform 1 0 16128 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_140
timestamp 1669390400
transform 1 0 17024 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_144
timestamp 1669390400
transform 1 0 17472 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_150
timestamp 1669390400
transform 1 0 18144 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_37_166
timestamp 1669390400
transform 1 0 19936 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_182
timestamp 1669390400
transform 1 0 21728 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_192
timestamp 1669390400
transform 1 0 22848 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_198
timestamp 1669390400
transform 1 0 23520 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_212
timestamp 1669390400
transform 1 0 25088 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_37_215
timestamp 1669390400
transform 1 0 25424 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_223
timestamp 1669390400
transform 1 0 26320 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_227
timestamp 1669390400
transform 1 0 26768 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_229
timestamp 1669390400
transform 1 0 26992 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_243
timestamp 1669390400
transform 1 0 28560 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_37_253
timestamp 1669390400
transform 1 0 29680 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_261
timestamp 1669390400
transform 1 0 30576 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_265
timestamp 1669390400
transform 1 0 31024 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_37_274
timestamp 1669390400
transform 1 0 32032 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_282
timestamp 1669390400
transform 1 0 32928 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_286
timestamp 1669390400
transform 1 0 33376 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_37_295
timestamp 1669390400
transform 1 0 34384 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_311
timestamp 1669390400
transform 1 0 36176 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_315
timestamp 1669390400
transform 1 0 36624 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_317
timestamp 1669390400
transform 1 0 36848 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_326
timestamp 1669390400
transform 1 0 37856 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_336
timestamp 1669390400
transform 1 0 38976 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_37_340
timestamp 1669390400
transform 1 0 39424 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_348
timestamp 1669390400
transform 1 0 40320 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_352
timestamp 1669390400
transform 1 0 40768 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_354
timestamp 1669390400
transform 1 0 40992 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_357
timestamp 1669390400
transform 1 0 41328 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_361
timestamp 1669390400
transform 1 0 41776 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_363
timestamp 1669390400
transform 1 0 42000 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_37_368
timestamp 1669390400
transform 1 0 42560 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_37_384
timestamp 1669390400
transform 1 0 44352 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_392
timestamp 1669390400
transform 1 0 45248 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_395
timestamp 1669390400
transform 1 0 45584 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_420
timestamp 1669390400
transform 1 0 48384 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_424
timestamp 1669390400
transform 1 0 48832 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_428
timestamp 1669390400
transform 1 0 49280 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_437
timestamp 1669390400
transform 1 0 50288 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_441
timestamp 1669390400
transform 1 0 50736 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_443
timestamp 1669390400
transform 1 0 50960 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_37_456
timestamp 1669390400
transform 1 0 52416 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_464
timestamp 1669390400
transform 1 0 53312 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_470
timestamp 1669390400
transform 1 0 53984 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_480
timestamp 1669390400
transform 1 0 55104 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_489
timestamp 1669390400
transform 1 0 56112 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_493
timestamp 1669390400
transform 1 0 56560 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_499
timestamp 1669390400
transform 1 0 57232 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_508
timestamp 1669390400
transform 1 0 58240 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_515
timestamp 1669390400
transform 1 0 59024 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_519
timestamp 1669390400
transform 1 0 59472 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_523
timestamp 1669390400
transform 1 0 59920 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_529
timestamp 1669390400
transform 1 0 60592 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_545
timestamp 1669390400
transform 1 0 62384 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_549
timestamp 1669390400
transform 1 0 62832 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_37_559
timestamp 1669390400
transform 1 0 63952 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_567
timestamp 1669390400
transform 1 0 64848 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_37_570
timestamp 1669390400
transform 1 0 65184 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_578
timestamp 1669390400
transform 1 0 66080 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_586
timestamp 1669390400
transform 1 0 66976 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_37_593
timestamp 1669390400
transform 1 0 67760 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_601
timestamp 1669390400
transform 1 0 68656 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_605
timestamp 1669390400
transform 1 0 69104 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_607
timestamp 1669390400
transform 1 0 69328 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_614
timestamp 1669390400
transform 1 0 70112 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_37_628
timestamp 1669390400
transform 1 0 71680 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_636
timestamp 1669390400
transform 1 0 72576 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_638
timestamp 1669390400
transform 1 0 72800 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_37_641
timestamp 1669390400
transform 1 0 73136 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_649
timestamp 1669390400
transform 1 0 74032 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_652
timestamp 1669390400
transform 1 0 74368 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_666
timestamp 1669390400
transform 1 0 75936 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_674
timestamp 1669390400
transform 1 0 76832 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_682
timestamp 1669390400
transform 1 0 77728 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_686
timestamp 1669390400
transform 1 0 78176 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_2
timestamp 1669390400
transform 1 0 1568 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_10
timestamp 1669390400
transform 1 0 2464 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_18
timestamp 1669390400
transform 1 0 3360 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_22
timestamp 1669390400
transform 1 0 3808 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_30
timestamp 1669390400
transform 1 0 4704 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_34
timestamp 1669390400
transform 1 0 5152 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_37
timestamp 1669390400
transform 1 0 5488 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_68
timestamp 1669390400
transform 1 0 8960 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_78
timestamp 1669390400
transform 1 0 10080 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_82
timestamp 1669390400
transform 1 0 10528 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_90
timestamp 1669390400
transform 1 0 11424 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_105
timestamp 1669390400
transform 1 0 13104 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_108
timestamp 1669390400
transform 1 0 13440 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_114
timestamp 1669390400
transform 1 0 14112 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_38_118
timestamp 1669390400
transform 1 0 14560 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_134
timestamp 1669390400
transform 1 0 16352 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_144
timestamp 1669390400
transform 1 0 17472 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_158
timestamp 1669390400
transform 1 0 19040 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_168
timestamp 1669390400
transform 1 0 20160 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_172
timestamp 1669390400
transform 1 0 20608 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_176
timestamp 1669390400
transform 1 0 21056 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_179
timestamp 1669390400
transform 1 0 21392 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_185
timestamp 1669390400
transform 1 0 22064 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_189
timestamp 1669390400
transform 1 0 22512 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_193
timestamp 1669390400
transform 1 0 22960 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_38_203
timestamp 1669390400
transform 1 0 24080 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_235
timestamp 1669390400
transform 1 0 27664 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_247
timestamp 1669390400
transform 1 0 29008 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_250
timestamp 1669390400
transform 1 0 29344 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_264
timestamp 1669390400
transform 1 0 30912 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_272
timestamp 1669390400
transform 1 0 31808 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_276
timestamp 1669390400
transform 1 0 32256 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_302
timestamp 1669390400
transform 1 0 35168 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_310
timestamp 1669390400
transform 1 0 36064 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_314
timestamp 1669390400
transform 1 0 36512 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_318
timestamp 1669390400
transform 1 0 36960 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_321
timestamp 1669390400
transform 1 0 37296 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_323
timestamp 1669390400
transform 1 0 37520 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_38_348
timestamp 1669390400
transform 1 0 40320 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_364
timestamp 1669390400
transform 1 0 42112 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_366
timestamp 1669390400
transform 1 0 42336 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_375
timestamp 1669390400
transform 1 0 43344 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_389
timestamp 1669390400
transform 1 0 44912 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_392
timestamp 1669390400
transform 1 0 45248 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_398
timestamp 1669390400
transform 1 0 45920 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_406
timestamp 1669390400
transform 1 0 46816 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_408
timestamp 1669390400
transform 1 0 47040 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_411
timestamp 1669390400
transform 1 0 47376 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_415
timestamp 1669390400
transform 1 0 47824 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_435
timestamp 1669390400
transform 1 0 50064 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_445
timestamp 1669390400
transform 1 0 51184 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_452
timestamp 1669390400
transform 1 0 51968 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_456
timestamp 1669390400
transform 1 0 52416 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_460
timestamp 1669390400
transform 1 0 52864 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_463
timestamp 1669390400
transform 1 0 53200 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_477
timestamp 1669390400
transform 1 0 54768 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_481
timestamp 1669390400
transform 1 0 55216 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_483
timestamp 1669390400
transform 1 0 55440 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_496
timestamp 1669390400
transform 1 0 56896 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_506
timestamp 1669390400
transform 1 0 58016 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_514
timestamp 1669390400
transform 1 0 58912 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_517
timestamp 1669390400
transform 1 0 59248 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_525
timestamp 1669390400
transform 1 0 60144 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_531
timestamp 1669390400
transform 1 0 60816 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_534
timestamp 1669390400
transform 1 0 61152 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_540
timestamp 1669390400
transform 1 0 61824 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_544
timestamp 1669390400
transform 1 0 62272 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_548
timestamp 1669390400
transform 1 0 62720 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_554
timestamp 1669390400
transform 1 0 63392 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_556
timestamp 1669390400
transform 1 0 63616 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_562
timestamp 1669390400
transform 1 0 64288 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_566
timestamp 1669390400
transform 1 0 64736 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_576
timestamp 1669390400
transform 1 0 65856 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_590
timestamp 1669390400
transform 1 0 67424 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_598
timestamp 1669390400
transform 1 0 68320 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_602
timestamp 1669390400
transform 1 0 68768 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_605
timestamp 1669390400
transform 1 0 69104 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_625
timestamp 1669390400
transform 1 0 71344 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_635
timestamp 1669390400
transform 1 0 72464 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_639
timestamp 1669390400
transform 1 0 72912 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_642
timestamp 1669390400
transform 1 0 73248 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_646
timestamp 1669390400
transform 1 0 73696 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_649
timestamp 1669390400
transform 1 0 74032 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_653
timestamp 1669390400
transform 1 0 74480 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_661
timestamp 1669390400
transform 1 0 75376 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_665
timestamp 1669390400
transform 1 0 75824 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_673
timestamp 1669390400
transform 1 0 76720 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_676
timestamp 1669390400
transform 1 0 77056 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_683
timestamp 1669390400
transform 1 0 77840 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_687
timestamp 1669390400
transform 1 0 78288 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_2
timestamp 1669390400
transform 1 0 1568 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_39_17
timestamp 1669390400
transform 1 0 3248 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_33
timestamp 1669390400
transform 1 0 5040 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_41
timestamp 1669390400
transform 1 0 5936 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_45
timestamp 1669390400
transform 1 0 6384 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_70
timestamp 1669390400
transform 1 0 9184 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_73
timestamp 1669390400
transform 1 0 9520 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_39_76
timestamp 1669390400
transform 1 0 9856 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_92
timestamp 1669390400
transform 1 0 11648 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_96
timestamp 1669390400
transform 1 0 12096 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_100
timestamp 1669390400
transform 1 0 12544 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_113
timestamp 1669390400
transform 1 0 14000 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_121
timestamp 1669390400
transform 1 0 14896 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_125
timestamp 1669390400
transform 1 0 15344 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_129
timestamp 1669390400
transform 1 0 15792 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_133
timestamp 1669390400
transform 1 0 16240 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_137
timestamp 1669390400
transform 1 0 16688 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_141
timestamp 1669390400
transform 1 0 17136 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_144
timestamp 1669390400
transform 1 0 17472 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_151
timestamp 1669390400
transform 1 0 18256 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_153
timestamp 1669390400
transform 1 0 18480 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_159
timestamp 1669390400
transform 1 0 19152 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_161
timestamp 1669390400
transform 1 0 19376 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_186
timestamp 1669390400
transform 1 0 22176 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_190
timestamp 1669390400
transform 1 0 22624 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_203
timestamp 1669390400
transform 1 0 24080 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_207
timestamp 1669390400
transform 1 0 24528 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_209
timestamp 1669390400
transform 1 0 24752 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_212
timestamp 1669390400
transform 1 0 25088 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_215
timestamp 1669390400
transform 1 0 25424 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_227
timestamp 1669390400
transform 1 0 26768 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_39_234
timestamp 1669390400
transform 1 0 27552 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_250
timestamp 1669390400
transform 1 0 29344 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_258
timestamp 1669390400
transform 1 0 30240 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_264
timestamp 1669390400
transform 1 0 30912 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_272
timestamp 1669390400
transform 1 0 31808 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_280
timestamp 1669390400
transform 1 0 32704 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_283
timestamp 1669390400
transform 1 0 33040 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_286
timestamp 1669390400
transform 1 0 33376 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_296
timestamp 1669390400
transform 1 0 34496 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_300
timestamp 1669390400
transform 1 0 34944 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_309
timestamp 1669390400
transform 1 0 35952 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_317
timestamp 1669390400
transform 1 0 36848 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_325
timestamp 1669390400
transform 1 0 37744 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_333
timestamp 1669390400
transform 1 0 38640 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_337
timestamp 1669390400
transform 1 0 39088 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_345
timestamp 1669390400
transform 1 0 39984 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_352
timestamp 1669390400
transform 1 0 40768 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_354
timestamp 1669390400
transform 1 0 40992 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_357
timestamp 1669390400
transform 1 0 41328 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_361
timestamp 1669390400
transform 1 0 41776 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_363
timestamp 1669390400
transform 1 0 42000 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_370
timestamp 1669390400
transform 1 0 42784 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_39_382
timestamp 1669390400
transform 1 0 44128 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_414
timestamp 1669390400
transform 1 0 47712 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_422
timestamp 1669390400
transform 1 0 48608 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_428
timestamp 1669390400
transform 1 0 49280 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_432
timestamp 1669390400
transform 1 0 49728 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_446
timestamp 1669390400
transform 1 0 51296 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_453
timestamp 1669390400
transform 1 0 52080 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_460
timestamp 1669390400
transform 1 0 52864 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_464
timestamp 1669390400
transform 1 0 53312 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_466
timestamp 1669390400
transform 1 0 53536 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_472
timestamp 1669390400
transform 1 0 54208 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_476
timestamp 1669390400
transform 1 0 54656 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_483
timestamp 1669390400
transform 1 0 55440 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_491
timestamp 1669390400
transform 1 0 56336 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_495
timestamp 1669390400
transform 1 0 56784 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_499
timestamp 1669390400
transform 1 0 57232 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_512
timestamp 1669390400
transform 1 0 58688 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_516
timestamp 1669390400
transform 1 0 59136 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_522
timestamp 1669390400
transform 1 0 59808 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_39_532
timestamp 1669390400
transform 1 0 60928 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_553
timestamp 1669390400
transform 1 0 63280 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_561
timestamp 1669390400
transform 1 0 64176 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_565
timestamp 1669390400
transform 1 0 64624 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_567
timestamp 1669390400
transform 1 0 64848 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_570
timestamp 1669390400
transform 1 0 65184 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_572
timestamp 1669390400
transform 1 0 65408 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_39_579
timestamp 1669390400
transform 1 0 66192 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_611
timestamp 1669390400
transform 1 0 69776 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_617
timestamp 1669390400
transform 1 0 70448 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_625
timestamp 1669390400
transform 1 0 71344 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_631
timestamp 1669390400
transform 1 0 72016 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_635
timestamp 1669390400
transform 1 0 72464 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_641
timestamp 1669390400
transform 1 0 73136 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_643
timestamp 1669390400
transform 1 0 73360 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_646
timestamp 1669390400
transform 1 0 73696 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_654
timestamp 1669390400
transform 1 0 74592 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_670
timestamp 1669390400
transform 1 0 76384 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_678
timestamp 1669390400
transform 1 0 77280 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_686
timestamp 1669390400
transform 1 0 78176 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_2
timestamp 1669390400
transform 1 0 1568 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_17
timestamp 1669390400
transform 1 0 3248 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_25
timestamp 1669390400
transform 1 0 4144 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_29
timestamp 1669390400
transform 1 0 4592 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_33
timestamp 1669390400
transform 1 0 5040 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_40_37
timestamp 1669390400
transform 1 0 5488 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_40_69
timestamp 1669390400
transform 1 0 9072 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_97
timestamp 1669390400
transform 1 0 12208 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_105
timestamp 1669390400
transform 1 0 13104 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_108
timestamp 1669390400
transform 1 0 13440 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_110
timestamp 1669390400
transform 1 0 13664 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_123
timestamp 1669390400
transform 1 0 15120 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_127
timestamp 1669390400
transform 1 0 15568 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_130
timestamp 1669390400
transform 1 0 15904 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_144
timestamp 1669390400
transform 1 0 17472 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_148
timestamp 1669390400
transform 1 0 17920 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_151
timestamp 1669390400
transform 1 0 18256 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_159
timestamp 1669390400
transform 1 0 19152 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_169
timestamp 1669390400
transform 1 0 20272 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_173
timestamp 1669390400
transform 1 0 20720 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_179
timestamp 1669390400
transform 1 0 21392 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_185
timestamp 1669390400
transform 1 0 22064 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_195
timestamp 1669390400
transform 1 0 23184 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_40_202
timestamp 1669390400
transform 1 0 23968 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_212
timestamp 1669390400
transform 1 0 25088 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_221
timestamp 1669390400
transform 1 0 26096 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_235
timestamp 1669390400
transform 1 0 27664 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_239
timestamp 1669390400
transform 1 0 28112 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_247
timestamp 1669390400
transform 1 0 29008 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_250
timestamp 1669390400
transform 1 0 29344 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_254
timestamp 1669390400
transform 1 0 29792 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_262
timestamp 1669390400
transform 1 0 30688 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_277
timestamp 1669390400
transform 1 0 32368 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_40_281
timestamp 1669390400
transform 1 0 32816 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_289
timestamp 1669390400
transform 1 0 33712 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_293
timestamp 1669390400
transform 1 0 34160 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_295
timestamp 1669390400
transform 1 0 34384 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_308
timestamp 1669390400
transform 1 0 35840 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_318
timestamp 1669390400
transform 1 0 36960 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_321
timestamp 1669390400
transform 1 0 37296 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_40_328
timestamp 1669390400
transform 1 0 38080 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_336
timestamp 1669390400
transform 1 0 38976 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_338
timestamp 1669390400
transform 1 0 39200 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_351
timestamp 1669390400
transform 1 0 40656 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_355
timestamp 1669390400
transform 1 0 41104 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_361
timestamp 1669390400
transform 1 0 41776 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_365
timestamp 1669390400
transform 1 0 42224 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_389
timestamp 1669390400
transform 1 0 44912 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_392
timestamp 1669390400
transform 1 0 45248 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_395
timestamp 1669390400
transform 1 0 45584 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_399
timestamp 1669390400
transform 1 0 46032 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_402
timestamp 1669390400
transform 1 0 46368 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_406
timestamp 1669390400
transform 1 0 46816 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_414
timestamp 1669390400
transform 1 0 47712 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_424
timestamp 1669390400
transform 1 0 48832 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_426
timestamp 1669390400
transform 1 0 49056 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_429
timestamp 1669390400
transform 1 0 49392 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_439
timestamp 1669390400
transform 1 0 50512 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_447
timestamp 1669390400
transform 1 0 51408 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_455
timestamp 1669390400
transform 1 0 52304 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_459
timestamp 1669390400
transform 1 0 52752 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_40_463
timestamp 1669390400
transform 1 0 53200 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_471
timestamp 1669390400
transform 1 0 54096 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_475
timestamp 1669390400
transform 1 0 54544 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_490
timestamp 1669390400
transform 1 0 56224 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_500
timestamp 1669390400
transform 1 0 57344 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_504
timestamp 1669390400
transform 1 0 57792 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_506
timestamp 1669390400
transform 1 0 58016 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_509
timestamp 1669390400
transform 1 0 58352 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_511
timestamp 1669390400
transform 1 0 58576 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_525
timestamp 1669390400
transform 1 0 60144 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_529
timestamp 1669390400
transform 1 0 60592 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_531
timestamp 1669390400
transform 1 0 60816 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_534
timestamp 1669390400
transform 1 0 61152 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_537
timestamp 1669390400
transform 1 0 61488 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_541
timestamp 1669390400
transform 1 0 61936 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_554
timestamp 1669390400
transform 1 0 63392 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_562
timestamp 1669390400
transform 1 0 64288 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_564
timestamp 1669390400
transform 1 0 64512 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_575
timestamp 1669390400
transform 1 0 65744 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_585
timestamp 1669390400
transform 1 0 66864 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_40_589
timestamp 1669390400
transform 1 0 67312 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_597
timestamp 1669390400
transform 1 0 68208 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_601
timestamp 1669390400
transform 1 0 68656 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_605
timestamp 1669390400
transform 1 0 69104 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_629
timestamp 1669390400
transform 1 0 71792 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_636
timestamp 1669390400
transform 1 0 72576 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_640
timestamp 1669390400
transform 1 0 73024 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_647
timestamp 1669390400
transform 1 0 73808 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_651
timestamp 1669390400
transform 1 0 74256 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_655
timestamp 1669390400
transform 1 0 74704 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_670
timestamp 1669390400
transform 1 0 76384 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_676
timestamp 1669390400
transform 1 0 77056 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_683
timestamp 1669390400
transform 1 0 77840 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_687
timestamp 1669390400
transform 1 0 78288 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_2
timestamp 1669390400
transform 1 0 1568 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_17
timestamp 1669390400
transform 1 0 3248 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_25
timestamp 1669390400
transform 1 0 4144 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_33
timestamp 1669390400
transform 1 0 5040 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_41_37
timestamp 1669390400
transform 1 0 5488 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_69
timestamp 1669390400
transform 1 0 9072 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_41_73
timestamp 1669390400
transform 1 0 9520 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_83
timestamp 1669390400
transform 1 0 10640 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_87
timestamp 1669390400
transform 1 0 11088 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_91
timestamp 1669390400
transform 1 0 11536 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_98
timestamp 1669390400
transform 1 0 12320 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_113
timestamp 1669390400
transform 1 0 14000 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_117
timestamp 1669390400
transform 1 0 14448 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_125
timestamp 1669390400
transform 1 0 15344 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_140
timestamp 1669390400
transform 1 0 17024 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_144
timestamp 1669390400
transform 1 0 17472 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_159
timestamp 1669390400
transform 1 0 19152 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_173
timestamp 1669390400
transform 1 0 20720 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_177
timestamp 1669390400
transform 1 0 21168 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_190
timestamp 1669390400
transform 1 0 22624 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_204
timestamp 1669390400
transform 1 0 24192 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_212
timestamp 1669390400
transform 1 0 25088 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_215
timestamp 1669390400
transform 1 0 25424 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_219
timestamp 1669390400
transform 1 0 25872 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_229
timestamp 1669390400
transform 1 0 26992 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_247
timestamp 1669390400
transform 1 0 29008 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_262
timestamp 1669390400
transform 1 0 30688 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_269
timestamp 1669390400
transform 1 0 31472 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_283
timestamp 1669390400
transform 1 0 33040 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_286
timestamp 1669390400
transform 1 0 33376 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_293
timestamp 1669390400
transform 1 0 34160 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_307
timestamp 1669390400
transform 1 0 35728 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_311
timestamp 1669390400
transform 1 0 36176 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_326
timestamp 1669390400
transform 1 0 37856 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_330
timestamp 1669390400
transform 1 0 38304 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_348
timestamp 1669390400
transform 1 0 40320 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_352
timestamp 1669390400
transform 1 0 40768 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_354
timestamp 1669390400
transform 1 0 40992 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_357
timestamp 1669390400
transform 1 0 41328 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_371
timestamp 1669390400
transform 1 0 42896 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_375
timestamp 1669390400
transform 1 0 43344 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_377
timestamp 1669390400
transform 1 0 43568 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_392
timestamp 1669390400
transform 1 0 45248 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_407
timestamp 1669390400
transform 1 0 46928 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_411
timestamp 1669390400
transform 1 0 47376 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_425
timestamp 1669390400
transform 1 0 48944 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_428
timestamp 1669390400
transform 1 0 49280 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_435
timestamp 1669390400
transform 1 0 50064 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_441
timestamp 1669390400
transform 1 0 50736 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_455
timestamp 1669390400
transform 1 0 52304 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_459
timestamp 1669390400
transform 1 0 52752 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_463
timestamp 1669390400
transform 1 0 53200 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_41_466
timestamp 1669390400
transform 1 0 53536 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_474
timestamp 1669390400
transform 1 0 54432 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_478
timestamp 1669390400
transform 1 0 54880 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_480
timestamp 1669390400
transform 1 0 55104 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_483
timestamp 1669390400
transform 1 0 55440 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_495
timestamp 1669390400
transform 1 0 56784 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_499
timestamp 1669390400
transform 1 0 57232 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_508
timestamp 1669390400
transform 1 0 58240 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_512
timestamp 1669390400
transform 1 0 58688 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_525
timestamp 1669390400
transform 1 0 60144 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_531
timestamp 1669390400
transform 1 0 60816 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_533
timestamp 1669390400
transform 1 0 61040 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_546
timestamp 1669390400
transform 1 0 62496 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_554
timestamp 1669390400
transform 1 0 63392 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_558
timestamp 1669390400
transform 1 0 63840 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_567
timestamp 1669390400
transform 1 0 64848 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_570
timestamp 1669390400
transform 1 0 65184 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_584
timestamp 1669390400
transform 1 0 66752 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_592
timestamp 1669390400
transform 1 0 67648 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_596
timestamp 1669390400
transform 1 0 68096 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_600
timestamp 1669390400
transform 1 0 68544 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_606
timestamp 1669390400
transform 1 0 69216 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_612
timestamp 1669390400
transform 1 0 69888 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_622
timestamp 1669390400
transform 1 0 71008 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_626
timestamp 1669390400
transform 1 0 71456 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_630
timestamp 1669390400
transform 1 0 71904 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_638
timestamp 1669390400
transform 1 0 72800 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_641
timestamp 1669390400
transform 1 0 73136 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_644
timestamp 1669390400
transform 1 0 73472 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_654
timestamp 1669390400
transform 1 0 74592 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_670
timestamp 1669390400
transform 1 0 76384 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_686
timestamp 1669390400
transform 1 0 78176 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_2
timestamp 1669390400
transform 1 0 1568 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_18
timestamp 1669390400
transform 1 0 3360 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_34
timestamp 1669390400
transform 1 0 5152 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_37
timestamp 1669390400
transform 1 0 5488 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_40
timestamp 1669390400
transform 1 0 5824 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_44
timestamp 1669390400
transform 1 0 6272 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_62
timestamp 1669390400
transform 1 0 8288 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_66
timestamp 1669390400
transform 1 0 8736 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_72
timestamp 1669390400
transform 1 0 9408 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_87
timestamp 1669390400
transform 1 0 11088 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_89
timestamp 1669390400
transform 1 0 11312 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_104
timestamp 1669390400
transform 1 0 12992 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_107
timestamp 1669390400
transform 1 0 13328 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_109
timestamp 1669390400
transform 1 0 13552 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_112
timestamp 1669390400
transform 1 0 13888 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_128
timestamp 1669390400
transform 1 0 15680 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_132
timestamp 1669390400
transform 1 0 16128 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_139
timestamp 1669390400
transform 1 0 16912 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_142
timestamp 1669390400
transform 1 0 17248 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_151
timestamp 1669390400
transform 1 0 18256 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_153
timestamp 1669390400
transform 1 0 18480 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_156
timestamp 1669390400
transform 1 0 18816 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_172
timestamp 1669390400
transform 1 0 20608 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_174
timestamp 1669390400
transform 1 0 20832 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_177
timestamp 1669390400
transform 1 0 21168 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_193
timestamp 1669390400
transform 1 0 22960 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_209
timestamp 1669390400
transform 1 0 24752 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_212
timestamp 1669390400
transform 1 0 25088 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_215
timestamp 1669390400
transform 1 0 25424 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_222
timestamp 1669390400
transform 1 0 26208 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_238
timestamp 1669390400
transform 1 0 28000 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_244
timestamp 1669390400
transform 1 0 28672 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_247
timestamp 1669390400
transform 1 0 29008 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_262
timestamp 1669390400
transform 1 0 30688 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_264
timestamp 1669390400
transform 1 0 30912 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_279
timestamp 1669390400
transform 1 0 32592 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_282
timestamp 1669390400
transform 1 0 32928 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_288
timestamp 1669390400
transform 1 0 33600 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_304
timestamp 1669390400
transform 1 0 35392 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_314
timestamp 1669390400
transform 1 0 36512 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_317
timestamp 1669390400
transform 1 0 36848 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_42_342
timestamp 1669390400
transform 1 0 39648 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_352
timestamp 1669390400
transform 1 0 40768 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_370
timestamp 1669390400
transform 1 0 42784 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_374
timestamp 1669390400
transform 1 0 43232 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_384
timestamp 1669390400
transform 1 0 44352 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_387
timestamp 1669390400
transform 1 0 44688 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_396
timestamp 1669390400
transform 1 0 45696 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_414
timestamp 1669390400
transform 1 0 47712 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_418
timestamp 1669390400
transform 1 0 48160 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_422
timestamp 1669390400
transform 1 0 48608 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_437
timestamp 1669390400
transform 1 0 50288 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_439
timestamp 1669390400
transform 1 0 50512 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_454
timestamp 1669390400
transform 1 0 52192 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_457
timestamp 1669390400
transform 1 0 52528 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_464
timestamp 1669390400
transform 1 0 53312 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_42_480
timestamp 1669390400
transform 1 0 55104 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_488
timestamp 1669390400
transform 1 0 56000 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_492
timestamp 1669390400
transform 1 0 56448 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_507
timestamp 1669390400
transform 1 0 58128 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_509
timestamp 1669390400
transform 1 0 58352 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_524
timestamp 1669390400
transform 1 0 60032 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_527
timestamp 1669390400
transform 1 0 60368 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_530
timestamp 1669390400
transform 1 0 60704 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_546
timestamp 1669390400
transform 1 0 62496 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_554
timestamp 1669390400
transform 1 0 63392 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_556
timestamp 1669390400
transform 1 0 63616 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_559
timestamp 1669390400
transform 1 0 63952 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_562
timestamp 1669390400
transform 1 0 64288 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_577
timestamp 1669390400
transform 1 0 65968 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_593
timestamp 1669390400
transform 1 0 67760 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_597
timestamp 1669390400
transform 1 0 68208 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_612
timestamp 1669390400
transform 1 0 69888 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_614
timestamp 1669390400
transform 1 0 70112 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_629
timestamp 1669390400
transform 1 0 71792 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_632
timestamp 1669390400
transform 1 0 72128 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_640
timestamp 1669390400
transform 1 0 73024 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_656
timestamp 1669390400
transform 1 0 74816 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_664
timestamp 1669390400
transform 1 0 75712 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_667
timestamp 1669390400
transform 1 0 76048 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_682
timestamp 1669390400
transform 1 0 77728 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_686
timestamp 1669390400
transform 1 0 78176 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_0 Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_1
timestamp 1669390400
transform -1 0 78624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_2
timestamp 1669390400
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_3
timestamp 1669390400
transform -1 0 78624 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_4
timestamp 1669390400
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_5
timestamp 1669390400
transform -1 0 78624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_6
timestamp 1669390400
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_7
timestamp 1669390400
transform -1 0 78624 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_8
timestamp 1669390400
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_9
timestamp 1669390400
transform -1 0 78624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_10
timestamp 1669390400
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_11
timestamp 1669390400
transform -1 0 78624 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_12
timestamp 1669390400
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_13
timestamp 1669390400
transform -1 0 78624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_14
timestamp 1669390400
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_15
timestamp 1669390400
transform -1 0 78624 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_16
timestamp 1669390400
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_17
timestamp 1669390400
transform -1 0 78624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_18
timestamp 1669390400
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_19
timestamp 1669390400
transform -1 0 78624 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_20
timestamp 1669390400
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_21
timestamp 1669390400
transform -1 0 78624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_22
timestamp 1669390400
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_23
timestamp 1669390400
transform -1 0 78624 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_24
timestamp 1669390400
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_25
timestamp 1669390400
transform -1 0 78624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_26
timestamp 1669390400
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_27
timestamp 1669390400
transform -1 0 78624 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_28
timestamp 1669390400
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_29
timestamp 1669390400
transform -1 0 78624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_30
timestamp 1669390400
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_31
timestamp 1669390400
transform -1 0 78624 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_32
timestamp 1669390400
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_33
timestamp 1669390400
transform -1 0 78624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_34
timestamp 1669390400
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_35
timestamp 1669390400
transform -1 0 78624 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_36
timestamp 1669390400
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_37
timestamp 1669390400
transform -1 0 78624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_38
timestamp 1669390400
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_39
timestamp 1669390400
transform -1 0 78624 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_40
timestamp 1669390400
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_41
timestamp 1669390400
transform -1 0 78624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_42
timestamp 1669390400
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_43
timestamp 1669390400
transform -1 0 78624 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_44
timestamp 1669390400
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_45
timestamp 1669390400
transform -1 0 78624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_46
timestamp 1669390400
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_47
timestamp 1669390400
transform -1 0 78624 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_48
timestamp 1669390400
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_49
timestamp 1669390400
transform -1 0 78624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_50
timestamp 1669390400
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_51
timestamp 1669390400
transform -1 0 78624 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_52
timestamp 1669390400
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_53
timestamp 1669390400
transform -1 0 78624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_54
timestamp 1669390400
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_55
timestamp 1669390400
transform -1 0 78624 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_56
timestamp 1669390400
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_57
timestamp 1669390400
transform -1 0 78624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_58
timestamp 1669390400
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_59
timestamp 1669390400
transform -1 0 78624 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_60
timestamp 1669390400
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_61
timestamp 1669390400
transform -1 0 78624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_62
timestamp 1669390400
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_63
timestamp 1669390400
transform -1 0 78624 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_64
timestamp 1669390400
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_65
timestamp 1669390400
transform -1 0 78624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_66
timestamp 1669390400
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_67
timestamp 1669390400
transform -1 0 78624 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_68
timestamp 1669390400
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_69
timestamp 1669390400
transform -1 0 78624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_70
timestamp 1669390400
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_71
timestamp 1669390400
transform -1 0 78624 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_72
timestamp 1669390400
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_73
timestamp 1669390400
transform -1 0 78624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_74
timestamp 1669390400
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_75
timestamp 1669390400
transform -1 0 78624 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_76
timestamp 1669390400
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_77
timestamp 1669390400
transform -1 0 78624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_78
timestamp 1669390400
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_79
timestamp 1669390400
transform -1 0 78624 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_80
timestamp 1669390400
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_81
timestamp 1669390400
transform -1 0 78624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_82
timestamp 1669390400
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_83
timestamp 1669390400
transform -1 0 78624 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_84
timestamp 1669390400
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_85
timestamp 1669390400
transform -1 0 78624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_86 Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 5264 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_87
timestamp 1669390400
transform 1 0 9184 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_88
timestamp 1669390400
transform 1 0 13104 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_89
timestamp 1669390400
transform 1 0 17024 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_90
timestamp 1669390400
transform 1 0 20944 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_91
timestamp 1669390400
transform 1 0 24864 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_92
timestamp 1669390400
transform 1 0 28784 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_93
timestamp 1669390400
transform 1 0 32704 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_94
timestamp 1669390400
transform 1 0 36624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_95
timestamp 1669390400
transform 1 0 40544 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_96
timestamp 1669390400
transform 1 0 44464 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_97
timestamp 1669390400
transform 1 0 48384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_98
timestamp 1669390400
transform 1 0 52304 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_99
timestamp 1669390400
transform 1 0 56224 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_100
timestamp 1669390400
transform 1 0 60144 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_101
timestamp 1669390400
transform 1 0 64064 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_102
timestamp 1669390400
transform 1 0 67984 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_103
timestamp 1669390400
transform 1 0 71904 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_104
timestamp 1669390400
transform 1 0 75824 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_105
timestamp 1669390400
transform 1 0 9296 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_106
timestamp 1669390400
transform 1 0 17248 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_107
timestamp 1669390400
transform 1 0 25200 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_108
timestamp 1669390400
transform 1 0 33152 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_109
timestamp 1669390400
transform 1 0 41104 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_110
timestamp 1669390400
transform 1 0 49056 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_111
timestamp 1669390400
transform 1 0 57008 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_112
timestamp 1669390400
transform 1 0 64960 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_113
timestamp 1669390400
transform 1 0 72912 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_114
timestamp 1669390400
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_115
timestamp 1669390400
transform 1 0 13216 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_116
timestamp 1669390400
transform 1 0 21168 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_117
timestamp 1669390400
transform 1 0 29120 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_118
timestamp 1669390400
transform 1 0 37072 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_119
timestamp 1669390400
transform 1 0 45024 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_120
timestamp 1669390400
transform 1 0 52976 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_121
timestamp 1669390400
transform 1 0 60928 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_122
timestamp 1669390400
transform 1 0 68880 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_123
timestamp 1669390400
transform 1 0 76832 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_124
timestamp 1669390400
transform 1 0 9296 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_125
timestamp 1669390400
transform 1 0 17248 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_126
timestamp 1669390400
transform 1 0 25200 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_127
timestamp 1669390400
transform 1 0 33152 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_128
timestamp 1669390400
transform 1 0 41104 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_129
timestamp 1669390400
transform 1 0 49056 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_130
timestamp 1669390400
transform 1 0 57008 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_131
timestamp 1669390400
transform 1 0 64960 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_132
timestamp 1669390400
transform 1 0 72912 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_133
timestamp 1669390400
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_134
timestamp 1669390400
transform 1 0 13216 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_135
timestamp 1669390400
transform 1 0 21168 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_136
timestamp 1669390400
transform 1 0 29120 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_137
timestamp 1669390400
transform 1 0 37072 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_138
timestamp 1669390400
transform 1 0 45024 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_139
timestamp 1669390400
transform 1 0 52976 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_140
timestamp 1669390400
transform 1 0 60928 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_141
timestamp 1669390400
transform 1 0 68880 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_142
timestamp 1669390400
transform 1 0 76832 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_143
timestamp 1669390400
transform 1 0 9296 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_144
timestamp 1669390400
transform 1 0 17248 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_145
timestamp 1669390400
transform 1 0 25200 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_146
timestamp 1669390400
transform 1 0 33152 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_147
timestamp 1669390400
transform 1 0 41104 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_148
timestamp 1669390400
transform 1 0 49056 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_149
timestamp 1669390400
transform 1 0 57008 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_150
timestamp 1669390400
transform 1 0 64960 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_151
timestamp 1669390400
transform 1 0 72912 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_152
timestamp 1669390400
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_153
timestamp 1669390400
transform 1 0 13216 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_154
timestamp 1669390400
transform 1 0 21168 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_155
timestamp 1669390400
transform 1 0 29120 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_156
timestamp 1669390400
transform 1 0 37072 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_157
timestamp 1669390400
transform 1 0 45024 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_158
timestamp 1669390400
transform 1 0 52976 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_159
timestamp 1669390400
transform 1 0 60928 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_160
timestamp 1669390400
transform 1 0 68880 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_161
timestamp 1669390400
transform 1 0 76832 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_162
timestamp 1669390400
transform 1 0 9296 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_163
timestamp 1669390400
transform 1 0 17248 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_164
timestamp 1669390400
transform 1 0 25200 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_165
timestamp 1669390400
transform 1 0 33152 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_166
timestamp 1669390400
transform 1 0 41104 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_167
timestamp 1669390400
transform 1 0 49056 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_168
timestamp 1669390400
transform 1 0 57008 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_169
timestamp 1669390400
transform 1 0 64960 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_170
timestamp 1669390400
transform 1 0 72912 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_171
timestamp 1669390400
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_172
timestamp 1669390400
transform 1 0 13216 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_173
timestamp 1669390400
transform 1 0 21168 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_174
timestamp 1669390400
transform 1 0 29120 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_175
timestamp 1669390400
transform 1 0 37072 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_176
timestamp 1669390400
transform 1 0 45024 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_177
timestamp 1669390400
transform 1 0 52976 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_178
timestamp 1669390400
transform 1 0 60928 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_179
timestamp 1669390400
transform 1 0 68880 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_180
timestamp 1669390400
transform 1 0 76832 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_181
timestamp 1669390400
transform 1 0 9296 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_182
timestamp 1669390400
transform 1 0 17248 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_183
timestamp 1669390400
transform 1 0 25200 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_184
timestamp 1669390400
transform 1 0 33152 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_185
timestamp 1669390400
transform 1 0 41104 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_186
timestamp 1669390400
transform 1 0 49056 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_187
timestamp 1669390400
transform 1 0 57008 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_188
timestamp 1669390400
transform 1 0 64960 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_189
timestamp 1669390400
transform 1 0 72912 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_190
timestamp 1669390400
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_191
timestamp 1669390400
transform 1 0 13216 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_192
timestamp 1669390400
transform 1 0 21168 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_193
timestamp 1669390400
transform 1 0 29120 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_194
timestamp 1669390400
transform 1 0 37072 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_195
timestamp 1669390400
transform 1 0 45024 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_196
timestamp 1669390400
transform 1 0 52976 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_197
timestamp 1669390400
transform 1 0 60928 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_198
timestamp 1669390400
transform 1 0 68880 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_199
timestamp 1669390400
transform 1 0 76832 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_200
timestamp 1669390400
transform 1 0 9296 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_201
timestamp 1669390400
transform 1 0 17248 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_202
timestamp 1669390400
transform 1 0 25200 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_203
timestamp 1669390400
transform 1 0 33152 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_204
timestamp 1669390400
transform 1 0 41104 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_205
timestamp 1669390400
transform 1 0 49056 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_206
timestamp 1669390400
transform 1 0 57008 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_207
timestamp 1669390400
transform 1 0 64960 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_208
timestamp 1669390400
transform 1 0 72912 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_209
timestamp 1669390400
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_210
timestamp 1669390400
transform 1 0 13216 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_211
timestamp 1669390400
transform 1 0 21168 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_212
timestamp 1669390400
transform 1 0 29120 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_213
timestamp 1669390400
transform 1 0 37072 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_214
timestamp 1669390400
transform 1 0 45024 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_215
timestamp 1669390400
transform 1 0 52976 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_216
timestamp 1669390400
transform 1 0 60928 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_217
timestamp 1669390400
transform 1 0 68880 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_218
timestamp 1669390400
transform 1 0 76832 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_219
timestamp 1669390400
transform 1 0 9296 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_220
timestamp 1669390400
transform 1 0 17248 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_221
timestamp 1669390400
transform 1 0 25200 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_222
timestamp 1669390400
transform 1 0 33152 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_223
timestamp 1669390400
transform 1 0 41104 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_224
timestamp 1669390400
transform 1 0 49056 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_225
timestamp 1669390400
transform 1 0 57008 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_226
timestamp 1669390400
transform 1 0 64960 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_227
timestamp 1669390400
transform 1 0 72912 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_228
timestamp 1669390400
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_229
timestamp 1669390400
transform 1 0 13216 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_230
timestamp 1669390400
transform 1 0 21168 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_231
timestamp 1669390400
transform 1 0 29120 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_232
timestamp 1669390400
transform 1 0 37072 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_233
timestamp 1669390400
transform 1 0 45024 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_234
timestamp 1669390400
transform 1 0 52976 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_235
timestamp 1669390400
transform 1 0 60928 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_236
timestamp 1669390400
transform 1 0 68880 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_237
timestamp 1669390400
transform 1 0 76832 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_238
timestamp 1669390400
transform 1 0 9296 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_239
timestamp 1669390400
transform 1 0 17248 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_240
timestamp 1669390400
transform 1 0 25200 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_241
timestamp 1669390400
transform 1 0 33152 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_242
timestamp 1669390400
transform 1 0 41104 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_243
timestamp 1669390400
transform 1 0 49056 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_244
timestamp 1669390400
transform 1 0 57008 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_245
timestamp 1669390400
transform 1 0 64960 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_246
timestamp 1669390400
transform 1 0 72912 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_247
timestamp 1669390400
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_248
timestamp 1669390400
transform 1 0 13216 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_249
timestamp 1669390400
transform 1 0 21168 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_250
timestamp 1669390400
transform 1 0 29120 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_251
timestamp 1669390400
transform 1 0 37072 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_252
timestamp 1669390400
transform 1 0 45024 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_253
timestamp 1669390400
transform 1 0 52976 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_254
timestamp 1669390400
transform 1 0 60928 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_255
timestamp 1669390400
transform 1 0 68880 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_256
timestamp 1669390400
transform 1 0 76832 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_257
timestamp 1669390400
transform 1 0 9296 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_258
timestamp 1669390400
transform 1 0 17248 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_259
timestamp 1669390400
transform 1 0 25200 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_260
timestamp 1669390400
transform 1 0 33152 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_261
timestamp 1669390400
transform 1 0 41104 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_262
timestamp 1669390400
transform 1 0 49056 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_263
timestamp 1669390400
transform 1 0 57008 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_264
timestamp 1669390400
transform 1 0 64960 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_265
timestamp 1669390400
transform 1 0 72912 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_266
timestamp 1669390400
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_267
timestamp 1669390400
transform 1 0 13216 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_268
timestamp 1669390400
transform 1 0 21168 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_269
timestamp 1669390400
transform 1 0 29120 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_270
timestamp 1669390400
transform 1 0 37072 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_271
timestamp 1669390400
transform 1 0 45024 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_272
timestamp 1669390400
transform 1 0 52976 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_273
timestamp 1669390400
transform 1 0 60928 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_274
timestamp 1669390400
transform 1 0 68880 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_275
timestamp 1669390400
transform 1 0 76832 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_276
timestamp 1669390400
transform 1 0 9296 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_277
timestamp 1669390400
transform 1 0 17248 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_278
timestamp 1669390400
transform 1 0 25200 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_279
timestamp 1669390400
transform 1 0 33152 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_280
timestamp 1669390400
transform 1 0 41104 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_281
timestamp 1669390400
transform 1 0 49056 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_282
timestamp 1669390400
transform 1 0 57008 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_283
timestamp 1669390400
transform 1 0 64960 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_284
timestamp 1669390400
transform 1 0 72912 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_285
timestamp 1669390400
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_286
timestamp 1669390400
transform 1 0 13216 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_287
timestamp 1669390400
transform 1 0 21168 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_288
timestamp 1669390400
transform 1 0 29120 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_289
timestamp 1669390400
transform 1 0 37072 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_290
timestamp 1669390400
transform 1 0 45024 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_291
timestamp 1669390400
transform 1 0 52976 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_292
timestamp 1669390400
transform 1 0 60928 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_293
timestamp 1669390400
transform 1 0 68880 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_294
timestamp 1669390400
transform 1 0 76832 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_295
timestamp 1669390400
transform 1 0 9296 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_296
timestamp 1669390400
transform 1 0 17248 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_297
timestamp 1669390400
transform 1 0 25200 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_298
timestamp 1669390400
transform 1 0 33152 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_299
timestamp 1669390400
transform 1 0 41104 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_300
timestamp 1669390400
transform 1 0 49056 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_301
timestamp 1669390400
transform 1 0 57008 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_302
timestamp 1669390400
transform 1 0 64960 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_303
timestamp 1669390400
transform 1 0 72912 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_304
timestamp 1669390400
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_305
timestamp 1669390400
transform 1 0 13216 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_306
timestamp 1669390400
transform 1 0 21168 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_307
timestamp 1669390400
transform 1 0 29120 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_308
timestamp 1669390400
transform 1 0 37072 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_309
timestamp 1669390400
transform 1 0 45024 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_310
timestamp 1669390400
transform 1 0 52976 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_311
timestamp 1669390400
transform 1 0 60928 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_312
timestamp 1669390400
transform 1 0 68880 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_313
timestamp 1669390400
transform 1 0 76832 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_314
timestamp 1669390400
transform 1 0 9296 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_315
timestamp 1669390400
transform 1 0 17248 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_316
timestamp 1669390400
transform 1 0 25200 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_317
timestamp 1669390400
transform 1 0 33152 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_318
timestamp 1669390400
transform 1 0 41104 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_319
timestamp 1669390400
transform 1 0 49056 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_320
timestamp 1669390400
transform 1 0 57008 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_321
timestamp 1669390400
transform 1 0 64960 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_322
timestamp 1669390400
transform 1 0 72912 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_323
timestamp 1669390400
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_324
timestamp 1669390400
transform 1 0 13216 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_325
timestamp 1669390400
transform 1 0 21168 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_326
timestamp 1669390400
transform 1 0 29120 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_327
timestamp 1669390400
transform 1 0 37072 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_328
timestamp 1669390400
transform 1 0 45024 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_329
timestamp 1669390400
transform 1 0 52976 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_330
timestamp 1669390400
transform 1 0 60928 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_331
timestamp 1669390400
transform 1 0 68880 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_332
timestamp 1669390400
transform 1 0 76832 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_333
timestamp 1669390400
transform 1 0 9296 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_334
timestamp 1669390400
transform 1 0 17248 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_335
timestamp 1669390400
transform 1 0 25200 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_336
timestamp 1669390400
transform 1 0 33152 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_337
timestamp 1669390400
transform 1 0 41104 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_338
timestamp 1669390400
transform 1 0 49056 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_339
timestamp 1669390400
transform 1 0 57008 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_340
timestamp 1669390400
transform 1 0 64960 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_341
timestamp 1669390400
transform 1 0 72912 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_342
timestamp 1669390400
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_343
timestamp 1669390400
transform 1 0 13216 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_344
timestamp 1669390400
transform 1 0 21168 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_345
timestamp 1669390400
transform 1 0 29120 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_346
timestamp 1669390400
transform 1 0 37072 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_347
timestamp 1669390400
transform 1 0 45024 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_348
timestamp 1669390400
transform 1 0 52976 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_349
timestamp 1669390400
transform 1 0 60928 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_350
timestamp 1669390400
transform 1 0 68880 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_351
timestamp 1669390400
transform 1 0 76832 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_352
timestamp 1669390400
transform 1 0 9296 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_353
timestamp 1669390400
transform 1 0 17248 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_354
timestamp 1669390400
transform 1 0 25200 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_355
timestamp 1669390400
transform 1 0 33152 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_356
timestamp 1669390400
transform 1 0 41104 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_357
timestamp 1669390400
transform 1 0 49056 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_358
timestamp 1669390400
transform 1 0 57008 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_359
timestamp 1669390400
transform 1 0 64960 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_360
timestamp 1669390400
transform 1 0 72912 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_361
timestamp 1669390400
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_362
timestamp 1669390400
transform 1 0 13216 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_363
timestamp 1669390400
transform 1 0 21168 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_364
timestamp 1669390400
transform 1 0 29120 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_365
timestamp 1669390400
transform 1 0 37072 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_366
timestamp 1669390400
transform 1 0 45024 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_367
timestamp 1669390400
transform 1 0 52976 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_368
timestamp 1669390400
transform 1 0 60928 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_369
timestamp 1669390400
transform 1 0 68880 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_370
timestamp 1669390400
transform 1 0 76832 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_371
timestamp 1669390400
transform 1 0 9296 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_372
timestamp 1669390400
transform 1 0 17248 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_373
timestamp 1669390400
transform 1 0 25200 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_374
timestamp 1669390400
transform 1 0 33152 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_375
timestamp 1669390400
transform 1 0 41104 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_376
timestamp 1669390400
transform 1 0 49056 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_377
timestamp 1669390400
transform 1 0 57008 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_378
timestamp 1669390400
transform 1 0 64960 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_379
timestamp 1669390400
transform 1 0 72912 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_380
timestamp 1669390400
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_381
timestamp 1669390400
transform 1 0 13216 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_382
timestamp 1669390400
transform 1 0 21168 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_383
timestamp 1669390400
transform 1 0 29120 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_384
timestamp 1669390400
transform 1 0 37072 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_385
timestamp 1669390400
transform 1 0 45024 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_386
timestamp 1669390400
transform 1 0 52976 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_387
timestamp 1669390400
transform 1 0 60928 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_388
timestamp 1669390400
transform 1 0 68880 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_389
timestamp 1669390400
transform 1 0 76832 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_390
timestamp 1669390400
transform 1 0 9296 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_391
timestamp 1669390400
transform 1 0 17248 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_392
timestamp 1669390400
transform 1 0 25200 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_393
timestamp 1669390400
transform 1 0 33152 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_394
timestamp 1669390400
transform 1 0 41104 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_395
timestamp 1669390400
transform 1 0 49056 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_396
timestamp 1669390400
transform 1 0 57008 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_397
timestamp 1669390400
transform 1 0 64960 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_398
timestamp 1669390400
transform 1 0 72912 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_399
timestamp 1669390400
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_400
timestamp 1669390400
transform 1 0 13216 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_401
timestamp 1669390400
transform 1 0 21168 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_402
timestamp 1669390400
transform 1 0 29120 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_403
timestamp 1669390400
transform 1 0 37072 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_404
timestamp 1669390400
transform 1 0 45024 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_405
timestamp 1669390400
transform 1 0 52976 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_406
timestamp 1669390400
transform 1 0 60928 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_407
timestamp 1669390400
transform 1 0 68880 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_408
timestamp 1669390400
transform 1 0 76832 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_409
timestamp 1669390400
transform 1 0 9296 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_410
timestamp 1669390400
transform 1 0 17248 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_411
timestamp 1669390400
transform 1 0 25200 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_412
timestamp 1669390400
transform 1 0 33152 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_413
timestamp 1669390400
transform 1 0 41104 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_414
timestamp 1669390400
transform 1 0 49056 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_415
timestamp 1669390400
transform 1 0 57008 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_416
timestamp 1669390400
transform 1 0 64960 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_417
timestamp 1669390400
transform 1 0 72912 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_418
timestamp 1669390400
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_419
timestamp 1669390400
transform 1 0 13216 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_420
timestamp 1669390400
transform 1 0 21168 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_421
timestamp 1669390400
transform 1 0 29120 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_422
timestamp 1669390400
transform 1 0 37072 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_423
timestamp 1669390400
transform 1 0 45024 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_424
timestamp 1669390400
transform 1 0 52976 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_425
timestamp 1669390400
transform 1 0 60928 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_426
timestamp 1669390400
transform 1 0 68880 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_427
timestamp 1669390400
transform 1 0 76832 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_428
timestamp 1669390400
transform 1 0 9296 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_429
timestamp 1669390400
transform 1 0 17248 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_430
timestamp 1669390400
transform 1 0 25200 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_431
timestamp 1669390400
transform 1 0 33152 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_432
timestamp 1669390400
transform 1 0 41104 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_433
timestamp 1669390400
transform 1 0 49056 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_434
timestamp 1669390400
transform 1 0 57008 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_435
timestamp 1669390400
transform 1 0 64960 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_436
timestamp 1669390400
transform 1 0 72912 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_437
timestamp 1669390400
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_438
timestamp 1669390400
transform 1 0 13216 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_439
timestamp 1669390400
transform 1 0 21168 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_440
timestamp 1669390400
transform 1 0 29120 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_441
timestamp 1669390400
transform 1 0 37072 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_442
timestamp 1669390400
transform 1 0 45024 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_443
timestamp 1669390400
transform 1 0 52976 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_444
timestamp 1669390400
transform 1 0 60928 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_445
timestamp 1669390400
transform 1 0 68880 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_446
timestamp 1669390400
transform 1 0 76832 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_447
timestamp 1669390400
transform 1 0 9296 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_448
timestamp 1669390400
transform 1 0 17248 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_449
timestamp 1669390400
transform 1 0 25200 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_450
timestamp 1669390400
transform 1 0 33152 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_451
timestamp 1669390400
transform 1 0 41104 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_452
timestamp 1669390400
transform 1 0 49056 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_453
timestamp 1669390400
transform 1 0 57008 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_454
timestamp 1669390400
transform 1 0 64960 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_455
timestamp 1669390400
transform 1 0 72912 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_456
timestamp 1669390400
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_457
timestamp 1669390400
transform 1 0 13216 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_458
timestamp 1669390400
transform 1 0 21168 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_459
timestamp 1669390400
transform 1 0 29120 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_460
timestamp 1669390400
transform 1 0 37072 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_461
timestamp 1669390400
transform 1 0 45024 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_462
timestamp 1669390400
transform 1 0 52976 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_463
timestamp 1669390400
transform 1 0 60928 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_464
timestamp 1669390400
transform 1 0 68880 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_465
timestamp 1669390400
transform 1 0 76832 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_466
timestamp 1669390400
transform 1 0 9296 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_467
timestamp 1669390400
transform 1 0 17248 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_468
timestamp 1669390400
transform 1 0 25200 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_469
timestamp 1669390400
transform 1 0 33152 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_470
timestamp 1669390400
transform 1 0 41104 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_471
timestamp 1669390400
transform 1 0 49056 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_472
timestamp 1669390400
transform 1 0 57008 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_473
timestamp 1669390400
transform 1 0 64960 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_474
timestamp 1669390400
transform 1 0 72912 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_475
timestamp 1669390400
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_476
timestamp 1669390400
transform 1 0 13216 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_477
timestamp 1669390400
transform 1 0 21168 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_478
timestamp 1669390400
transform 1 0 29120 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_479
timestamp 1669390400
transform 1 0 37072 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_480
timestamp 1669390400
transform 1 0 45024 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_481
timestamp 1669390400
transform 1 0 52976 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_482
timestamp 1669390400
transform 1 0 60928 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_483
timestamp 1669390400
transform 1 0 68880 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_484
timestamp 1669390400
transform 1 0 76832 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_485
timestamp 1669390400
transform 1 0 9296 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_486
timestamp 1669390400
transform 1 0 17248 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_487
timestamp 1669390400
transform 1 0 25200 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_488
timestamp 1669390400
transform 1 0 33152 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_489
timestamp 1669390400
transform 1 0 41104 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_490
timestamp 1669390400
transform 1 0 49056 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_491
timestamp 1669390400
transform 1 0 57008 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_492
timestamp 1669390400
transform 1 0 64960 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_493
timestamp 1669390400
transform 1 0 72912 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_494
timestamp 1669390400
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_495
timestamp 1669390400
transform 1 0 9184 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_496
timestamp 1669390400
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_497
timestamp 1669390400
transform 1 0 17024 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_498
timestamp 1669390400
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_499
timestamp 1669390400
transform 1 0 24864 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_500
timestamp 1669390400
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_501
timestamp 1669390400
transform 1 0 32704 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_502
timestamp 1669390400
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_503
timestamp 1669390400
transform 1 0 40544 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_504
timestamp 1669390400
transform 1 0 44464 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_505
timestamp 1669390400
transform 1 0 48384 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_506
timestamp 1669390400
transform 1 0 52304 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_507
timestamp 1669390400
transform 1 0 56224 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_508
timestamp 1669390400
transform 1 0 60144 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_509
timestamp 1669390400
transform 1 0 64064 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_510
timestamp 1669390400
transform 1 0 67984 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_511
timestamp 1669390400
transform 1 0 71904 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_512
timestamp 1669390400
transform 1 0 75824 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1387_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 2128 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1388_
timestamp 1669390400
transform 1 0 36624 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1389_
timestamp 1669390400
transform -1 0 22848 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1390_
timestamp 1669390400
transform 1 0 21504 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1391_
timestamp 1669390400
transform 1 0 22064 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1392_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 20160 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1393_
timestamp 1669390400
transform 1 0 46144 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1394_
timestamp 1669390400
transform 1 0 19264 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1395_
timestamp 1669390400
transform 1 0 20048 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1396_
timestamp 1669390400
transform 1 0 21952 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1397_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 23408 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1398_
timestamp 1669390400
transform 1 0 23632 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1399_
timestamp 1669390400
transform -1 0 19264 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1400_
timestamp 1669390400
transform -1 0 44352 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1401_
timestamp 1669390400
transform 1 0 16576 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1402_
timestamp 1669390400
transform 1 0 14560 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1403_
timestamp 1669390400
transform 1 0 22848 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1404_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 17584 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _1405_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 18368 0 1 28224
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1406_
timestamp 1669390400
transform 1 0 23296 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1407_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 24416 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1408_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 23072 0 -1 28224
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1409_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 21952 0 -1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1410_
timestamp 1669390400
transform 1 0 23520 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1411_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 21728 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1412_
timestamp 1669390400
transform -1 0 15792 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1413_
timestamp 1669390400
transform -1 0 14784 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1414_
timestamp 1669390400
transform -1 0 15232 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1415_
timestamp 1669390400
transform -1 0 18592 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1416_
timestamp 1669390400
transform -1 0 19376 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1417_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 18144 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1418_
timestamp 1669390400
transform 1 0 17920 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1419_
timestamp 1669390400
transform 1 0 16576 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1420_
timestamp 1669390400
transform 1 0 6944 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1421_
timestamp 1669390400
transform 1 0 23968 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1422_
timestamp 1669390400
transform -1 0 20720 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1423_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 17584 0 -1 26656
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1424_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 18480 0 1 29792
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1425_
timestamp 1669390400
transform 1 0 19488 0 -1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1426_
timestamp 1669390400
transform 1 0 21504 0 1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1427_
timestamp 1669390400
transform 1 0 22176 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1428_
timestamp 1669390400
transform -1 0 21056 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1429_
timestamp 1669390400
transform 1 0 13104 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1430_
timestamp 1669390400
transform -1 0 46704 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1431_
timestamp 1669390400
transform 1 0 48272 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1432_
timestamp 1669390400
transform -1 0 15344 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1433_
timestamp 1669390400
transform -1 0 14448 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1434_
timestamp 1669390400
transform -1 0 14560 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1435_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 15008 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1436_
timestamp 1669390400
transform 1 0 13888 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1437_
timestamp 1669390400
transform -1 0 20944 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1438_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 22512 0 1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _1439_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 17808 0 1 25088
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1440_
timestamp 1669390400
transform 1 0 18144 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1441_
timestamp 1669390400
transform 1 0 13552 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1442_
timestamp 1669390400
transform 1 0 25536 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1443_
timestamp 1669390400
transform -1 0 20944 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _1444_
timestamp 1669390400
transform -1 0 20944 0 -1 25088
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1445_
timestamp 1669390400
transform 1 0 15680 0 -1 31360
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1446_
timestamp 1669390400
transform 1 0 16576 0 1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1447_
timestamp 1669390400
transform 1 0 18816 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1448_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 18368 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1449_
timestamp 1669390400
transform 1 0 17696 0 1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1450_
timestamp 1669390400
transform 1 0 18592 0 -1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1451_
timestamp 1669390400
transform 1 0 19488 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1452_
timestamp 1669390400
transform -1 0 15904 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1453_
timestamp 1669390400
transform -1 0 16352 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1454_
timestamp 1669390400
transform 1 0 14560 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1455_
timestamp 1669390400
transform -1 0 55216 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1456_
timestamp 1669390400
transform -1 0 12992 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1457_
timestamp 1669390400
transform -1 0 9184 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1458_
timestamp 1669390400
transform -1 0 11872 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1459_
timestamp 1669390400
transform -1 0 11648 0 -1 28224
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1460_
timestamp 1669390400
transform 1 0 9968 0 1 28224
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1461_
timestamp 1669390400
transform -1 0 21728 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1462_
timestamp 1669390400
transform -1 0 23408 0 -1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1463_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 19152 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1464_
timestamp 1669390400
transform 1 0 18928 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1465_
timestamp 1669390400
transform 1 0 3808 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1466_
timestamp 1669390400
transform 1 0 47488 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1467_
timestamp 1669390400
transform -1 0 21056 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _1468_
timestamp 1669390400
transform -1 0 22400 0 -1 23520
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1469_
timestamp 1669390400
transform -1 0 11872 0 -1 29792
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1470_
timestamp 1669390400
transform 1 0 11312 0 1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1471_
timestamp 1669390400
transform -1 0 15008 0 1 31360
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1472_
timestamp 1669390400
transform 1 0 13664 0 -1 32928
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1473_
timestamp 1669390400
transform -1 0 18144 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1474_
timestamp 1669390400
transform -1 0 19152 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1475_
timestamp 1669390400
transform 1 0 11760 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1476_
timestamp 1669390400
transform -1 0 14000 0 -1 36064
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1477_
timestamp 1669390400
transform 1 0 12432 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1478_
timestamp 1669390400
transform 1 0 17584 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1479_
timestamp 1669390400
transform -1 0 11760 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1480_
timestamp 1669390400
transform 1 0 9968 0 1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1481_
timestamp 1669390400
transform -1 0 56112 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1482_
timestamp 1669390400
transform 1 0 6496 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1483_
timestamp 1669390400
transform 1 0 7168 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1484_
timestamp 1669390400
transform 1 0 7616 0 -1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1485_
timestamp 1669390400
transform -1 0 12656 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1486_
timestamp 1669390400
transform 1 0 10192 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1487_
timestamp 1669390400
transform -1 0 20384 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1488_
timestamp 1669390400
transform -1 0 22512 0 1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1489_
timestamp 1669390400
transform -1 0 20832 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1490_
timestamp 1669390400
transform 1 0 16576 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1491_
timestamp 1669390400
transform 1 0 8288 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1492_
timestamp 1669390400
transform -1 0 17136 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _1493_
timestamp 1669390400
transform -1 0 18368 0 1 20384
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1494_
timestamp 1669390400
transform -1 0 17136 0 -1 23520
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1495_
timestamp 1669390400
transform -1 0 10976 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1496_
timestamp 1669390400
transform 1 0 10080 0 1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1497_
timestamp 1669390400
transform -1 0 14224 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1498_
timestamp 1669390400
transform 1 0 12544 0 -1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1499_
timestamp 1669390400
transform -1 0 15456 0 -1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _1500_
timestamp 1669390400
transform 1 0 8960 0 1 31360
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1501_
timestamp 1669390400
transform -1 0 14000 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1502_
timestamp 1669390400
transform -1 0 13440 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1503_
timestamp 1669390400
transform 1 0 11648 0 1 32928
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1504_
timestamp 1669390400
transform 1 0 16128 0 1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1505_
timestamp 1669390400
transform 1 0 14672 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1506_
timestamp 1669390400
transform 1 0 15568 0 -1 36064
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1507_
timestamp 1669390400
transform -1 0 16912 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1508_
timestamp 1669390400
transform 1 0 11424 0 -1 26656
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1509_
timestamp 1669390400
transform 1 0 10192 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1510_
timestamp 1669390400
transform -1 0 58240 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1511_
timestamp 1669390400
transform 1 0 3136 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1512_
timestamp 1669390400
transform -1 0 14336 0 -1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1513_
timestamp 1669390400
transform -1 0 4592 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1514_
timestamp 1669390400
transform 1 0 4144 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1515_
timestamp 1669390400
transform 1 0 5600 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1516_
timestamp 1669390400
transform 1 0 3920 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1517_
timestamp 1669390400
transform 1 0 3472 0 -1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1518_
timestamp 1669390400
transform 1 0 16240 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1519_
timestamp 1669390400
transform 1 0 15680 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1520_
timestamp 1669390400
transform 1 0 17584 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1521_
timestamp 1669390400
transform -1 0 18928 0 1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1522_
timestamp 1669390400
transform 1 0 17584 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1523_
timestamp 1669390400
transform 1 0 16576 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1524_
timestamp 1669390400
transform -1 0 8400 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1525_
timestamp 1669390400
transform 1 0 67536 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1526_
timestamp 1669390400
transform 1 0 18928 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _1527_
timestamp 1669390400
transform -1 0 20272 0 -1 20384
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1528_
timestamp 1669390400
transform -1 0 7392 0 -1 23520
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1529_
timestamp 1669390400
transform -1 0 10192 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1530_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 11312 0 1 23520
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1531_
timestamp 1669390400
transform -1 0 23744 0 1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1532_
timestamp 1669390400
transform -1 0 8512 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1533_
timestamp 1669390400
transform -1 0 7616 0 -1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1534_
timestamp 1669390400
transform 1 0 5936 0 1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1535_
timestamp 1669390400
transform -1 0 7728 0 -1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1536_
timestamp 1669390400
transform -1 0 7504 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1537_
timestamp 1669390400
transform -1 0 7280 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1538_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 8064 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1539_
timestamp 1669390400
transform 1 0 7504 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1540_
timestamp 1669390400
transform -1 0 62720 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1541_
timestamp 1669390400
transform 1 0 8624 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1542_
timestamp 1669390400
transform 1 0 2464 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1543_
timestamp 1669390400
transform -1 0 4032 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1544_
timestamp 1669390400
transform -1 0 3920 0 -1 23520
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1545_
timestamp 1669390400
transform 1 0 2352 0 -1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1546_
timestamp 1669390400
transform 1 0 2464 0 1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1547_
timestamp 1669390400
transform 1 0 3024 0 1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1548_
timestamp 1669390400
transform -1 0 7056 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1549_
timestamp 1669390400
transform 1 0 5936 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1550_
timestamp 1669390400
transform -1 0 9184 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1551_
timestamp 1669390400
transform 1 0 9072 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1552_
timestamp 1669390400
transform -1 0 12768 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1553_
timestamp 1669390400
transform 1 0 9632 0 -1 20384
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1554_
timestamp 1669390400
transform -1 0 18928 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1555_
timestamp 1669390400
transform -1 0 48720 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1556_
timestamp 1669390400
transform -1 0 20384 0 1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1557_
timestamp 1669390400
transform -1 0 17696 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1558_
timestamp 1669390400
transform 1 0 16576 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1559_
timestamp 1669390400
transform -1 0 28448 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1560_
timestamp 1669390400
transform 1 0 14448 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1561_
timestamp 1669390400
transform -1 0 19712 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _1562_
timestamp 1669390400
transform -1 0 18704 0 1 17248
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1563_
timestamp 1669390400
transform -1 0 14560 0 -1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1564_
timestamp 1669390400
transform -1 0 13776 0 -1 21952
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1565_
timestamp 1669390400
transform 1 0 2352 0 -1 28224
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _1566_
timestamp 1669390400
transform 1 0 3472 0 -1 31360
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1567_
timestamp 1669390400
transform 1 0 8512 0 1 26656
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1568_
timestamp 1669390400
transform 1 0 8512 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1569_
timestamp 1669390400
transform 1 0 9296 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1570_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 9632 0 -1 31360
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1571_
timestamp 1669390400
transform 1 0 6496 0 1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1572_
timestamp 1669390400
transform 1 0 7952 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1573_
timestamp 1669390400
transform 1 0 7168 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1574_
timestamp 1669390400
transform -1 0 10080 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1575_
timestamp 1669390400
transform 1 0 13552 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1576_
timestamp 1669390400
transform 1 0 6384 0 1 32928
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1577_
timestamp 1669390400
transform 1 0 14224 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _1578_
timestamp 1669390400
transform 1 0 19488 0 -1 34496
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _1579_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 13776 0 1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1580_
timestamp 1669390400
transform 1 0 21280 0 -1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1581_
timestamp 1669390400
transform 1 0 17360 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _1582_
timestamp 1669390400
transform 1 0 6496 0 -1 34496
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1583_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 14000 0 -1 34496
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1584_
timestamp 1669390400
transform 1 0 10864 0 1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1585_
timestamp 1669390400
transform 1 0 19376 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1586_
timestamp 1669390400
transform 1 0 22848 0 -1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1587_
timestamp 1669390400
transform 1 0 24416 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1588_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 3472 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1589_
timestamp 1669390400
transform -1 0 5712 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1590_
timestamp 1669390400
transform -1 0 28336 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1591_
timestamp 1669390400
transform 1 0 25088 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1592_
timestamp 1669390400
transform -1 0 26096 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1593_
timestamp 1669390400
transform -1 0 25312 0 1 28224
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1594_
timestamp 1669390400
transform 1 0 4480 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1595_
timestamp 1669390400
transform -1 0 6832 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1596_
timestamp 1669390400
transform 1 0 5152 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1597_
timestamp 1669390400
transform 1 0 3360 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1598_
timestamp 1669390400
transform 1 0 3472 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1599_
timestamp 1669390400
transform 1 0 4144 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1600_
timestamp 1669390400
transform -1 0 10864 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1601_
timestamp 1669390400
transform 1 0 8400 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1602_
timestamp 1669390400
transform 1 0 8176 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1603_
timestamp 1669390400
transform 1 0 9296 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1604_
timestamp 1669390400
transform -1 0 4816 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1605_
timestamp 1669390400
transform -1 0 5152 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1606_
timestamp 1669390400
transform -1 0 7504 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1607_
timestamp 1669390400
transform 1 0 3248 0 -1 21952
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1608_
timestamp 1669390400
transform 1 0 7392 0 1 21952
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1609_
timestamp 1669390400
transform 1 0 8960 0 1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1610_
timestamp 1669390400
transform -1 0 15344 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1611_
timestamp 1669390400
transform 1 0 13552 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1612_
timestamp 1669390400
transform 1 0 9632 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1613_
timestamp 1669390400
transform -1 0 14112 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1614_
timestamp 1669390400
transform 1 0 11088 0 -1 18816
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1615_
timestamp 1669390400
transform 1 0 17584 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1616_
timestamp 1669390400
transform -1 0 18592 0 1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1617_
timestamp 1669390400
transform 1 0 17584 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1618_
timestamp 1669390400
transform 1 0 16576 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1619_
timestamp 1669390400
transform -1 0 30912 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1620_
timestamp 1669390400
transform 1 0 18256 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _1621_
timestamp 1669390400
transform 1 0 17360 0 1 14112
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1622_
timestamp 1669390400
transform 1 0 21168 0 -1 17248
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1623_
timestamp 1669390400
transform -1 0 22624 0 -1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _1624_
timestamp 1669390400
transform 1 0 12768 0 -1 23520
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1625_
timestamp 1669390400
transform 1 0 14336 0 -1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1626_
timestamp 1669390400
transform 1 0 23184 0 -1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1627_
timestamp 1669390400
transform 1 0 4032 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1628_
timestamp 1669390400
transform 1 0 4256 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1629_
timestamp 1669390400
transform -1 0 6496 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1630_
timestamp 1669390400
transform 1 0 23744 0 -1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1631_
timestamp 1669390400
transform 1 0 22736 0 -1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1632_
timestamp 1669390400
transform 1 0 23184 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1633_
timestamp 1669390400
transform 1 0 25872 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1634_
timestamp 1669390400
transform 1 0 26320 0 1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1635_
timestamp 1669390400
transform 1 0 22288 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1636_
timestamp 1669390400
transform 1 0 23408 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1637_
timestamp 1669390400
transform 1 0 25648 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1638_
timestamp 1669390400
transform -1 0 30688 0 -1 36064
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1639_
timestamp 1669390400
transform -1 0 29008 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1640_
timestamp 1669390400
transform 1 0 25312 0 1 34496
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1641_
timestamp 1669390400
transform 1 0 26096 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1642_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 27216 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1643_
timestamp 1669390400
transform 1 0 26432 0 1 28224
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1644_
timestamp 1669390400
transform 1 0 14672 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1645_
timestamp 1669390400
transform -1 0 24304 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1646_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 8736 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1647_
timestamp 1669390400
transform 1 0 9632 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1648_
timestamp 1669390400
transform 1 0 9632 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1649_
timestamp 1669390400
transform 1 0 26432 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1650_
timestamp 1669390400
transform -1 0 58240 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1651_
timestamp 1669390400
transform -1 0 58240 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1652_
timestamp 1669390400
transform 1 0 27440 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1653_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 26432 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1654_
timestamp 1669390400
transform 1 0 28112 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1655_
timestamp 1669390400
transform 1 0 28448 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1656_
timestamp 1669390400
transform -1 0 28112 0 -1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1657_
timestamp 1669390400
transform 1 0 12432 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1658_
timestamp 1669390400
transform -1 0 15232 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1659_
timestamp 1669390400
transform 1 0 13552 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1660_
timestamp 1669390400
transform -1 0 6160 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1661_
timestamp 1669390400
transform -1 0 4368 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1662_
timestamp 1669390400
transform -1 0 4368 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1663_
timestamp 1669390400
transform -1 0 10192 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1664_
timestamp 1669390400
transform -1 0 10528 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1665_
timestamp 1669390400
transform -1 0 10304 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1666_
timestamp 1669390400
transform -1 0 5040 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1667_
timestamp 1669390400
transform -1 0 4032 0 1 15680
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1668_
timestamp 1669390400
transform -1 0 4144 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1669_
timestamp 1669390400
transform 1 0 2800 0 1 17248
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1670_
timestamp 1669390400
transform 1 0 4704 0 -1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1671_
timestamp 1669390400
transform 1 0 5600 0 1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1672_
timestamp 1669390400
transform 1 0 21728 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1673_
timestamp 1669390400
transform -1 0 23744 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1674_
timestamp 1669390400
transform -1 0 13776 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1675_
timestamp 1669390400
transform 1 0 13552 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1676_
timestamp 1669390400
transform 1 0 12208 0 -1 15680
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1677_
timestamp 1669390400
transform -1 0 19600 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1678_
timestamp 1669390400
transform 1 0 14784 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1679_
timestamp 1669390400
transform 1 0 17920 0 -1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1680_
timestamp 1669390400
transform 1 0 18256 0 -1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1681_
timestamp 1669390400
transform 1 0 18816 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1682_
timestamp 1669390400
transform -1 0 42336 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1683_
timestamp 1669390400
transform -1 0 66304 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1684_
timestamp 1669390400
transform 1 0 22064 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _1685_
timestamp 1669390400
transform 1 0 20608 0 -1 14112
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1686_
timestamp 1669390400
transform 1 0 23296 0 -1 15680
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1687_
timestamp 1669390400
transform 1 0 23744 0 1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _1688_
timestamp 1669390400
transform 1 0 23072 0 1 18816
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1689_
timestamp 1669390400
transform 1 0 25536 0 -1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1690_
timestamp 1669390400
transform 1 0 26432 0 1 31360
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1691_
timestamp 1669390400
transform 1 0 27104 0 -1 32928
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1692_
timestamp 1669390400
transform 1 0 29456 0 1 32928
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1693_
timestamp 1669390400
transform 1 0 24416 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1694_
timestamp 1669390400
transform 1 0 26992 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1695_
timestamp 1669390400
transform 1 0 30912 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1696_
timestamp 1669390400
transform 1 0 30912 0 1 34496
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1697_
timestamp 1669390400
transform 1 0 31696 0 -1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1698_
timestamp 1669390400
transform 1 0 33488 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1699_
timestamp 1669390400
transform 1 0 28336 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1700_
timestamp 1669390400
transform 1 0 25648 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1701_
timestamp 1669390400
transform -1 0 28000 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1702_
timestamp 1669390400
transform 1 0 4704 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1703_
timestamp 1669390400
transform 1 0 5600 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1704_
timestamp 1669390400
transform 1 0 6272 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1705_
timestamp 1669390400
transform 1 0 5600 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1706_
timestamp 1669390400
transform -1 0 68208 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1707_
timestamp 1669390400
transform 1 0 63728 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1708_
timestamp 1669390400
transform 1 0 26544 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1709_
timestamp 1669390400
transform -1 0 29008 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1710_
timestamp 1669390400
transform -1 0 28000 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1711_
timestamp 1669390400
transform 1 0 25984 0 -1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1712_
timestamp 1669390400
transform 1 0 27216 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1713_
timestamp 1669390400
transform 1 0 27216 0 -1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1714_
timestamp 1669390400
transform 1 0 29456 0 1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1715_
timestamp 1669390400
transform 1 0 30016 0 -1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1716_
timestamp 1669390400
transform -1 0 24640 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1717_
timestamp 1669390400
transform -1 0 26544 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1718_
timestamp 1669390400
transform 1 0 23968 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1719_
timestamp 1669390400
transform 1 0 2912 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1720_
timestamp 1669390400
transform 1 0 4256 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1721_
timestamp 1669390400
transform -1 0 4144 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1722_
timestamp 1669390400
transform 1 0 4368 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1723_
timestamp 1669390400
transform -1 0 12880 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1724_
timestamp 1669390400
transform 1 0 10864 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1725_
timestamp 1669390400
transform -1 0 12096 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1726_
timestamp 1669390400
transform 1 0 2128 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1727_
timestamp 1669390400
transform 1 0 2352 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1728_
timestamp 1669390400
transform 1 0 2352 0 1 10976
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1729_
timestamp 1669390400
transform 1 0 2912 0 -1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1730_
timestamp 1669390400
transform 1 0 5824 0 1 15680
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1731_
timestamp 1669390400
transform 1 0 6608 0 -1 17248
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1732_
timestamp 1669390400
transform 1 0 23744 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1733_
timestamp 1669390400
transform -1 0 25088 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1734_
timestamp 1669390400
transform -1 0 14112 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1735_
timestamp 1669390400
transform 1 0 13552 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1736_
timestamp 1669390400
transform 1 0 12432 0 -1 14112
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1737_
timestamp 1669390400
transform -1 0 20832 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1738_
timestamp 1669390400
transform -1 0 21056 0 1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1739_
timestamp 1669390400
transform -1 0 20944 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1740_
timestamp 1669390400
transform 1 0 18032 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1741_
timestamp 1669390400
transform -1 0 66192 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1742_
timestamp 1669390400
transform 1 0 64960 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1743_
timestamp 1669390400
transform 1 0 19264 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _1744_
timestamp 1669390400
transform 1 0 18368 0 1 10976
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1745_
timestamp 1669390400
transform 1 0 24640 0 1 12544
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1746_
timestamp 1669390400
transform 1 0 24976 0 1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _1747_
timestamp 1669390400
transform 1 0 25536 0 -1 17248
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1748_
timestamp 1669390400
transform 1 0 29792 0 1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1749_
timestamp 1669390400
transform 1 0 30912 0 1 31360
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _1750_
timestamp 1669390400
transform 1 0 32480 0 1 32928
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1751_
timestamp 1669390400
transform 1 0 28784 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1752_
timestamp 1669390400
transform 1 0 28112 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1753_
timestamp 1669390400
transform 1 0 34496 0 1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1754_
timestamp 1669390400
transform 1 0 31136 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1755_
timestamp 1669390400
transform -1 0 30688 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1756_
timestamp 1669390400
transform 1 0 35616 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _1757_
timestamp 1669390400
transform 1 0 36960 0 1 36064
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1758_
timestamp 1669390400
transform 1 0 39312 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1759_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 34608 0 -1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1760_
timestamp 1669390400
transform 1 0 37072 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1761_
timestamp 1669390400
transform -1 0 36960 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1762_
timestamp 1669390400
transform 1 0 37408 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1763_
timestamp 1669390400
transform -1 0 47712 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1764_
timestamp 1669390400
transform 1 0 35056 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1765_
timestamp 1669390400
transform 1 0 33040 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1766_
timestamp 1669390400
transform 1 0 33488 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1767_
timestamp 1669390400
transform 1 0 33600 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1768_
timestamp 1669390400
transform 1 0 31360 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1769_
timestamp 1669390400
transform -1 0 32480 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1770_
timestamp 1669390400
transform 1 0 31136 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1771_
timestamp 1669390400
transform 1 0 28336 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1772_
timestamp 1669390400
transform 1 0 7504 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1773_
timestamp 1669390400
transform 1 0 6720 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1774_
timestamp 1669390400
transform -1 0 66192 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1775_
timestamp 1669390400
transform 1 0 63616 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1776_
timestamp 1669390400
transform -1 0 31024 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1777_
timestamp 1669390400
transform 1 0 27328 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1778_
timestamp 1669390400
transform 1 0 29568 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1779_
timestamp 1669390400
transform -1 0 27776 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1780_
timestamp 1669390400
transform 1 0 26208 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1781_
timestamp 1669390400
transform 1 0 27440 0 -1 23520
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1782_
timestamp 1669390400
transform 1 0 30240 0 -1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1783_
timestamp 1669390400
transform 1 0 31248 0 -1 28224
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1784_
timestamp 1669390400
transform -1 0 33264 0 1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1785_
timestamp 1669390400
transform 1 0 31584 0 -1 29792
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1786_
timestamp 1669390400
transform -1 0 26656 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1787_
timestamp 1669390400
transform -1 0 27440 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1788_
timestamp 1669390400
transform 1 0 26096 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1789_
timestamp 1669390400
transform -1 0 4816 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1790_
timestamp 1669390400
transform 1 0 3248 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1791_
timestamp 1669390400
transform -1 0 14896 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1792_
timestamp 1669390400
transform 1 0 11312 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1793_
timestamp 1669390400
transform -1 0 13104 0 1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1794_
timestamp 1669390400
transform 1 0 3136 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1795_
timestamp 1669390400
transform -1 0 8736 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1796_
timestamp 1669390400
transform 1 0 3696 0 -1 12544
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1797_
timestamp 1669390400
transform 1 0 7392 0 -1 14112
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1798_
timestamp 1669390400
transform 1 0 7616 0 1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1799_
timestamp 1669390400
transform 1 0 24528 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1800_
timestamp 1669390400
transform -1 0 26432 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1801_
timestamp 1669390400
transform 1 0 12208 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1802_
timestamp 1669390400
transform -1 0 15456 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1803_
timestamp 1669390400
transform 1 0 12992 0 -1 12544
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1804_
timestamp 1669390400
transform 1 0 21056 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1805_
timestamp 1669390400
transform 1 0 20944 0 -1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1806_
timestamp 1669390400
transform 1 0 21504 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1807_
timestamp 1669390400
transform 1 0 17136 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1808_
timestamp 1669390400
transform 1 0 29792 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1809_
timestamp 1669390400
transform -1 0 18816 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1810_
timestamp 1669390400
transform 1 0 22736 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _1811_
timestamp 1669390400
transform 1 0 21840 0 -1 10976
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1812_
timestamp 1669390400
transform 1 0 24528 0 1 10976
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1813_
timestamp 1669390400
transform 1 0 25536 0 -1 12544
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _1814_
timestamp 1669390400
transform 1 0 27776 0 -1 14112
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1815_
timestamp 1669390400
transform 1 0 34720 0 -1 31360
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _1816_
timestamp 1669390400
transform 1 0 37632 0 1 32928
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1817_
timestamp 1669390400
transform 1 0 39312 0 1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1818_
timestamp 1669390400
transform 1 0 41440 0 -1 36064
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1819_
timestamp 1669390400
transform 1 0 47600 0 -1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1820_
timestamp 1669390400
transform 1 0 50736 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1821_
timestamp 1669390400
transform 1 0 41216 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1822_
timestamp 1669390400
transform -1 0 45696 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1823_
timestamp 1669390400
transform 1 0 40208 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1824_
timestamp 1669390400
transform 1 0 33488 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1825_
timestamp 1669390400
transform 1 0 32592 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1826_
timestamp 1669390400
transform 1 0 33488 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1827_
timestamp 1669390400
transform 1 0 34272 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1828_
timestamp 1669390400
transform -1 0 36848 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1829_
timestamp 1669390400
transform 1 0 35168 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1830_
timestamp 1669390400
transform 1 0 27552 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1831_
timestamp 1669390400
transform -1 0 29008 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1832_
timestamp 1669390400
transform 1 0 27888 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1833_
timestamp 1669390400
transform -1 0 5152 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1834_
timestamp 1669390400
transform -1 0 4816 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1835_
timestamp 1669390400
transform -1 0 6272 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1836_
timestamp 1669390400
transform -1 0 4928 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1837_
timestamp 1669390400
transform 1 0 12320 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1838_
timestamp 1669390400
transform -1 0 14112 0 -1 10976
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1839_
timestamp 1669390400
transform 1 0 13552 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1840_
timestamp 1669390400
transform -1 0 8400 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1841_
timestamp 1669390400
transform -1 0 9184 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _1842_
timestamp 1669390400
transform 1 0 5376 0 -1 10976
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1843_
timestamp 1669390400
transform 1 0 7952 0 1 10976
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1844_
timestamp 1669390400
transform 1 0 9632 0 -1 12544
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1845_
timestamp 1669390400
transform 1 0 25536 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1846_
timestamp 1669390400
transform -1 0 27104 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1847_
timestamp 1669390400
transform 1 0 13552 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1848_
timestamp 1669390400
transform -1 0 15120 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1849_
timestamp 1669390400
transform 1 0 13552 0 1 7840
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1850_
timestamp 1669390400
transform 1 0 17024 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1851_
timestamp 1669390400
transform 1 0 18032 0 -1 10976
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1852_
timestamp 1669390400
transform -1 0 19040 0 1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1853_
timestamp 1669390400
transform -1 0 18816 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1854_
timestamp 1669390400
transform 1 0 63728 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1855_
timestamp 1669390400
transform 1 0 59024 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1856_
timestamp 1669390400
transform -1 0 25424 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _1857_
timestamp 1669390400
transform 1 0 17024 0 1 6272
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1858_
timestamp 1669390400
transform 1 0 17808 0 1 7840
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1859_
timestamp 1669390400
transform 1 0 18032 0 -1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _1860_
timestamp 1669390400
transform 1 0 28336 0 -1 12544
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1861_
timestamp 1669390400
transform 1 0 35952 0 -1 28224
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1862_
timestamp 1669390400
transform -1 0 32144 0 1 26656
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1863_
timestamp 1669390400
transform -1 0 32704 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1864_
timestamp 1669390400
transform 1 0 6944 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1865_
timestamp 1669390400
transform 1 0 9632 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1866_
timestamp 1669390400
transform 1 0 9184 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1867_
timestamp 1669390400
transform 1 0 64848 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1868_
timestamp 1669390400
transform -1 0 64848 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1869_
timestamp 1669390400
transform -1 0 40544 0 1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1870_
timestamp 1669390400
transform 1 0 39648 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1871_
timestamp 1669390400
transform -1 0 39424 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1872_
timestamp 1669390400
transform -1 0 38864 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1873_
timestamp 1669390400
transform 1 0 26320 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1874_
timestamp 1669390400
transform 1 0 26320 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1875_
timestamp 1669390400
transform 1 0 25312 0 1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1876_
timestamp 1669390400
transform -1 0 27664 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1877_
timestamp 1669390400
transform -1 0 27888 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1878_
timestamp 1669390400
transform 1 0 27328 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _1879_
timestamp 1669390400
transform 1 0 27216 0 -1 21952
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1880_
timestamp 1669390400
transform 1 0 29792 0 -1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1881_
timestamp 1669390400
transform 1 0 33600 0 1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1882_
timestamp 1669390400
transform 1 0 34272 0 -1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1883_
timestamp 1669390400
transform 1 0 35168 0 1 26656
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1884_
timestamp 1669390400
transform 1 0 36736 0 -1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _1885_
timestamp 1669390400
transform 1 0 39312 0 1 31360
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1886_
timestamp 1669390400
transform 1 0 42112 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1887_
timestamp 1669390400
transform 1 0 37408 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1888_
timestamp 1669390400
transform 1 0 36960 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1889_
timestamp 1669390400
transform -1 0 38976 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1890_
timestamp 1669390400
transform 1 0 42336 0 1 34496
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1891_
timestamp 1669390400
transform -1 0 46928 0 -1 36064
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1892_
timestamp 1669390400
transform -1 0 44352 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1893_
timestamp 1669390400
transform 1 0 42448 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1894_
timestamp 1669390400
transform 1 0 38976 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1895_
timestamp 1669390400
transform 1 0 40096 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1896_
timestamp 1669390400
transform -1 0 42336 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1897_
timestamp 1669390400
transform 1 0 35840 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1898_
timestamp 1669390400
transform -1 0 34944 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1899_
timestamp 1669390400
transform 1 0 39648 0 -1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1900_
timestamp 1669390400
transform 1 0 36400 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1901_
timestamp 1669390400
transform -1 0 38304 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1902_
timestamp 1669390400
transform 1 0 30128 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1903_
timestamp 1669390400
transform -1 0 33376 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1904_
timestamp 1669390400
transform -1 0 33040 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1905_
timestamp 1669390400
transform 1 0 8512 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1906_
timestamp 1669390400
transform -1 0 9184 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1907_
timestamp 1669390400
transform -1 0 69664 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1908_
timestamp 1669390400
transform -1 0 40768 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1909_
timestamp 1669390400
transform 1 0 39872 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1910_
timestamp 1669390400
transform 1 0 40208 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1911_
timestamp 1669390400
transform -1 0 41328 0 1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1912_
timestamp 1669390400
transform -1 0 39984 0 -1 23520
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1913_
timestamp 1669390400
transform -1 0 28560 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1914_
timestamp 1669390400
transform 1 0 25536 0 -1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1915_
timestamp 1669390400
transform 1 0 27104 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1916_
timestamp 1669390400
transform 1 0 29456 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1917_
timestamp 1669390400
transform 1 0 31248 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1918_
timestamp 1669390400
transform 1 0 29904 0 1 20384
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1919_
timestamp 1669390400
transform 1 0 31808 0 1 21952
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1920_
timestamp 1669390400
transform 1 0 33488 0 -1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1921_
timestamp 1669390400
transform 1 0 32928 0 1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1922_
timestamp 1669390400
transform 1 0 33488 0 -1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1923_
timestamp 1669390400
transform 1 0 27440 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1924_
timestamp 1669390400
transform 1 0 29456 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1925_
timestamp 1669390400
transform 1 0 29456 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1926_
timestamp 1669390400
transform -1 0 10304 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1927_
timestamp 1669390400
transform 1 0 4256 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1928_
timestamp 1669390400
transform 1 0 7504 0 1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1929_
timestamp 1669390400
transform -1 0 16800 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1930_
timestamp 1669390400
transform 1 0 13104 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1931_
timestamp 1669390400
transform -1 0 14336 0 -1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1932_
timestamp 1669390400
transform -1 0 6048 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1933_
timestamp 1669390400
transform -1 0 9856 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1934_
timestamp 1669390400
transform -1 0 9184 0 -1 7840
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1935_
timestamp 1669390400
transform 1 0 3696 0 1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1936_
timestamp 1669390400
transform 1 0 10080 0 -1 9408
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1937_
timestamp 1669390400
transform 1 0 10528 0 1 9408
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1938_
timestamp 1669390400
transform 1 0 19040 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1939_
timestamp 1669390400
transform -1 0 20384 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1940_
timestamp 1669390400
transform 1 0 12432 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1941_
timestamp 1669390400
transform -1 0 16352 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1942_
timestamp 1669390400
transform 1 0 12320 0 -1 6272
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1943_
timestamp 1669390400
transform -1 0 24304 0 -1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1944_
timestamp 1669390400
transform -1 0 24528 0 1 6272
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1945_
timestamp 1669390400
transform 1 0 22736 0 -1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1946_
timestamp 1669390400
transform -1 0 25088 0 -1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1947_
timestamp 1669390400
transform -1 0 55776 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1948_
timestamp 1669390400
transform -1 0 40656 0 -1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _1949_
timestamp 1669390400
transform 1 0 23520 0 1 4704
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1950_
timestamp 1669390400
transform -1 0 22960 0 1 4704
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1951_
timestamp 1669390400
transform 1 0 21504 0 1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1952_
timestamp 1669390400
transform 1 0 23072 0 -1 9408
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1953_
timestamp 1669390400
transform 1 0 25760 0 1 9408
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1954_
timestamp 1669390400
transform 1 0 37408 0 1 12544
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1955_
timestamp 1669390400
transform 1 0 36624 0 -1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _1956_
timestamp 1669390400
transform 1 0 41440 0 -1 29792
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1957_
timestamp 1669390400
transform 1 0 42896 0 1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1958_
timestamp 1669390400
transform 1 0 43568 0 1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1959_
timestamp 1669390400
transform 1 0 47936 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1960_
timestamp 1669390400
transform 1 0 42112 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1961_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 44128 0 -1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1962_
timestamp 1669390400
transform 1 0 49616 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1963_
timestamp 1669390400
transform 1 0 50960 0 -1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1964_
timestamp 1669390400
transform 1 0 52640 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1965_
timestamp 1669390400
transform 1 0 45360 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1966_
timestamp 1669390400
transform 1 0 52304 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1967_
timestamp 1669390400
transform -1 0 52080 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1968_
timestamp 1669390400
transform 1 0 41440 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1969_
timestamp 1669390400
transform 1 0 43456 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1970_
timestamp 1669390400
transform 1 0 38976 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1971_
timestamp 1669390400
transform -1 0 41328 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1972_
timestamp 1669390400
transform 1 0 40096 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1973_
timestamp 1669390400
transform 1 0 68768 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1974_
timestamp 1669390400
transform -1 0 44128 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1975_
timestamp 1669390400
transform 1 0 34496 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1976_
timestamp 1669390400
transform 1 0 35168 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1977_
timestamp 1669390400
transform 1 0 35280 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1978_
timestamp 1669390400
transform 1 0 41440 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1979_
timestamp 1669390400
transform 1 0 39984 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1980_
timestamp 1669390400
transform 1 0 40880 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1981_
timestamp 1669390400
transform 1 0 42224 0 -1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1982_
timestamp 1669390400
transform -1 0 44576 0 1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1983_
timestamp 1669390400
transform 1 0 36400 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1984_
timestamp 1669390400
transform -1 0 38416 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1985_
timestamp 1669390400
transform 1 0 31808 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1986_
timestamp 1669390400
transform 1 0 32480 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1987_
timestamp 1669390400
transform -1 0 34272 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1988_
timestamp 1669390400
transform 1 0 10304 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1989_
timestamp 1669390400
transform 1 0 11760 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1990_
timestamp 1669390400
transform 1 0 10976 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1991_
timestamp 1669390400
transform -1 0 40096 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1992_
timestamp 1669390400
transform -1 0 41888 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1993_
timestamp 1669390400
transform -1 0 40992 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1994_
timestamp 1669390400
transform 1 0 38528 0 1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1995_
timestamp 1669390400
transform -1 0 42336 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1996_
timestamp 1669390400
transform -1 0 41216 0 1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1997_
timestamp 1669390400
transform 1 0 29456 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1998_
timestamp 1669390400
transform 1 0 30128 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1999_
timestamp 1669390400
transform 1 0 30240 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2000_
timestamp 1669390400
transform 1 0 27552 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2001_
timestamp 1669390400
transform 1 0 30016 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2002_
timestamp 1669390400
transform 1 0 29120 0 -1 18816
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2003_
timestamp 1669390400
transform 1 0 33600 0 1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2004_
timestamp 1669390400
transform -1 0 36512 0 1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2005_
timestamp 1669390400
transform 1 0 34832 0 -1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2006_
timestamp 1669390400
transform 1 0 35392 0 1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2007_
timestamp 1669390400
transform 1 0 23520 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2008_
timestamp 1669390400
transform -1 0 26544 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2009_
timestamp 1669390400
transform 1 0 9632 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2010_
timestamp 1669390400
transform 1 0 4144 0 -1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2011_
timestamp 1669390400
transform 1 0 18368 0 1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2012_
timestamp 1669390400
transform -1 0 14448 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2013_
timestamp 1669390400
transform 1 0 13552 0 1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2014_
timestamp 1669390400
transform -1 0 8960 0 1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2015_
timestamp 1669390400
transform -1 0 10640 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2016_
timestamp 1669390400
transform -1 0 7168 0 -1 6272
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2017_
timestamp 1669390400
transform 1 0 2800 0 -1 6272
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2018_
timestamp 1669390400
transform 1 0 3472 0 -1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2019_
timestamp 1669390400
transform 1 0 21840 0 -1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2020_
timestamp 1669390400
transform -1 0 22400 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2021_
timestamp 1669390400
transform -1 0 35840 0 -1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2022_
timestamp 1669390400
transform -1 0 16800 0 1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2023_
timestamp 1669390400
transform 1 0 14112 0 -1 4704
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2024_
timestamp 1669390400
transform 1 0 42672 0 1 3136
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2025_
timestamp 1669390400
transform 1 0 53536 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2026_
timestamp 1669390400
transform -1 0 27888 0 -1 4704
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2027_
timestamp 1669390400
transform 1 0 25536 0 -1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2028_
timestamp 1669390400
transform -1 0 40432 0 1 3136
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2029_
timestamp 1669390400
transform -1 0 54656 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2030_
timestamp 1669390400
transform -1 0 31024 0 1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2031_
timestamp 1669390400
transform -1 0 30912 0 -1 4704
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2032_
timestamp 1669390400
transform -1 0 20832 0 -1 4704
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2033_
timestamp 1669390400
transform 1 0 19376 0 1 3136
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2034_
timestamp 1669390400
transform 1 0 21952 0 -1 7840
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2035_
timestamp 1669390400
transform 1 0 23072 0 1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2036_
timestamp 1669390400
transform 1 0 28672 0 -1 10976
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2037_
timestamp 1669390400
transform 1 0 37408 0 1 21952
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2038_
timestamp 1669390400
transform 1 0 38192 0 -1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2039_
timestamp 1669390400
transform 1 0 39088 0 -1 26656
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2040_
timestamp 1669390400
transform 1 0 44800 0 -1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2041_
timestamp 1669390400
transform 1 0 45808 0 -1 32928
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2042_
timestamp 1669390400
transform 1 0 49952 0 -1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2043_
timestamp 1669390400
transform 1 0 51632 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2044_
timestamp 1669390400
transform 1 0 41776 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2045_
timestamp 1669390400
transform 1 0 59920 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2046_
timestamp 1669390400
transform 1 0 43904 0 -1 25088
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2047_
timestamp 1669390400
transform 1 0 45360 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2048_
timestamp 1669390400
transform 1 0 38640 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2049_
timestamp 1669390400
transform -1 0 42336 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2050_
timestamp 1669390400
transform 1 0 34272 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2051_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 37072 0 -1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2052_
timestamp 1669390400
transform 1 0 41440 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2053_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 41552 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2054_
timestamp 1669390400
transform -1 0 46816 0 1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2055_
timestamp 1669390400
transform 1 0 29456 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2056_
timestamp 1669390400
transform -1 0 38192 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2057_
timestamp 1669390400
transform 1 0 34160 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2058_
timestamp 1669390400
transform 1 0 34384 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2059_
timestamp 1669390400
transform -1 0 36064 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2060_
timestamp 1669390400
transform -1 0 6608 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2061_
timestamp 1669390400
transform 1 0 4256 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2062_
timestamp 1669390400
transform -1 0 5936 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2063_
timestamp 1669390400
transform 1 0 39424 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2064_
timestamp 1669390400
transform 1 0 40432 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2065_
timestamp 1669390400
transform -1 0 43120 0 -1 18816
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2066_
timestamp 1669390400
transform -1 0 40992 0 -1 18816
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2067_
timestamp 1669390400
transform 1 0 30016 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2068_
timestamp 1669390400
transform 1 0 31920 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _2069_
timestamp 1669390400
transform -1 0 32928 0 1 17248
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2070_
timestamp 1669390400
transform -1 0 35504 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2071_
timestamp 1669390400
transform -1 0 33040 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2072_
timestamp 1669390400
transform 1 0 30800 0 -1 17248
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2073_
timestamp 1669390400
transform 1 0 31472 0 1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2074_
timestamp 1669390400
transform 1 0 31696 0 1 14112
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2075_
timestamp 1669390400
transform 1 0 31920 0 1 12544
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2076_
timestamp 1669390400
transform -1 0 24192 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2077_
timestamp 1669390400
transform -1 0 22848 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2078_
timestamp 1669390400
transform -1 0 57120 0 1 3136
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2079_
timestamp 1669390400
transform 1 0 8288 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2080_
timestamp 1669390400
transform 1 0 9632 0 -1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2081_
timestamp 1669390400
transform 1 0 29568 0 1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2082_
timestamp 1669390400
transform 1 0 14784 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2083_
timestamp 1669390400
transform -1 0 15904 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2084_
timestamp 1669390400
transform 1 0 26656 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2085_
timestamp 1669390400
transform 1 0 26768 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2086_
timestamp 1669390400
transform -1 0 29232 0 -1 6272
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2087_
timestamp 1669390400
transform -1 0 11872 0 -1 4704
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2088_
timestamp 1669390400
transform 1 0 10192 0 1 4704
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2089_
timestamp 1669390400
transform -1 0 21616 0 -1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2090_
timestamp 1669390400
transform 1 0 19712 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2091_
timestamp 1669390400
transform -1 0 54992 0 1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2092_
timestamp 1669390400
transform 1 0 36064 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2093_
timestamp 1669390400
transform 1 0 34384 0 1 4704
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2094_
timestamp 1669390400
transform -1 0 46704 0 1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2095_
timestamp 1669390400
transform -1 0 42448 0 -1 4704
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2096_
timestamp 1669390400
transform 1 0 39648 0 1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2097_
timestamp 1669390400
transform 1 0 47264 0 -1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2098_
timestamp 1669390400
transform -1 0 51072 0 -1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2099_
timestamp 1669390400
transform 1 0 47264 0 1 4704
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2100_
timestamp 1669390400
transform -1 0 39872 0 -1 4704
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2101_
timestamp 1669390400
transform -1 0 37408 0 -1 4704
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2102_
timestamp 1669390400
transform -1 0 34944 0 -1 4704
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2103_
timestamp 1669390400
transform 1 0 31696 0 -1 4704
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2104_
timestamp 1669390400
transform 1 0 33488 0 -1 10976
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2105_
timestamp 1669390400
transform 1 0 33600 0 -1 12544
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2106_
timestamp 1669390400
transform 1 0 43456 0 1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2107_
timestamp 1669390400
transform 1 0 43568 0 1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2108_
timestamp 1669390400
transform 1 0 43568 0 1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2109_
timestamp 1669390400
transform 1 0 44240 0 -1 28224
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2110_
timestamp 1669390400
transform -1 0 48048 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2111_
timestamp 1669390400
transform 1 0 44240 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2112_
timestamp 1669390400
transform 1 0 45920 0 1 29792
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2113_
timestamp 1669390400
transform 1 0 48048 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2114_
timestamp 1669390400
transform 1 0 48160 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2115_
timestamp 1669390400
transform -1 0 51632 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2116_
timestamp 1669390400
transform -1 0 51184 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2117_
timestamp 1669390400
transform 1 0 45808 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2118_
timestamp 1669390400
transform -1 0 47824 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2119_
timestamp 1669390400
transform -1 0 47040 0 1 31360
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2120_
timestamp 1669390400
transform -1 0 50288 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2121_
timestamp 1669390400
transform 1 0 49392 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2122_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 48048 0 1 32928
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2123_
timestamp 1669390400
transform 1 0 49616 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2124_
timestamp 1669390400
transform -1 0 50960 0 1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2125_
timestamp 1669390400
transform -1 0 48944 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2126_
timestamp 1669390400
transform 1 0 44352 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2127_
timestamp 1669390400
transform -1 0 46816 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2128_
timestamp 1669390400
transform -1 0 48384 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2129_
timestamp 1669390400
transform 1 0 44016 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2130_
timestamp 1669390400
transform 1 0 44688 0 -1 23520
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2131_
timestamp 1669390400
transform 1 0 35616 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2132_
timestamp 1669390400
transform 1 0 34608 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2133_
timestamp 1669390400
transform -1 0 35392 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2134_
timestamp 1669390400
transform 1 0 43344 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2135_
timestamp 1669390400
transform 1 0 42224 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2136_
timestamp 1669390400
transform 1 0 43456 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2137_
timestamp 1669390400
transform 1 0 43792 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2138_
timestamp 1669390400
transform 1 0 46032 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2139_
timestamp 1669390400
transform -1 0 44912 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2140_
timestamp 1669390400
transform 1 0 33040 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2141_
timestamp 1669390400
transform -1 0 34608 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2142_
timestamp 1669390400
transform 1 0 33376 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2143_
timestamp 1669390400
transform 1 0 34272 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2144_
timestamp 1669390400
transform 1 0 34048 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2145_
timestamp 1669390400
transform 1 0 9744 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2146_
timestamp 1669390400
transform -1 0 12320 0 1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2147_
timestamp 1669390400
transform 1 0 11312 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2148_
timestamp 1669390400
transform 1 0 63952 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2149_
timestamp 1669390400
transform 1 0 38304 0 -1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2150_
timestamp 1669390400
transform 1 0 40096 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2151_
timestamp 1669390400
transform -1 0 42224 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2152_
timestamp 1669390400
transform -1 0 39872 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2153_
timestamp 1669390400
transform 1 0 30688 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2154_
timestamp 1669390400
transform -1 0 32592 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2155_
timestamp 1669390400
transform 1 0 36288 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2156_
timestamp 1669390400
transform -1 0 35616 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2157_
timestamp 1669390400
transform 1 0 34608 0 -1 17248
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2158_
timestamp 1669390400
transform 1 0 37408 0 1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2159_
timestamp 1669390400
transform 1 0 37968 0 1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2160_
timestamp 1669390400
transform -1 0 39424 0 -1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2161_
timestamp 1669390400
transform 1 0 37968 0 1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2162_
timestamp 1669390400
transform 1 0 38416 0 -1 14112
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2163_
timestamp 1669390400
transform -1 0 34496 0 1 3136
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2164_
timestamp 1669390400
transform 1 0 32704 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2165_
timestamp 1669390400
transform -1 0 29232 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2166_
timestamp 1669390400
transform -1 0 28448 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2167_
timestamp 1669390400
transform 1 0 27440 0 1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2168_
timestamp 1669390400
transform 1 0 35952 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2169_
timestamp 1669390400
transform 1 0 34720 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2170_
timestamp 1669390400
transform -1 0 35728 0 1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2171_
timestamp 1669390400
transform -1 0 33040 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2172_
timestamp 1669390400
transform 1 0 28560 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2173_
timestamp 1669390400
transform 1 0 27552 0 1 7840
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2174_
timestamp 1669390400
transform 1 0 31136 0 1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2175_
timestamp 1669390400
transform 1 0 31584 0 1 6272
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2176_
timestamp 1669390400
transform 1 0 31584 0 -1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2177_
timestamp 1669390400
transform 1 0 37632 0 -1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2178_
timestamp 1669390400
transform -1 0 39424 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2179_
timestamp 1669390400
transform 1 0 34720 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2180_
timestamp 1669390400
transform 1 0 35504 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2181_
timestamp 1669390400
transform 1 0 36064 0 -1 7840
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2182_
timestamp 1669390400
transform -1 0 51856 0 -1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2183_
timestamp 1669390400
transform -1 0 53200 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2184_
timestamp 1669390400
transform -1 0 44912 0 1 4704
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2185_
timestamp 1669390400
transform 1 0 44800 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2186_
timestamp 1669390400
transform -1 0 48944 0 -1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2187_
timestamp 1669390400
transform 1 0 51184 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2188_
timestamp 1669390400
transform -1 0 52864 0 1 4704
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2189_
timestamp 1669390400
transform -1 0 45360 0 -1 6272
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2190_
timestamp 1669390400
transform -1 0 43792 0 1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2191_
timestamp 1669390400
transform -1 0 40768 0 1 6272
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2192_
timestamp 1669390400
transform -1 0 40320 0 -1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2193_
timestamp 1669390400
transform 1 0 38864 0 -1 12544
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2194_
timestamp 1669390400
transform 1 0 39648 0 1 12544
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2195_
timestamp 1669390400
transform 1 0 43120 0 1 12544
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2196_
timestamp 1669390400
transform 1 0 45360 0 1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2197_
timestamp 1669390400
transform -1 0 48944 0 -1 25088
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2198_
timestamp 1669390400
transform 1 0 49392 0 -1 28224
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2199_
timestamp 1669390400
transform -1 0 50736 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2200_
timestamp 1669390400
transform -1 0 50848 0 -1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2201_
timestamp 1669390400
transform -1 0 47040 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2202_
timestamp 1669390400
transform 1 0 42336 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2203_
timestamp 1669390400
transform -1 0 45808 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2204_
timestamp 1669390400
transform -1 0 38192 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2205_
timestamp 1669390400
transform -1 0 40880 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2206_
timestamp 1669390400
transform -1 0 40096 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2207_
timestamp 1669390400
transform 1 0 45360 0 1 17248
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2208_
timestamp 1669390400
transform 1 0 39536 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2209_
timestamp 1669390400
transform -1 0 40992 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2210_
timestamp 1669390400
transform 1 0 39536 0 1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2211_
timestamp 1669390400
transform 1 0 30912 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2212_
timestamp 1669390400
transform 1 0 31360 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2213_
timestamp 1669390400
transform -1 0 33040 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2214_
timestamp 1669390400
transform 1 0 36400 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _2215_
timestamp 1669390400
transform -1 0 38416 0 -1 17248
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2216_
timestamp 1669390400
transform 1 0 51184 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _2217_
timestamp 1669390400
transform 1 0 49392 0 -1 17248
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2218_
timestamp 1669390400
transform -1 0 52080 0 -1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2219_
timestamp 1669390400
transform 1 0 51184 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2220_
timestamp 1669390400
transform -1 0 52304 0 -1 17248
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2221_
timestamp 1669390400
transform 1 0 41664 0 -1 17248
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2222_
timestamp 1669390400
transform 1 0 42000 0 1 14112
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2223_
timestamp 1669390400
transform -1 0 41552 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2224_
timestamp 1669390400
transform 1 0 39760 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2225_
timestamp 1669390400
transform 1 0 30352 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2226_
timestamp 1669390400
transform -1 0 32256 0 -1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2227_
timestamp 1669390400
transform 1 0 36288 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2228_
timestamp 1669390400
transform 1 0 36064 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2229_
timestamp 1669390400
transform 1 0 37408 0 1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2230_
timestamp 1669390400
transform 1 0 35392 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2231_
timestamp 1669390400
transform 1 0 30352 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2232_
timestamp 1669390400
transform 1 0 31136 0 -1 10976
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2233_
timestamp 1669390400
transform 1 0 35168 0 -1 10976
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2234_
timestamp 1669390400
transform 1 0 37968 0 -1 10976
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2235_
timestamp 1669390400
transform 1 0 39648 0 -1 10976
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2236_
timestamp 1669390400
transform -1 0 45920 0 1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2237_
timestamp 1669390400
transform 1 0 44128 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2238_
timestamp 1669390400
transform 1 0 40432 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2239_
timestamp 1669390400
transform 1 0 36288 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2240_
timestamp 1669390400
transform 1 0 41104 0 1 7840
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2241_
timestamp 1669390400
transform -1 0 49952 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2242_
timestamp 1669390400
transform 1 0 45584 0 -1 6272
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2243_
timestamp 1669390400
transform 1 0 47824 0 -1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2244_
timestamp 1669390400
transform 1 0 49840 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2245_
timestamp 1669390400
transform -1 0 53872 0 1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2246_
timestamp 1669390400
transform 1 0 49392 0 -1 7840
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2247_
timestamp 1669390400
transform -1 0 47824 0 -1 7840
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2248_
timestamp 1669390400
transform -1 0 47040 0 1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2249_
timestamp 1669390400
transform -1 0 46816 0 1 9408
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2250_
timestamp 1669390400
transform 1 0 43232 0 -1 10976
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2251_
timestamp 1669390400
transform 1 0 43456 0 -1 12544
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2252_
timestamp 1669390400
transform 1 0 44240 0 -1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2253_
timestamp 1669390400
transform 1 0 45584 0 1 14112
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2254_
timestamp 1669390400
transform 1 0 46480 0 -1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2255_
timestamp 1669390400
transform 1 0 47936 0 1 20384
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2256_
timestamp 1669390400
transform 1 0 46816 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2257_
timestamp 1669390400
transform 1 0 47600 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _2258_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 49840 0 1 21952
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2259_
timestamp 1669390400
transform 1 0 52080 0 -1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2260_
timestamp 1669390400
transform 1 0 47264 0 1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2261_
timestamp 1669390400
transform 1 0 48048 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2262_
timestamp 1669390400
transform 1 0 49392 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2263_
timestamp 1669390400
transform 1 0 45360 0 1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai33_1  _2264_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 47936 0 1 26656
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2265_
timestamp 1669390400
transform 1 0 46144 0 1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2266_
timestamp 1669390400
transform 1 0 52192 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2267_
timestamp 1669390400
transform 1 0 54208 0 -1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2268_
timestamp 1669390400
transform -1 0 55104 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2269_
timestamp 1669390400
transform -1 0 54656 0 1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2270_
timestamp 1669390400
transform -1 0 52864 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2271_
timestamp 1669390400
transform 1 0 48272 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2272_
timestamp 1669390400
transform 1 0 48384 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2273_
timestamp 1669390400
transform -1 0 50288 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2274_
timestamp 1669390400
transform 1 0 45360 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2275_
timestamp 1669390400
transform 1 0 46032 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2276_
timestamp 1669390400
transform -1 0 47936 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2277_
timestamp 1669390400
transform -1 0 43568 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2278_
timestamp 1669390400
transform -1 0 44352 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2279_
timestamp 1669390400
transform 1 0 43008 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2280_
timestamp 1669390400
transform 1 0 44016 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2281_
timestamp 1669390400
transform -1 0 46256 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2282_
timestamp 1669390400
transform -1 0 47264 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2283_
timestamp 1669390400
transform -1 0 46480 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2284_
timestamp 1669390400
transform 1 0 46032 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2285_
timestamp 1669390400
transform 1 0 46032 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2286_
timestamp 1669390400
transform -1 0 40768 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2287_
timestamp 1669390400
transform 1 0 38416 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2288_
timestamp 1669390400
transform -1 0 40320 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2289_
timestamp 1669390400
transform 1 0 50400 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2290_
timestamp 1669390400
transform 1 0 47488 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2291_
timestamp 1669390400
transform 1 0 54096 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2292_
timestamp 1669390400
transform 1 0 52080 0 -1 15680
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2293_
timestamp 1669390400
transform 1 0 52528 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2294_
timestamp 1669390400
transform -1 0 52640 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2295_
timestamp 1669390400
transform 1 0 53312 0 1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2296_
timestamp 1669390400
transform 1 0 53312 0 1 12544
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2297_
timestamp 1669390400
transform -1 0 54768 0 -1 12544
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2298_
timestamp 1669390400
transform -1 0 44912 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2299_
timestamp 1669390400
transform -1 0 45696 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2300_
timestamp 1669390400
transform -1 0 57680 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2301_
timestamp 1669390400
transform -1 0 43680 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2302_
timestamp 1669390400
transform 1 0 35392 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2303_
timestamp 1669390400
transform 1 0 42336 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2304_
timestamp 1669390400
transform 1 0 37072 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2305_
timestamp 1669390400
transform 1 0 40992 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2306_
timestamp 1669390400
transform 1 0 41440 0 -1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2307_
timestamp 1669390400
transform 1 0 56336 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2308_
timestamp 1669390400
transform -1 0 69328 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2309_
timestamp 1669390400
transform 1 0 56336 0 1 9408
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2310_
timestamp 1669390400
transform -1 0 57568 0 1 10976
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2311_
timestamp 1669390400
transform -1 0 54768 0 1 10976
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2312_
timestamp 1669390400
transform -1 0 52864 0 1 10976
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2313_
timestamp 1669390400
transform -1 0 48608 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2314_
timestamp 1669390400
transform 1 0 47264 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2315_
timestamp 1669390400
transform 1 0 50736 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2316_
timestamp 1669390400
transform 1 0 42784 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2317_
timestamp 1669390400
transform 1 0 50400 0 -1 9408
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2318_
timestamp 1669390400
transform -1 0 52080 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2319_
timestamp 1669390400
transform -1 0 56672 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2320_
timestamp 1669390400
transform -1 0 56896 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2321_
timestamp 1669390400
transform 1 0 49728 0 -1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2322_
timestamp 1669390400
transform 1 0 50736 0 1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2323_
timestamp 1669390400
transform 1 0 54432 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2324_
timestamp 1669390400
transform 1 0 56560 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2325_
timestamp 1669390400
transform 1 0 54208 0 -1 7840
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2326_
timestamp 1669390400
transform -1 0 56112 0 1 7840
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2327_
timestamp 1669390400
transform -1 0 55552 0 -1 9408
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2328_
timestamp 1669390400
transform 1 0 46256 0 -1 10976
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2329_
timestamp 1669390400
transform 1 0 49392 0 -1 12544
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2330_
timestamp 1669390400
transform -1 0 50176 0 1 12544
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2331_
timestamp 1669390400
transform -1 0 50736 0 -1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2332_
timestamp 1669390400
transform 1 0 48272 0 1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2333_
timestamp 1669390400
transform 1 0 47824 0 1 18816
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2334_
timestamp 1669390400
transform 1 0 51744 0 -1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2335_
timestamp 1669390400
transform 1 0 52304 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2336_
timestamp 1669390400
transform -1 0 54208 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2337_
timestamp 1669390400
transform -1 0 53872 0 -1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2338_
timestamp 1669390400
transform -1 0 50960 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2339_
timestamp 1669390400
transform -1 0 48944 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2340_
timestamp 1669390400
transform 1 0 49840 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2341_
timestamp 1669390400
transform 1 0 50624 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2342_
timestamp 1669390400
transform -1 0 55440 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2343_
timestamp 1669390400
transform 1 0 54992 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2344_
timestamp 1669390400
transform 1 0 54768 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2345_
timestamp 1669390400
transform 1 0 48384 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2346_
timestamp 1669390400
transform -1 0 51296 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2347_
timestamp 1669390400
transform 1 0 53648 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2348_
timestamp 1669390400
transform -1 0 54544 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2349_
timestamp 1669390400
transform 1 0 52864 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2350_
timestamp 1669390400
transform 1 0 61264 0 1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _2351_
timestamp 1669390400
transform 1 0 61152 0 -1 17248
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2352_
timestamp 1669390400
transform 1 0 62496 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2353_
timestamp 1669390400
transform 1 0 55440 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2354_
timestamp 1669390400
transform -1 0 58016 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2355_
timestamp 1669390400
transform 1 0 56224 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2356_
timestamp 1669390400
transform -1 0 64064 0 -1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2357_
timestamp 1669390400
transform -1 0 63840 0 -1 14112
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2358_
timestamp 1669390400
transform -1 0 60592 0 -1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2359_
timestamp 1669390400
transform 1 0 48160 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2360_
timestamp 1669390400
transform -1 0 49952 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2361_
timestamp 1669390400
transform 1 0 48496 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2362_
timestamp 1669390400
transform -1 0 68544 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2363_
timestamp 1669390400
transform -1 0 56896 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2364_
timestamp 1669390400
transform 1 0 57792 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2365_
timestamp 1669390400
transform -1 0 58016 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2366_
timestamp 1669390400
transform 1 0 48384 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2367_
timestamp 1669390400
transform 1 0 49616 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2368_
timestamp 1669390400
transform -1 0 51296 0 1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2369_
timestamp 1669390400
transform 1 0 66528 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2370_
timestamp 1669390400
transform -1 0 67760 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2371_
timestamp 1669390400
transform 1 0 66640 0 1 9408
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2372_
timestamp 1669390400
transform -1 0 67872 0 -1 10976
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2373_
timestamp 1669390400
transform -1 0 64512 0 1 10976
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2374_
timestamp 1669390400
transform -1 0 62832 0 1 10976
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2375_
timestamp 1669390400
transform -1 0 56896 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2376_
timestamp 1669390400
transform 1 0 55776 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2377_
timestamp 1669390400
transform -1 0 56896 0 1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2378_
timestamp 1669390400
transform 1 0 52304 0 -1 7840
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2379_
timestamp 1669390400
transform 1 0 55216 0 1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2380_
timestamp 1669390400
transform 1 0 57568 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2381_
timestamp 1669390400
transform 1 0 58464 0 1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2382_
timestamp 1669390400
transform 1 0 59696 0 -1 6272
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2383_
timestamp 1669390400
transform 1 0 61712 0 1 6272
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2384_
timestamp 1669390400
transform -1 0 62272 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2385_
timestamp 1669390400
transform -1 0 65520 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2386_
timestamp 1669390400
transform 1 0 59248 0 1 7840
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2387_
timestamp 1669390400
transform 1 0 61264 0 1 7840
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2388_
timestamp 1669390400
transform -1 0 64288 0 1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2389_
timestamp 1669390400
transform -1 0 61936 0 -1 9408
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2390_
timestamp 1669390400
transform 1 0 59024 0 -1 12544
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2391_
timestamp 1669390400
transform -1 0 60480 0 1 12544
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2392_
timestamp 1669390400
transform -1 0 57568 0 1 14112
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2393_
timestamp 1669390400
transform -1 0 56672 0 -1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2394_
timestamp 1669390400
transform -1 0 54432 0 -1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2395_
timestamp 1669390400
transform -1 0 50064 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2396_
timestamp 1669390400
transform -1 0 51296 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2397_
timestamp 1669390400
transform 1 0 49392 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2398_
timestamp 1669390400
transform 1 0 53312 0 1 18816
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2399_
timestamp 1669390400
transform -1 0 55104 0 -1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _2400_
timestamp 1669390400
transform -1 0 53984 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2401_
timestamp 1669390400
transform 1 0 52640 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2402_
timestamp 1669390400
transform 1 0 53312 0 1 28224
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2403_
timestamp 1669390400
transform 1 0 52192 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2404_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 53312 0 -1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2405_
timestamp 1669390400
transform 1 0 53312 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2406_
timestamp 1669390400
transform -1 0 55776 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2407_
timestamp 1669390400
transform -1 0 54992 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2408_
timestamp 1669390400
transform -1 0 54656 0 1 21952
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2409_
timestamp 1669390400
transform -1 0 51968 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2410_
timestamp 1669390400
transform 1 0 52864 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2411_
timestamp 1669390400
transform -1 0 53984 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2412_
timestamp 1669390400
transform 1 0 53984 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2413_
timestamp 1669390400
transform 1 0 54656 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2414_
timestamp 1669390400
transform -1 0 58352 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2415_
timestamp 1669390400
transform 1 0 57344 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2416_
timestamp 1669390400
transform -1 0 62944 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2417_
timestamp 1669390400
transform 1 0 61264 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2418_
timestamp 1669390400
transform 1 0 60592 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2419_
timestamp 1669390400
transform 1 0 61264 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2420_
timestamp 1669390400
transform 1 0 63504 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2421_
timestamp 1669390400
transform -1 0 63728 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2422_
timestamp 1669390400
transform -1 0 63728 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2423_
timestamp 1669390400
transform 1 0 64288 0 1 15680
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2424_
timestamp 1669390400
transform 1 0 65296 0 -1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2425_
timestamp 1669390400
transform 1 0 65744 0 1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2426_
timestamp 1669390400
transform -1 0 62944 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2427_
timestamp 1669390400
transform -1 0 63728 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2428_
timestamp 1669390400
transform -1 0 62608 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2429_
timestamp 1669390400
transform -1 0 63168 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2430_
timestamp 1669390400
transform -1 0 63504 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2431_
timestamp 1669390400
transform -1 0 60144 0 -1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2432_
timestamp 1669390400
transform 1 0 55440 0 -1 6272
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2433_
timestamp 1669390400
transform 1 0 58352 0 -1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2434_
timestamp 1669390400
transform -1 0 63952 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2435_
timestamp 1669390400
transform 1 0 58800 0 -1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2436_
timestamp 1669390400
transform 1 0 65296 0 -1 4704
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2437_
timestamp 1669390400
transform 1 0 75152 0 1 4704
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2438_
timestamp 1669390400
transform 1 0 67200 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2439_
timestamp 1669390400
transform 1 0 64288 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2440_
timestamp 1669390400
transform 1 0 65296 0 1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2441_
timestamp 1669390400
transform 1 0 65296 0 1 6272
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2442_
timestamp 1669390400
transform 1 0 71344 0 -1 7840
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2443_
timestamp 1669390400
transform -1 0 77728 0 -1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2444_
timestamp 1669390400
transform 1 0 75824 0 -1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2445_
timestamp 1669390400
transform 1 0 70112 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2446_
timestamp 1669390400
transform -1 0 69888 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2447_
timestamp 1669390400
transform 1 0 68096 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2448_
timestamp 1669390400
transform 1 0 69104 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2449_
timestamp 1669390400
transform 1 0 62160 0 -1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2450_
timestamp 1669390400
transform 1 0 73248 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2451_
timestamp 1669390400
transform 1 0 70896 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2452_
timestamp 1669390400
transform 1 0 71344 0 -1 10976
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2453_
timestamp 1669390400
transform 1 0 74480 0 -1 10976
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2454_
timestamp 1669390400
transform -1 0 77504 0 -1 10976
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2455_
timestamp 1669390400
transform 1 0 75376 0 1 10976
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2456_
timestamp 1669390400
transform -1 0 77952 0 -1 12544
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2457_
timestamp 1669390400
transform -1 0 67536 0 1 12544
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2458_
timestamp 1669390400
transform -1 0 67424 0 1 14112
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2459_
timestamp 1669390400
transform -1 0 60816 0 1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2460_
timestamp 1669390400
transform -1 0 60368 0 1 15680
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2461_
timestamp 1669390400
transform -1 0 58800 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2462_
timestamp 1669390400
transform -1 0 58576 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2463_
timestamp 1669390400
transform 1 0 57568 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2464_
timestamp 1669390400
transform -1 0 57120 0 1 18816
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2465_
timestamp 1669390400
transform -1 0 54656 0 1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2466_
timestamp 1669390400
transform -1 0 52864 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _2467_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 63840 0 -1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2468_
timestamp 1669390400
transform -1 0 67760 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2469_
timestamp 1669390400
transform 1 0 67760 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2470_
timestamp 1669390400
transform 1 0 67648 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2471_
timestamp 1669390400
transform 1 0 76272 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2472_
timestamp 1669390400
transform -1 0 78288 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2473_
timestamp 1669390400
transform -1 0 75152 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2474_
timestamp 1669390400
transform 1 0 75712 0 -1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2475_
timestamp 1669390400
transform 1 0 77168 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2476_
timestamp 1669390400
transform 1 0 77168 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2477_
timestamp 1669390400
transform 1 0 74032 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2478_
timestamp 1669390400
transform 1 0 77168 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2479_
timestamp 1669390400
transform 1 0 59360 0 1 3136
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2480_
timestamp 1669390400
transform 1 0 57568 0 -1 4704
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2481_
timestamp 1669390400
transform -1 0 62160 0 -1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2482_
timestamp 1669390400
transform 1 0 66080 0 1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2483_
timestamp 1669390400
transform 1 0 60256 0 1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2484_
timestamp 1669390400
transform 1 0 68880 0 -1 4704
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2485_
timestamp 1669390400
transform 1 0 71344 0 1 4704
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2486_
timestamp 1669390400
transform 1 0 66416 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2487_
timestamp 1669390400
transform -1 0 69104 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2488_
timestamp 1669390400
transform 1 0 66528 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2489_
timestamp 1669390400
transform 1 0 69216 0 1 6272
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2490_
timestamp 1669390400
transform 1 0 71456 0 -1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2491_
timestamp 1669390400
transform 1 0 74816 0 -1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2492_
timestamp 1669390400
transform 1 0 71904 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2493_
timestamp 1669390400
transform 1 0 73248 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2494_
timestamp 1669390400
transform -1 0 73472 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2495_
timestamp 1669390400
transform 1 0 69216 0 -1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2496_
timestamp 1669390400
transform 1 0 70000 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2497_
timestamp 1669390400
transform -1 0 70336 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2498_
timestamp 1669390400
transform 1 0 70000 0 -1 12544
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2499_
timestamp 1669390400
transform 1 0 70000 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2500_
timestamp 1669390400
transform -1 0 72016 0 1 10976
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2501_
timestamp 1669390400
transform 1 0 70896 0 1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2502_
timestamp 1669390400
transform 1 0 72464 0 1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2503_
timestamp 1669390400
transform -1 0 76608 0 1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2504_
timestamp 1669390400
transform 1 0 75264 0 1 12544
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2505_
timestamp 1669390400
transform -1 0 77392 0 -1 14112
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2506_
timestamp 1669390400
transform 1 0 69216 0 1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2507_
timestamp 1669390400
transform -1 0 70672 0 1 17248
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2508_
timestamp 1669390400
transform -1 0 61488 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2509_
timestamp 1669390400
transform 1 0 60032 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2510_
timestamp 1669390400
transform -1 0 62608 0 -1 18816
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2511_
timestamp 1669390400
transform 1 0 59024 0 1 18816
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2512_
timestamp 1669390400
transform 1 0 55664 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2513_
timestamp 1669390400
transform -1 0 56560 0 1 20384
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2514_
timestamp 1669390400
transform -1 0 59136 0 1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2515_
timestamp 1669390400
transform -1 0 58352 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2516_
timestamp 1669390400
transform 1 0 58800 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2517_
timestamp 1669390400
transform 1 0 59584 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2518_
timestamp 1669390400
transform 1 0 61600 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2519_
timestamp 1669390400
transform 1 0 77168 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2520_
timestamp 1669390400
transform -1 0 77616 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2521_
timestamp 1669390400
transform 1 0 75152 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2522_
timestamp 1669390400
transform 1 0 77280 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2523_
timestamp 1669390400
transform -1 0 77728 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2524_
timestamp 1669390400
transform 1 0 70224 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2525_
timestamp 1669390400
transform 1 0 71456 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2526_
timestamp 1669390400
transform 1 0 73248 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2527_
timestamp 1669390400
transform 1 0 75040 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2528_
timestamp 1669390400
transform 1 0 74480 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2529_
timestamp 1669390400
transform 1 0 76608 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2530_
timestamp 1669390400
transform 1 0 71792 0 -1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2531_
timestamp 1669390400
transform -1 0 72912 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2532_
timestamp 1669390400
transform 1 0 62944 0 1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2533_
timestamp 1669390400
transform 1 0 66976 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2534_
timestamp 1669390400
transform 1 0 67536 0 1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2535_
timestamp 1669390400
transform 1 0 65296 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2536_
timestamp 1669390400
transform 1 0 58128 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2537_
timestamp 1669390400
transform 1 0 65072 0 1 18816
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2538_
timestamp 1669390400
transform 1 0 70000 0 1 18816
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2539_
timestamp 1669390400
transform 1 0 65296 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2540_
timestamp 1669390400
transform 1 0 65072 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2541_
timestamp 1669390400
transform 1 0 65408 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2542_
timestamp 1669390400
transform 1 0 65856 0 1 20384
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2543_
timestamp 1669390400
transform 1 0 70784 0 -1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2544_
timestamp 1669390400
transform 1 0 72016 0 1 15680
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2545_
timestamp 1669390400
transform 1 0 70784 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2546_
timestamp 1669390400
transform 1 0 71008 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2547_
timestamp 1669390400
transform -1 0 68320 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2548_
timestamp 1669390400
transform -1 0 68544 0 1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2549_
timestamp 1669390400
transform 1 0 66976 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2550_
timestamp 1669390400
transform 1 0 69216 0 1 14112
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2551_
timestamp 1669390400
transform 1 0 71232 0 1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2552_
timestamp 1669390400
transform 1 0 72800 0 1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2553_
timestamp 1669390400
transform 1 0 73696 0 1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2554_
timestamp 1669390400
transform -1 0 77952 0 -1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2555_
timestamp 1669390400
transform -1 0 76384 0 1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2556_
timestamp 1669390400
transform -1 0 77168 0 -1 18816
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2557_
timestamp 1669390400
transform -1 0 70560 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2558_
timestamp 1669390400
transform 1 0 70896 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2559_
timestamp 1669390400
transform -1 0 71232 0 -1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2560_
timestamp 1669390400
transform -1 0 62832 0 -1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2561_
timestamp 1669390400
transform 1 0 59360 0 1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2562_
timestamp 1669390400
transform -1 0 61040 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2563_
timestamp 1669390400
transform 1 0 69328 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2564_
timestamp 1669390400
transform 1 0 71456 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2565_
timestamp 1669390400
transform 1 0 75824 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2566_
timestamp 1669390400
transform -1 0 74816 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2567_
timestamp 1669390400
transform 1 0 71232 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2568_
timestamp 1669390400
transform 1 0 72352 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2569_
timestamp 1669390400
transform -1 0 73808 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2570_
timestamp 1669390400
transform 1 0 71904 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2571_
timestamp 1669390400
transform 1 0 73248 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2572_
timestamp 1669390400
transform -1 0 74368 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2573_
timestamp 1669390400
transform 1 0 69216 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2574_
timestamp 1669390400
transform -1 0 72464 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2575_
timestamp 1669390400
transform 1 0 58912 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2576_
timestamp 1669390400
transform 1 0 63952 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2577_
timestamp 1669390400
transform -1 0 66416 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2578_
timestamp 1669390400
transform 1 0 59584 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2579_
timestamp 1669390400
transform 1 0 58800 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2580_
timestamp 1669390400
transform 1 0 61040 0 -1 23520
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2581_
timestamp 1669390400
transform 1 0 70896 0 -1 23520
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2582_
timestamp 1669390400
transform 1 0 65296 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2583_
timestamp 1669390400
transform 1 0 64624 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2584_
timestamp 1669390400
transform 1 0 65184 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2585_
timestamp 1669390400
transform 1 0 66864 0 -1 23520
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2586_
timestamp 1669390400
transform 1 0 71792 0 1 21952
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2587_
timestamp 1669390400
transform -1 0 76720 0 1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2588_
timestamp 1669390400
transform 1 0 66192 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2589_
timestamp 1669390400
transform 1 0 66528 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2590_
timestamp 1669390400
transform 1 0 69216 0 1 20384
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2591_
timestamp 1669390400
transform 1 0 70560 0 -1 21952
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2592_
timestamp 1669390400
transform 1 0 73696 0 1 21952
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2593_
timestamp 1669390400
transform -1 0 75936 0 1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2594_
timestamp 1669390400
transform 1 0 74928 0 -1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2595_
timestamp 1669390400
transform -1 0 74704 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2596_
timestamp 1669390400
transform 1 0 76608 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2597_
timestamp 1669390400
transform -1 0 77840 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2598_
timestamp 1669390400
transform -1 0 74256 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2599_
timestamp 1669390400
transform 1 0 77168 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2600_
timestamp 1669390400
transform 1 0 77392 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2601_
timestamp 1669390400
transform -1 0 75040 0 1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2602_
timestamp 1669390400
transform -1 0 67312 0 1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2603_
timestamp 1669390400
transform -1 0 61824 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2604_
timestamp 1669390400
transform 1 0 55328 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2605_
timestamp 1669390400
transform -1 0 55216 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _2606_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 50176 0 -1 31360
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2607_
timestamp 1669390400
transform 1 0 61376 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _2608_
timestamp 1669390400
transform -1 0 63616 0 1 20384
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2609_
timestamp 1669390400
transform -1 0 62160 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2610_
timestamp 1669390400
transform -1 0 62608 0 1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2611_
timestamp 1669390400
transform -1 0 61264 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2612_
timestamp 1669390400
transform -1 0 68768 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2613_
timestamp 1669390400
transform -1 0 68096 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2614_
timestamp 1669390400
transform 1 0 62384 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _2615_
timestamp 1669390400
transform -1 0 63616 0 -1 31360
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2616_
timestamp 1669390400
transform 1 0 70112 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2617_
timestamp 1669390400
transform -1 0 71344 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2618_
timestamp 1669390400
transform 1 0 74592 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2619_
timestamp 1669390400
transform 1 0 76608 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2620_
timestamp 1669390400
transform 1 0 77168 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2621_
timestamp 1669390400
transform 1 0 64288 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2622_
timestamp 1669390400
transform 1 0 65744 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2623_
timestamp 1669390400
transform 1 0 66528 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2624_
timestamp 1669390400
transform 1 0 71008 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2625_
timestamp 1669390400
transform 1 0 73248 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2626_
timestamp 1669390400
transform 1 0 57344 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2627_
timestamp 1669390400
transform 1 0 58576 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2628_
timestamp 1669390400
transform -1 0 60816 0 -1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2629_
timestamp 1669390400
transform 1 0 57344 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2630_
timestamp 1669390400
transform 1 0 56896 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2631_
timestamp 1669390400
transform -1 0 58800 0 -1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2632_
timestamp 1669390400
transform 1 0 57232 0 1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2633_
timestamp 1669390400
transform 1 0 61152 0 -1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2634_
timestamp 1669390400
transform 1 0 66192 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2635_
timestamp 1669390400
transform 1 0 65296 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2636_
timestamp 1669390400
transform 1 0 65632 0 1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2637_
timestamp 1669390400
transform 1 0 67312 0 1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2638_
timestamp 1669390400
transform 1 0 70224 0 -1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2639_
timestamp 1669390400
transform 1 0 71456 0 1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2640_
timestamp 1669390400
transform 1 0 75264 0 -1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2641_
timestamp 1669390400
transform 1 0 75712 0 -1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2642_
timestamp 1669390400
transform 1 0 75376 0 1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2643_
timestamp 1669390400
transform 1 0 77168 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2644_
timestamp 1669390400
transform -1 0 74368 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2645_
timestamp 1669390400
transform 1 0 76608 0 -1 26656
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2646_
timestamp 1669390400
transform 1 0 76272 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2647_
timestamp 1669390400
transform -1 0 76720 0 1 28224
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2648_
timestamp 1669390400
transform -1 0 66976 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2649_
timestamp 1669390400
transform -1 0 67648 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2650_
timestamp 1669390400
transform -1 0 66528 0 -1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2651_
timestamp 1669390400
transform -1 0 66192 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2652_
timestamp 1669390400
transform -1 0 76048 0 -1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2653_
timestamp 1669390400
transform -1 0 71232 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2654_
timestamp 1669390400
transform -1 0 75488 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2655_
timestamp 1669390400
transform -1 0 77840 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2656_
timestamp 1669390400
transform 1 0 66416 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2657_
timestamp 1669390400
transform 1 0 66640 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2658_
timestamp 1669390400
transform 1 0 67536 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2659_
timestamp 1669390400
transform 1 0 61600 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2660_
timestamp 1669390400
transform -1 0 70112 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2661_
timestamp 1669390400
transform 1 0 62048 0 1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2662_
timestamp 1669390400
transform -1 0 65408 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2663_
timestamp 1669390400
transform 1 0 65632 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2664_
timestamp 1669390400
transform -1 0 65744 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2665_
timestamp 1669390400
transform -1 0 63504 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2666_
timestamp 1669390400
transform -1 0 59584 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2667_
timestamp 1669390400
transform 1 0 57680 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2668_
timestamp 1669390400
transform 1 0 58016 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2669_
timestamp 1669390400
transform 1 0 56336 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2670_
timestamp 1669390400
transform 1 0 56000 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2671_
timestamp 1669390400
transform -1 0 58352 0 -1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2672_
timestamp 1669390400
transform 1 0 56896 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2673_
timestamp 1669390400
transform 1 0 58016 0 1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2674_
timestamp 1669390400
transform 1 0 61040 0 -1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2675_
timestamp 1669390400
transform 1 0 62608 0 -1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2676_
timestamp 1669390400
transform 1 0 69216 0 1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2677_
timestamp 1669390400
transform 1 0 70224 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2678_
timestamp 1669390400
transform 1 0 70784 0 1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2679_
timestamp 1669390400
transform 1 0 71792 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2680_
timestamp 1669390400
transform -1 0 73808 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2681_
timestamp 1669390400
transform -1 0 72688 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2682_
timestamp 1669390400
transform 1 0 71344 0 -1 26656
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2683_
timestamp 1669390400
transform -1 0 74592 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2684_
timestamp 1669390400
transform 1 0 75488 0 1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2685_
timestamp 1669390400
transform 1 0 77392 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2686_
timestamp 1669390400
transform -1 0 77616 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2687_
timestamp 1669390400
transform 1 0 74592 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2688_
timestamp 1669390400
transform -1 0 78064 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2689_
timestamp 1669390400
transform -1 0 74704 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2690_
timestamp 1669390400
transform -1 0 76272 0 1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2691_
timestamp 1669390400
transform -1 0 71456 0 -1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2692_
timestamp 1669390400
transform -1 0 70112 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2693_
timestamp 1669390400
transform 1 0 61488 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2694_
timestamp 1669390400
transform 1 0 62608 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2695_
timestamp 1669390400
transform 1 0 63728 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2696_
timestamp 1669390400
transform 1 0 58016 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2697_
timestamp 1669390400
transform 1 0 58912 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2698_
timestamp 1669390400
transform -1 0 60032 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2699_
timestamp 1669390400
transform 1 0 54544 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2700_
timestamp 1669390400
transform 1 0 55440 0 -1 29792
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2701_
timestamp 1669390400
transform 1 0 57792 0 -1 29792
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2702_
timestamp 1669390400
transform 1 0 59472 0 1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2703_
timestamp 1669390400
transform 1 0 63952 0 1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2704_
timestamp 1669390400
transform 1 0 65520 0 1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2705_
timestamp 1669390400
transform 1 0 67088 0 1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2706_
timestamp 1669390400
transform 1 0 68208 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2707_
timestamp 1669390400
transform -1 0 70000 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2708_
timestamp 1669390400
transform 1 0 68880 0 -1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2709_
timestamp 1669390400
transform 1 0 72352 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2710_
timestamp 1669390400
transform -1 0 71792 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2711_
timestamp 1669390400
transform 1 0 70672 0 1 28224
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2712_
timestamp 1669390400
transform -1 0 78064 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2713_
timestamp 1669390400
transform -1 0 76496 0 -1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2714_
timestamp 1669390400
transform -1 0 74592 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2715_
timestamp 1669390400
transform -1 0 72240 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2716_
timestamp 1669390400
transform 1 0 71680 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2717_
timestamp 1669390400
transform -1 0 75152 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2718_
timestamp 1669390400
transform -1 0 73696 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2719_
timestamp 1669390400
transform -1 0 75936 0 -1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2720_
timestamp 1669390400
transform -1 0 75376 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2721_
timestamp 1669390400
transform 1 0 71232 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2722_
timestamp 1669390400
transform -1 0 64848 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2723_
timestamp 1669390400
transform -1 0 64176 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2724_
timestamp 1669390400
transform -1 0 66192 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2725_
timestamp 1669390400
transform 1 0 53760 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2726_
timestamp 1669390400
transform 1 0 53648 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2727_
timestamp 1669390400
transform -1 0 55888 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2728_
timestamp 1669390400
transform 1 0 54432 0 1 31360
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2729_
timestamp 1669390400
transform 1 0 57008 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2730_
timestamp 1669390400
transform 1 0 58016 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2731_
timestamp 1669390400
transform 1 0 58240 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2732_
timestamp 1669390400
transform -1 0 59920 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2733_
timestamp 1669390400
transform 1 0 60144 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2734_
timestamp 1669390400
transform -1 0 60592 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2735_
timestamp 1669390400
transform 1 0 61264 0 -1 28224
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2736_
timestamp 1669390400
transform 1 0 61264 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2737_
timestamp 1669390400
transform 1 0 61040 0 -1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2738_
timestamp 1669390400
transform -1 0 63952 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2739_
timestamp 1669390400
transform 1 0 62944 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2740_
timestamp 1669390400
transform 1 0 63280 0 1 31360
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2741_
timestamp 1669390400
transform 1 0 63728 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2742_
timestamp 1669390400
transform -1 0 69776 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2743_
timestamp 1669390400
transform -1 0 71008 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2744_
timestamp 1669390400
transform -1 0 67760 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2745_
timestamp 1669390400
transform 1 0 66080 0 1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2746_
timestamp 1669390400
transform -1 0 71680 0 -1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2747_
timestamp 1669390400
transform -1 0 72464 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2748_
timestamp 1669390400
transform -1 0 68768 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2749_
timestamp 1669390400
transform 1 0 76160 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2750_
timestamp 1669390400
transform 1 0 77168 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2751_
timestamp 1669390400
transform 1 0 69216 0 1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2752_
timestamp 1669390400
transform -1 0 69888 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2753_
timestamp 1669390400
transform 1 0 69440 0 1 31360
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2754_
timestamp 1669390400
transform 1 0 70000 0 1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2755_
timestamp 1669390400
transform 1 0 70672 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2756_
timestamp 1669390400
transform 1 0 66304 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2757_
timestamp 1669390400
transform 1 0 60368 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2758_
timestamp 1669390400
transform -1 0 61824 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2759_
timestamp 1669390400
transform 1 0 59248 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2760_
timestamp 1669390400
transform 1 0 50960 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2761_
timestamp 1669390400
transform 1 0 54208 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2762_
timestamp 1669390400
transform -1 0 55104 0 -1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2763_
timestamp 1669390400
transform -1 0 51968 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2764_
timestamp 1669390400
transform 1 0 51072 0 -1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2765_
timestamp 1669390400
transform 1 0 53312 0 1 32928
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2766_
timestamp 1669390400
transform -1 0 60144 0 1 34496
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2767_
timestamp 1669390400
transform 1 0 60368 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2768_
timestamp 1669390400
transform -1 0 65856 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2769_
timestamp 1669390400
transform -1 0 63280 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2770_
timestamp 1669390400
transform 1 0 62048 0 1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2771_
timestamp 1669390400
transform 1 0 63840 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2772_
timestamp 1669390400
transform 1 0 71568 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2773_
timestamp 1669390400
transform -1 0 70448 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2774_
timestamp 1669390400
transform 1 0 72016 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2775_
timestamp 1669390400
transform 1 0 69216 0 1 34496
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2776_
timestamp 1669390400
transform -1 0 71008 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2777_
timestamp 1669390400
transform -1 0 63392 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2778_
timestamp 1669390400
transform 1 0 54768 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2779_
timestamp 1669390400
transform 1 0 55328 0 -1 32928
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2780_
timestamp 1669390400
transform 1 0 53648 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2781_
timestamp 1669390400
transform -1 0 58016 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2782_
timestamp 1669390400
transform -1 0 56896 0 1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2783_
timestamp 1669390400
transform 1 0 54768 0 1 34496
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2784_
timestamp 1669390400
transform 1 0 55664 0 -1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2785_
timestamp 1669390400
transform -1 0 57344 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2786_
timestamp 1669390400
transform 1 0 57344 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2787_
timestamp 1669390400
transform 1 0 61152 0 -1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2788_
timestamp 1669390400
transform -1 0 69888 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2789_
timestamp 1669390400
transform 1 0 65968 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2790_
timestamp 1669390400
transform 1 0 65520 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2791_
timestamp 1669390400
transform -1 0 64848 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2792_
timestamp 1669390400
transform 1 0 65296 0 -1 36064
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2793_
timestamp 1669390400
transform 1 0 66976 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2794_
timestamp 1669390400
transform -1 0 60928 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2795_
timestamp 1669390400
transform -1 0 65744 0 1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2796_
timestamp 1669390400
transform -1 0 58240 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2797_
timestamp 1669390400
transform -1 0 59024 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _2798_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 57344 0 -1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _2799_
timestamp 1669390400
transform 1 0 58800 0 -1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2800_
timestamp 1669390400
transform 1 0 62720 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2801_
timestamp 1669390400
transform -1 0 20720 0 -1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2802_
timestamp 1669390400
transform -1 0 19152 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2803_
timestamp 1669390400
transform 1 0 22736 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2804_
timestamp 1669390400
transform 1 0 22400 0 1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2805_
timestamp 1669390400
transform 1 0 23296 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2806_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 1904 0 1 3136
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2807_
timestamp 1669390400
transform -1 0 78176 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2808_
timestamp 1669390400
transform -1 0 77280 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2809_
timestamp 1669390400
transform -1 0 78064 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2810_
timestamp 1669390400
transform -1 0 77392 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2811_
timestamp 1669390400
transform -1 0 77840 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2812_
timestamp 1669390400
transform 1 0 73920 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2813_
timestamp 1669390400
transform -1 0 77280 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2814_
timestamp 1669390400
transform -1 0 77728 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2815_
timestamp 1669390400
transform 1 0 73136 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2816_
timestamp 1669390400
transform -1 0 78176 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2817_
timestamp 1669390400
transform 1 0 77168 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2818_
timestamp 1669390400
transform -1 0 75712 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2819_
timestamp 1669390400
transform -1 0 76720 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2820_
timestamp 1669390400
transform 1 0 73920 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2821_
timestamp 1669390400
transform 1 0 72352 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2822_
timestamp 1669390400
transform 1 0 72128 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2823_
timestamp 1669390400
transform -1 0 4144 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2824_
timestamp 1669390400
transform -1 0 4144 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2825_
timestamp 1669390400
transform 1 0 2576 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2826_
timestamp 1669390400
transform 1 0 2240 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2827_
timestamp 1669390400
transform -1 0 3360 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2828_
timestamp 1669390400
transform -1 0 3360 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2829_
timestamp 1669390400
transform -1 0 2576 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2830_
timestamp 1669390400
transform -1 0 4144 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2831_
timestamp 1669390400
transform -1 0 3360 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2832_
timestamp 1669390400
transform -1 0 3248 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2833_
timestamp 1669390400
transform -1 0 3360 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2834_
timestamp 1669390400
transform -1 0 3360 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2835_
timestamp 1669390400
transform -1 0 3360 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2836_
timestamp 1669390400
transform -1 0 4144 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2837_
timestamp 1669390400
transform -1 0 4144 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2838_
timestamp 1669390400
transform -1 0 5040 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input1
timestamp 1669390400
transform 1 0 12096 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input2
timestamp 1669390400
transform 1 0 33040 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input3
timestamp 1669390400
transform 1 0 34720 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input4 Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 36960 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input5
timestamp 1669390400
transform 1 0 38976 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input6
timestamp 1669390400
transform 1 0 41104 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dlyd_1  input7 Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 43232 0 -1 4704
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input8
timestamp 1669390400
transform 1 0 13440 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input9
timestamp 1669390400
transform -1 0 16800 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input10
timestamp 1669390400
transform 1 0 17696 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input11
timestamp 1669390400
transform -1 0 19152 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input12
timestamp 1669390400
transform 1 0 21952 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input13
timestamp 1669390400
transform -1 0 24752 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input14
timestamp 1669390400
transform 1 0 26208 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input15
timestamp 1669390400
transform 1 0 29120 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input16
timestamp 1669390400
transform 1 0 30464 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input17
timestamp 1669390400
transform -1 0 48160 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input18
timestamp 1669390400
transform -1 0 66752 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input19 Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 70560 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input20
timestamp 1669390400
transform -1 0 71568 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input21
timestamp 1669390400
transform -1 0 73696 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input22
timestamp 1669390400
transform -1 0 74592 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input23
timestamp 1669390400
transform -1 0 77056 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  input24 Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 51520 0 1 3136
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input25
timestamp 1669390400
transform 1 0 49616 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input26
timestamp 1669390400
transform 1 0 52640 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input27
timestamp 1669390400
transform -1 0 55328 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input28
timestamp 1669390400
transform 1 0 56000 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input29
timestamp 1669390400
transform -1 0 59136 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  input30
timestamp 1669390400
transform -1 0 63280 0 1 3136
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input31
timestamp 1669390400
transform -1 0 64176 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input32
timestamp 1669390400
transform 1 0 64512 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input33
timestamp 1669390400
transform -1 0 8848 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output34 Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 3360 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output35
timestamp 1669390400
transform -1 0 28000 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output36
timestamp 1669390400
transform -1 0 30688 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output37
timestamp 1669390400
transform -1 0 32592 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output38
timestamp 1669390400
transform -1 0 35392 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output39
timestamp 1669390400
transform -1 0 37856 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output40
timestamp 1669390400
transform -1 0 40320 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output41
timestamp 1669390400
transform -1 0 42784 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output42
timestamp 1669390400
transform -1 0 45248 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output43
timestamp 1669390400
transform -1 0 47712 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output44
timestamp 1669390400
transform -1 0 50288 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output45
timestamp 1669390400
transform -1 0 5152 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output46
timestamp 1669390400
transform -1 0 52192 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output47
timestamp 1669390400
transform 1 0 53536 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output48
timestamp 1669390400
transform -1 0 58128 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output49
timestamp 1669390400
transform -1 0 60032 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output50
timestamp 1669390400
transform 1 0 60928 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output51
timestamp 1669390400
transform -1 0 65968 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output52
timestamp 1669390400
transform -1 0 67760 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output53
timestamp 1669390400
transform -1 0 69888 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output54
timestamp 1669390400
transform -1 0 71792 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output55
timestamp 1669390400
transform 1 0 73248 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output56
timestamp 1669390400
transform -1 0 8288 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output57
timestamp 1669390400
transform 1 0 76160 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output58
timestamp 1669390400
transform 1 0 74816 0 1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output59
timestamp 1669390400
transform -1 0 11088 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output60
timestamp 1669390400
transform -1 0 12992 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output61
timestamp 1669390400
transform -1 0 15680 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output62
timestamp 1669390400
transform -1 0 19152 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output63
timestamp 1669390400
transform -1 0 20608 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output64
timestamp 1669390400
transform -1 0 22960 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output65
timestamp 1669390400
transform -1 0 24752 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output66
timestamp 1669390400
transform 1 0 9520 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output67
timestamp 1669390400
transform -1 0 75712 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output68
timestamp 1669390400
transform -1 0 76384 0 -1 26656
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output69
timestamp 1669390400
transform 1 0 74816 0 -1 29792
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output70
timestamp 1669390400
transform -1 0 76384 0 1 31360
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output71
timestamp 1669390400
transform 1 0 74816 0 -1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output72
timestamp 1669390400
transform 1 0 74816 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output73
timestamp 1669390400
transform 1 0 76608 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output74
timestamp 1669390400
transform -1 0 76384 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output75
timestamp 1669390400
transform -1 0 76384 0 1 6272
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output76
timestamp 1669390400
transform -1 0 76384 0 -1 9408
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output77
timestamp 1669390400
transform -1 0 76384 0 -1 12544
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output78
timestamp 1669390400
transform 1 0 74816 0 1 14112
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output79
timestamp 1669390400
transform 1 0 74816 0 -1 17248
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output80
timestamp 1669390400
transform -1 0 76384 0 1 18816
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output81
timestamp 1669390400
transform 1 0 74816 0 -1 21952
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output82
timestamp 1669390400
transform -1 0 76384 0 1 23520
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output83
timestamp 1669390400
transform -1 0 3248 0 1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output84
timestamp 1669390400
transform -1 0 3248 0 -1 26656
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output85
timestamp 1669390400
transform -1 0 3248 0 -1 29792
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output86
timestamp 1669390400
transform -1 0 3248 0 1 31360
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output87
timestamp 1669390400
transform -1 0 3248 0 -1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output88
timestamp 1669390400
transform -1 0 3248 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output89
timestamp 1669390400
transform -1 0 3248 0 1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output90
timestamp 1669390400
transform -1 0 3248 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output91
timestamp 1669390400
transform -1 0 3248 0 1 6272
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output92
timestamp 1669390400
transform -1 0 3248 0 -1 9408
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output93
timestamp 1669390400
transform -1 0 3248 0 -1 12544
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output94
timestamp 1669390400
transform -1 0 3248 0 1 14112
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output95
timestamp 1669390400
transform 1 0 1680 0 -1 17248
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output96
timestamp 1669390400
transform -1 0 3248 0 1 18816
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output97
timestamp 1669390400
transform -1 0 3248 0 1 20384
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output98
timestamp 1669390400
transform -1 0 3248 0 1 23520
box -86 -86 1654 870
<< labels >>
flabel metal2 s 1680 39200 1792 40000 0 FreeSans 448 90 0 0 Y[0]
port 0 nsew signal tristate
flabel metal2 s 26320 39200 26432 40000 0 FreeSans 448 90 0 0 Y[10]
port 1 nsew signal tristate
flabel metal2 s 28784 39200 28896 40000 0 FreeSans 448 90 0 0 Y[11]
port 2 nsew signal tristate
flabel metal2 s 31248 39200 31360 40000 0 FreeSans 448 90 0 0 Y[12]
port 3 nsew signal tristate
flabel metal2 s 33712 39200 33824 40000 0 FreeSans 448 90 0 0 Y[13]
port 4 nsew signal tristate
flabel metal2 s 36176 39200 36288 40000 0 FreeSans 448 90 0 0 Y[14]
port 5 nsew signal tristate
flabel metal2 s 38640 39200 38752 40000 0 FreeSans 448 90 0 0 Y[15]
port 6 nsew signal tristate
flabel metal2 s 41104 39200 41216 40000 0 FreeSans 448 90 0 0 Y[16]
port 7 nsew signal tristate
flabel metal2 s 43568 39200 43680 40000 0 FreeSans 448 90 0 0 Y[17]
port 8 nsew signal tristate
flabel metal2 s 46032 39200 46144 40000 0 FreeSans 448 90 0 0 Y[18]
port 9 nsew signal tristate
flabel metal2 s 48496 39200 48608 40000 0 FreeSans 448 90 0 0 Y[19]
port 10 nsew signal tristate
flabel metal2 s 4144 39200 4256 40000 0 FreeSans 448 90 0 0 Y[1]
port 11 nsew signal tristate
flabel metal2 s 50960 39200 51072 40000 0 FreeSans 448 90 0 0 Y[20]
port 12 nsew signal tristate
flabel metal2 s 53424 39200 53536 40000 0 FreeSans 448 90 0 0 Y[21]
port 13 nsew signal tristate
flabel metal2 s 55888 39200 56000 40000 0 FreeSans 448 90 0 0 Y[22]
port 14 nsew signal tristate
flabel metal2 s 58352 39200 58464 40000 0 FreeSans 448 90 0 0 Y[23]
port 15 nsew signal tristate
flabel metal2 s 60816 39200 60928 40000 0 FreeSans 448 90 0 0 Y[24]
port 16 nsew signal tristate
flabel metal2 s 63280 39200 63392 40000 0 FreeSans 448 90 0 0 Y[25]
port 17 nsew signal tristate
flabel metal2 s 65744 39200 65856 40000 0 FreeSans 448 90 0 0 Y[26]
port 18 nsew signal tristate
flabel metal2 s 68208 39200 68320 40000 0 FreeSans 448 90 0 0 Y[27]
port 19 nsew signal tristate
flabel metal2 s 70672 39200 70784 40000 0 FreeSans 448 90 0 0 Y[28]
port 20 nsew signal tristate
flabel metal2 s 73136 39200 73248 40000 0 FreeSans 448 90 0 0 Y[29]
port 21 nsew signal tristate
flabel metal2 s 6608 39200 6720 40000 0 FreeSans 448 90 0 0 Y[2]
port 22 nsew signal tristate
flabel metal2 s 75600 39200 75712 40000 0 FreeSans 448 90 0 0 Y[30]
port 23 nsew signal tristate
flabel metal2 s 78064 39200 78176 40000 0 FreeSans 448 90 0 0 Y[31]
port 24 nsew signal tristate
flabel metal2 s 9072 39200 9184 40000 0 FreeSans 448 90 0 0 Y[3]
port 25 nsew signal tristate
flabel metal2 s 11536 39200 11648 40000 0 FreeSans 448 90 0 0 Y[4]
port 26 nsew signal tristate
flabel metal2 s 14000 39200 14112 40000 0 FreeSans 448 90 0 0 Y[5]
port 27 nsew signal tristate
flabel metal2 s 16464 39200 16576 40000 0 FreeSans 448 90 0 0 Y[6]
port 28 nsew signal tristate
flabel metal2 s 18928 39200 19040 40000 0 FreeSans 448 90 0 0 Y[7]
port 29 nsew signal tristate
flabel metal2 s 21392 39200 21504 40000 0 FreeSans 448 90 0 0 Y[8]
port 30 nsew signal tristate
flabel metal2 s 23856 39200 23968 40000 0 FreeSans 448 90 0 0 Y[9]
port 31 nsew signal tristate
flabel metal2 s 2688 0 2800 800 0 FreeSans 448 90 0 0 clk
port 32 nsew signal input
flabel metal2 s 11200 0 11312 800 0 FreeSans 448 90 0 0 dba[0]
port 33 nsew signal input
flabel metal2 s 32480 0 32592 800 0 FreeSans 448 90 0 0 dba[10]
port 34 nsew signal input
flabel metal2 s 34608 0 34720 800 0 FreeSans 448 90 0 0 dba[11]
port 35 nsew signal input
flabel metal2 s 36736 0 36848 800 0 FreeSans 448 90 0 0 dba[12]
port 36 nsew signal input
flabel metal2 s 38864 0 38976 800 0 FreeSans 448 90 0 0 dba[13]
port 37 nsew signal input
flabel metal2 s 40992 0 41104 800 0 FreeSans 448 90 0 0 dba[14]
port 38 nsew signal input
flabel metal2 s 43120 0 43232 800 0 FreeSans 448 90 0 0 dba[15]
port 39 nsew signal input
flabel metal2 s 13328 0 13440 800 0 FreeSans 448 90 0 0 dba[1]
port 40 nsew signal input
flabel metal2 s 15456 0 15568 800 0 FreeSans 448 90 0 0 dba[2]
port 41 nsew signal input
flabel metal2 s 17584 0 17696 800 0 FreeSans 448 90 0 0 dba[3]
port 42 nsew signal input
flabel metal2 s 19712 0 19824 800 0 FreeSans 448 90 0 0 dba[4]
port 43 nsew signal input
flabel metal2 s 21840 0 21952 800 0 FreeSans 448 90 0 0 dba[5]
port 44 nsew signal input
flabel metal2 s 23968 0 24080 800 0 FreeSans 448 90 0 0 dba[6]
port 45 nsew signal input
flabel metal2 s 26096 0 26208 800 0 FreeSans 448 90 0 0 dba[7]
port 46 nsew signal input
flabel metal2 s 28224 0 28336 800 0 FreeSans 448 90 0 0 dba[8]
port 47 nsew signal input
flabel metal2 s 30352 0 30464 800 0 FreeSans 448 90 0 0 dba[9]
port 48 nsew signal input
flabel metal2 s 45248 0 45360 800 0 FreeSans 448 90 0 0 dbb[0]
port 49 nsew signal input
flabel metal2 s 66528 0 66640 800 0 FreeSans 448 90 0 0 dbb[10]
port 50 nsew signal input
flabel metal2 s 68656 0 68768 800 0 FreeSans 448 90 0 0 dbb[11]
port 51 nsew signal input
flabel metal2 s 70784 0 70896 800 0 FreeSans 448 90 0 0 dbb[12]
port 52 nsew signal input
flabel metal2 s 72912 0 73024 800 0 FreeSans 448 90 0 0 dbb[13]
port 53 nsew signal input
flabel metal2 s 75040 0 75152 800 0 FreeSans 448 90 0 0 dbb[14]
port 54 nsew signal input
flabel metal2 s 77168 0 77280 800 0 FreeSans 448 90 0 0 dbb[15]
port 55 nsew signal input
flabel metal2 s 47376 0 47488 800 0 FreeSans 448 90 0 0 dbb[1]
port 56 nsew signal input
flabel metal2 s 49504 0 49616 800 0 FreeSans 448 90 0 0 dbb[2]
port 57 nsew signal input
flabel metal2 s 51632 0 51744 800 0 FreeSans 448 90 0 0 dbb[3]
port 58 nsew signal input
flabel metal2 s 53760 0 53872 800 0 FreeSans 448 90 0 0 dbb[4]
port 59 nsew signal input
flabel metal2 s 55888 0 56000 800 0 FreeSans 448 90 0 0 dbb[5]
port 60 nsew signal input
flabel metal2 s 58016 0 58128 800 0 FreeSans 448 90 0 0 dbb[6]
port 61 nsew signal input
flabel metal2 s 60144 0 60256 800 0 FreeSans 448 90 0 0 dbb[7]
port 62 nsew signal input
flabel metal2 s 62272 0 62384 800 0 FreeSans 448 90 0 0 dbb[8]
port 63 nsew signal input
flabel metal2 s 64400 0 64512 800 0 FreeSans 448 90 0 0 dbb[9]
port 64 nsew signal input
flabel metal2 s 9072 0 9184 800 0 FreeSans 448 90 0 0 done
port 65 nsew signal tristate
flabel metal2 s 6944 0 7056 800 0 FreeSans 448 90 0 0 enable
port 66 nsew signal input
flabel metal2 s 4816 0 4928 800 0 FreeSans 448 90 0 0 rst
port 67 nsew signal input
flabel metal4 s 10844 3076 11164 36908 0 FreeSans 1280 90 0 0 vdd
port 68 nsew power bidirectional
flabel metal4 s 30164 3076 30484 36908 0 FreeSans 1280 90 0 0 vdd
port 68 nsew power bidirectional
flabel metal4 s 49484 3076 49804 36908 0 FreeSans 1280 90 0 0 vdd
port 68 nsew power bidirectional
flabel metal4 s 68804 3076 69124 36908 0 FreeSans 1280 90 0 0 vdd
port 68 nsew power bidirectional
flabel metal4 s 20504 3076 20824 36908 0 FreeSans 1280 90 0 0 vss
port 69 nsew ground bidirectional
flabel metal4 s 39824 3076 40144 36908 0 FreeSans 1280 90 0 0 vss
port 69 nsew ground bidirectional
flabel metal4 s 59144 3076 59464 36908 0 FreeSans 1280 90 0 0 vss
port 69 nsew ground bidirectional
flabel metal4 s 78464 3076 78784 36908 0 FreeSans 1280 90 0 0 vss
port 69 nsew ground bidirectional
flabel metal3 s 79200 1456 80000 1568 0 FreeSans 448 0 0 0 yA[0]
port 70 nsew signal tristate
flabel metal3 s 79200 26096 80000 26208 0 FreeSans 448 0 0 0 yA[10]
port 71 nsew signal tristate
flabel metal3 s 79200 28560 80000 28672 0 FreeSans 448 0 0 0 yA[11]
port 72 nsew signal tristate
flabel metal3 s 79200 31024 80000 31136 0 FreeSans 448 0 0 0 yA[12]
port 73 nsew signal tristate
flabel metal3 s 79200 33488 80000 33600 0 FreeSans 448 0 0 0 yA[13]
port 74 nsew signal tristate
flabel metal3 s 79200 35952 80000 36064 0 FreeSans 448 0 0 0 yA[14]
port 75 nsew signal tristate
flabel metal3 s 79200 38416 80000 38528 0 FreeSans 448 0 0 0 yA[15]
port 76 nsew signal tristate
flabel metal3 s 79200 3920 80000 4032 0 FreeSans 448 0 0 0 yA[1]
port 77 nsew signal tristate
flabel metal3 s 79200 6384 80000 6496 0 FreeSans 448 0 0 0 yA[2]
port 78 nsew signal tristate
flabel metal3 s 79200 8848 80000 8960 0 FreeSans 448 0 0 0 yA[3]
port 79 nsew signal tristate
flabel metal3 s 79200 11312 80000 11424 0 FreeSans 448 0 0 0 yA[4]
port 80 nsew signal tristate
flabel metal3 s 79200 13776 80000 13888 0 FreeSans 448 0 0 0 yA[5]
port 81 nsew signal tristate
flabel metal3 s 79200 16240 80000 16352 0 FreeSans 448 0 0 0 yA[6]
port 82 nsew signal tristate
flabel metal3 s 79200 18704 80000 18816 0 FreeSans 448 0 0 0 yA[7]
port 83 nsew signal tristate
flabel metal3 s 79200 21168 80000 21280 0 FreeSans 448 0 0 0 yA[8]
port 84 nsew signal tristate
flabel metal3 s 79200 23632 80000 23744 0 FreeSans 448 0 0 0 yA[9]
port 85 nsew signal tristate
flabel metal3 s 0 1456 800 1568 0 FreeSans 448 0 0 0 yB[0]
port 86 nsew signal tristate
flabel metal3 s 0 26096 800 26208 0 FreeSans 448 0 0 0 yB[10]
port 87 nsew signal tristate
flabel metal3 s 0 28560 800 28672 0 FreeSans 448 0 0 0 yB[11]
port 88 nsew signal tristate
flabel metal3 s 0 31024 800 31136 0 FreeSans 448 0 0 0 yB[12]
port 89 nsew signal tristate
flabel metal3 s 0 33488 800 33600 0 FreeSans 448 0 0 0 yB[13]
port 90 nsew signal tristate
flabel metal3 s 0 35952 800 36064 0 FreeSans 448 0 0 0 yB[14]
port 91 nsew signal tristate
flabel metal3 s 0 38416 800 38528 0 FreeSans 448 0 0 0 yB[15]
port 92 nsew signal tristate
flabel metal3 s 0 3920 800 4032 0 FreeSans 448 0 0 0 yB[1]
port 93 nsew signal tristate
flabel metal3 s 0 6384 800 6496 0 FreeSans 448 0 0 0 yB[2]
port 94 nsew signal tristate
flabel metal3 s 0 8848 800 8960 0 FreeSans 448 0 0 0 yB[3]
port 95 nsew signal tristate
flabel metal3 s 0 11312 800 11424 0 FreeSans 448 0 0 0 yB[4]
port 96 nsew signal tristate
flabel metal3 s 0 13776 800 13888 0 FreeSans 448 0 0 0 yB[5]
port 97 nsew signal tristate
flabel metal3 s 0 16240 800 16352 0 FreeSans 448 0 0 0 yB[6]
port 98 nsew signal tristate
flabel metal3 s 0 18704 800 18816 0 FreeSans 448 0 0 0 yB[7]
port 99 nsew signal tristate
flabel metal3 s 0 21168 800 21280 0 FreeSans 448 0 0 0 yB[8]
port 100 nsew signal tristate
flabel metal3 s 0 23632 800 23744 0 FreeSans 448 0 0 0 yB[9]
port 101 nsew signal tristate
rlabel metal1 39984 36848 39984 36848 0 vdd
rlabel via1 40064 36064 40064 36064 0 vss
rlabel metal2 2072 37240 2072 37240 0 Y[0]
rlabel metal2 26712 37240 26712 37240 0 Y[10]
rlabel metal2 29400 37240 29400 37240 0 Y[11]
rlabel metal2 31304 37898 31304 37898 0 Y[12]
rlabel metal2 34104 37352 34104 37352 0 Y[13]
rlabel metal2 36568 36624 36568 36624 0 Y[14]
rlabel metal2 39032 36624 39032 36624 0 Y[15]
rlabel metal2 41496 37240 41496 37240 0 Y[16]
rlabel metal2 43792 35784 43792 35784 0 Y[17]
rlabel metal2 46424 37240 46424 37240 0 Y[18]
rlabel metal3 48776 36568 48776 36568 0 Y[19]
rlabel metal2 4200 37898 4200 37898 0 Y[1]
rlabel metal2 51016 37898 51016 37898 0 Y[20]
rlabel metal3 53928 36568 53928 36568 0 Y[21]
rlabel metal2 56840 37912 56840 37912 0 Y[22]
rlabel metal3 58632 36568 58632 36568 0 Y[23]
rlabel metal2 61768 37912 61768 37912 0 Y[24]
rlabel metal3 64008 36568 64008 36568 0 Y[25]
rlabel metal2 66472 37912 66472 37912 0 Y[26]
rlabel metal2 68600 37352 68600 37352 0 Y[27]
rlabel metal2 70728 37898 70728 37898 0 Y[28]
rlabel metal3 73640 36568 73640 36568 0 Y[29]
rlabel metal2 6832 36568 6832 36568 0 Y[2]
rlabel metal2 77000 37912 77000 37912 0 Y[30]
rlabel metal3 77112 35000 77112 35000 0 Y[31]
rlabel metal2 9800 37912 9800 37912 0 Y[3]
rlabel metal2 11704 36568 11704 36568 0 Y[4]
rlabel metal2 14224 36568 14224 36568 0 Y[5]
rlabel metal3 17192 35784 17192 35784 0 Y[6]
rlabel metal2 19152 36568 19152 36568 0 Y[7]
rlabel metal2 21560 36568 21560 36568 0 Y[8]
rlabel metal2 23912 37898 23912 37898 0 Y[9]
rlabel metal2 55496 7392 55496 7392 0 _0000_
rlabel metal2 54712 7112 54712 7112 0 _0001_
rlabel metal2 57064 6272 57064 6272 0 _0002_
rlabel metal2 56728 8288 56728 8288 0 _0003_
rlabel metal2 54824 8456 54824 8456 0 _0004_
rlabel metal2 49840 10584 49840 10584 0 _0005_
rlabel metal2 48496 12152 48496 12152 0 _0006_
rlabel metal2 50120 12432 50120 12432 0 _0007_
rlabel metal2 48776 13664 48776 13664 0 _0008_
rlabel metal2 49448 13832 49448 13832 0 _0009_
rlabel metal2 20216 25872 20216 25872 0 _0010_
rlabel metal2 49392 14728 49392 14728 0 _0011_
rlabel metal2 50344 20496 50344 20496 0 _0012_
rlabel metal2 52584 27496 52584 27496 0 _0013_
rlabel metal2 52808 25256 52808 25256 0 _0014_
rlabel metal2 53816 27048 53816 27048 0 _0015_
rlabel metal3 51744 26264 51744 26264 0 _0016_
rlabel metal2 48440 14112 48440 14112 0 _0017_
rlabel metal3 50568 14392 50568 14392 0 _0018_
rlabel metal3 52472 18424 52472 18424 0 _0019_
rlabel metal2 19264 29176 19264 29176 0 _0020_
rlabel metal2 55048 12040 55048 12040 0 _0021_
rlabel metal2 55720 13440 55720 13440 0 _0022_
rlabel metal3 55552 16856 55552 16856 0 _0023_
rlabel metal2 48888 12544 48888 12544 0 _0024_
rlabel metal2 57176 13776 57176 13776 0 _0025_
rlabel metal2 59864 13608 59864 13608 0 _0026_
rlabel metal2 53872 10584 53872 10584 0 _0027_
rlabel metal2 53144 10920 53144 10920 0 _0028_
rlabel metal3 62328 16184 62328 16184 0 _0029_
rlabel metal3 63280 16184 63280 16184 0 _0030_
rlabel metal2 19208 30520 19208 30520 0 _0031_
rlabel metal2 63280 15288 63280 15288 0 _0032_
rlabel metal2 56616 16128 56616 16128 0 _0033_
rlabel metal2 57512 16128 57512 16128 0 _0034_
rlabel metal2 63000 15344 63000 15344 0 _0035_
rlabel metal2 62776 14056 62776 14056 0 _0036_
rlabel metal3 60872 14280 60872 14280 0 _0037_
rlabel metal2 59976 12880 59976 12880 0 _0038_
rlabel metal2 48552 10528 48552 10528 0 _0039_
rlabel metal2 49392 10808 49392 10808 0 _0040_
rlabel metal2 59528 11704 59528 11704 0 _0041_
rlabel metal3 21224 31752 21224 31752 0 _0042_
rlabel metal2 68376 10192 68376 10192 0 _0043_
rlabel metal3 57064 10584 57064 10584 0 _0044_
rlabel metal2 57960 10696 57960 10696 0 _0045_
rlabel metal2 62216 11088 62216 11088 0 _0046_
rlabel metal2 50456 7784 50456 7784 0 _0047_
rlabel metal3 50568 8232 50568 8232 0 _0048_
rlabel metal3 51688 9688 51688 9688 0 _0049_
rlabel metal3 67984 10584 67984 10584 0 _0050_
rlabel metal2 67256 9576 67256 9576 0 _0051_
rlabel metal2 67592 10416 67592 10416 0 _0052_
rlabel metal2 22624 31864 22624 31864 0 _0053_
rlabel metal3 65240 11480 65240 11480 0 _0054_
rlabel metal3 62832 11480 62832 11480 0 _0055_
rlabel metal2 61544 10136 61544 10136 0 _0056_
rlabel metal2 56616 8736 56616 8736 0 _0057_
rlabel metal2 60872 8960 60872 8960 0 _0058_
rlabel metal3 58352 5320 58352 5320 0 _0059_
rlabel metal2 52808 7000 52808 7000 0 _0060_
rlabel metal2 62104 6832 62104 6832 0 _0061_
rlabel metal3 59248 5768 59248 5768 0 _0062_
rlabel metal2 61544 4704 61544 4704 0 _0063_
rlabel metal2 62216 6384 62216 6384 0 _0064_
rlabel metal3 63336 7672 63336 7672 0 _0065_
rlabel metal2 62216 9016 62216 9016 0 _0066_
rlabel metal2 69776 7672 69776 7672 0 _0067_
rlabel metal3 61040 8344 61040 8344 0 _0068_
rlabel metal2 63336 7896 63336 7896 0 _0069_
rlabel metal2 62776 9576 62776 9576 0 _0070_
rlabel metal2 59752 10416 59752 10416 0 _0071_
rlabel metal3 60760 12936 60760 12936 0 _0072_
rlabel metal2 58184 14112 58184 14112 0 _0073_
rlabel metal2 20328 32200 20328 32200 0 _0074_
rlabel metal3 57064 16744 57064 16744 0 _0075_
rlabel metal3 54600 18312 54600 18312 0 _0076_
rlabel metal2 53704 19264 53704 19264 0 _0077_
rlabel metal2 49560 18816 49560 18816 0 _0078_
rlabel metal2 50232 18704 50232 18704 0 _0079_
rlabel metal2 49672 19040 49672 19040 0 _0080_
rlabel metal2 53592 21112 53592 21112 0 _0081_
rlabel metal2 53816 27608 53816 27608 0 _0082_
rlabel metal2 52752 29176 52752 29176 0 _0083_
rlabel metal3 53872 28504 53872 28504 0 _0084_
rlabel metal3 12096 27832 12096 27832 0 _0085_
rlabel metal2 54040 28504 54040 28504 0 _0086_
rlabel metal2 52696 22624 52696 22624 0 _0087_
rlabel metal2 53648 23912 53648 23912 0 _0088_
rlabel metal3 54880 27160 54880 27160 0 _0089_
rlabel metal2 55048 28504 55048 28504 0 _0090_
rlabel metal2 54768 28056 54768 28056 0 _0091_
rlabel metal3 52640 22232 52640 22232 0 _0092_
rlabel metal3 55160 19992 55160 19992 0 _0093_
rlabel metal2 54152 20048 54152 20048 0 _0094_
rlabel metal2 45976 6720 45976 6720 0 _0095_
rlabel metal2 54208 20216 54208 20216 0 _0096_
rlabel metal2 56280 18928 56280 18928 0 _0097_
rlabel metal2 58072 14924 58072 14924 0 _0098_
rlabel metal2 58632 17416 58632 17416 0 _0099_
rlabel metal2 62272 14504 62272 14504 0 _0100_
rlabel metal2 60424 15680 60424 15680 0 _0101_
rlabel metal2 61600 12376 61600 12376 0 _0102_
rlabel metal3 61320 13832 61320 13832 0 _0103_
rlabel metal2 67368 16464 67368 16464 0 _0104_
rlabel metal2 63112 11480 63112 11480 0 _0105_
rlabel metal2 16240 26936 16240 26936 0 _0106_
rlabel metal3 64344 15176 64344 15176 0 _0107_
rlabel metal3 65296 16296 65296 16296 0 _0108_
rlabel metal2 66472 16464 66472 16464 0 _0109_
rlabel metal2 66920 15232 66920 15232 0 _0110_
rlabel metal2 62440 10304 62440 10304 0 _0111_
rlabel metal3 62720 10024 62720 10024 0 _0112_
rlabel metal2 66808 12712 66808 12712 0 _0113_
rlabel metal2 62664 6776 62664 6776 0 _0114_
rlabel metal3 74928 8120 74928 8120 0 _0115_
rlabel metal2 59640 4816 59640 4816 0 _0116_
rlabel metal2 14840 27440 14840 27440 0 _0117_
rlabel metal3 57400 5880 57400 5880 0 _0118_
rlabel metal2 74312 6440 74312 6440 0 _0119_
rlabel metal3 64792 5656 64792 5656 0 _0120_
rlabel metal2 70280 4816 70280 4816 0 _0121_
rlabel via2 74200 4984 74200 4984 0 _0122_
rlabel metal2 77000 5600 77000 5600 0 _0123_
rlabel metal3 70560 7448 70560 7448 0 _0124_
rlabel metal3 64288 6664 64288 6664 0 _0125_
rlabel metal2 65800 5936 65800 5936 0 _0126_
rlabel metal2 69608 7112 69608 7112 0 _0127_
rlabel metal2 13944 28224 13944 28224 0 _0128_
rlabel metal3 74816 6552 74816 6552 0 _0129_
rlabel metal2 76888 7840 76888 7840 0 _0130_
rlabel metal3 77336 11256 77336 11256 0 _0131_
rlabel metal2 72240 9688 72240 9688 0 _0132_
rlabel metal2 69496 10304 69496 10304 0 _0133_
rlabel metal3 68936 10360 68936 10360 0 _0134_
rlabel metal2 74760 10976 74760 10976 0 _0135_
rlabel metal2 75880 9464 75880 9464 0 _0136_
rlabel metal3 74312 10584 74312 10584 0 _0137_
rlabel metal2 71848 10640 71848 10640 0 _0138_
rlabel metal2 14056 27328 14056 27328 0 _0139_
rlabel metal3 74200 10472 74200 10472 0 _0140_
rlabel metal2 76440 10640 76440 10640 0 _0141_
rlabel metal3 75320 11368 75320 11368 0 _0142_
rlabel metal2 77448 11256 77448 11256 0 _0143_
rlabel metal3 72800 12264 72800 12264 0 _0144_
rlabel metal2 67704 14560 67704 14560 0 _0145_
rlabel metal2 61320 13944 61320 13944 0 _0146_
rlabel metal2 59640 14868 59640 14868 0 _0147_
rlabel metal2 59528 17248 59528 17248 0 _0148_
rlabel metal3 58744 19208 58744 19208 0 _0149_
rlabel metal2 14168 30184 14168 30184 0 _0150_
rlabel metal2 57680 18648 57680 18648 0 _0151_
rlabel metal3 57232 19320 57232 19320 0 _0152_
rlabel metal2 55608 19992 55608 19992 0 _0153_
rlabel metal2 53088 20664 53088 20664 0 _0154_
rlabel metal2 64792 16800 64792 16800 0 _0155_
rlabel metal3 68488 16856 68488 16856 0 _0156_
rlabel metal2 68432 13160 68432 13160 0 _0157_
rlabel metal3 68992 15288 68992 15288 0 _0158_
rlabel metal2 76552 10304 76552 10304 0 _0159_
rlabel metal2 14952 31248 14952 31248 0 _0160_
rlabel metal3 76272 10360 76272 10360 0 _0161_
rlabel metal2 75040 14056 75040 14056 0 _0162_
rlabel metal3 77224 15400 77224 15400 0 _0163_
rlabel metal2 77840 8344 77840 8344 0 _0164_
rlabel metal2 77448 12152 77448 12152 0 _0165_
rlabel metal3 76160 6104 76160 6104 0 _0166_
rlabel metal2 75320 6720 75320 6720 0 _0167_
rlabel metal3 73976 4536 73976 4536 0 _0168_
rlabel metal3 59864 4312 59864 4312 0 _0169_
rlabel metal2 72072 4368 72072 4368 0 _0170_
rlabel metal3 19992 25592 19992 25592 0 _0171_
rlabel metal2 67704 5040 67704 5040 0 _0172_
rlabel metal2 72408 4256 72408 4256 0 _0173_
rlabel metal2 71568 5208 71568 5208 0 _0174_
rlabel metal3 72296 5880 72296 5880 0 _0175_
rlabel metal2 69720 6216 69720 6216 0 _0176_
rlabel metal3 69216 6664 69216 6664 0 _0177_
rlabel metal2 67704 5880 67704 5880 0 _0178_
rlabel metal2 72408 6160 72408 6160 0 _0179_
rlabel metal3 73864 5768 73864 5768 0 _0180_
rlabel metal2 75992 7112 75992 7112 0 _0181_
rlabel metal3 20216 25480 20216 25480 0 _0182_
rlabel metal2 72968 9744 72968 9744 0 _0183_
rlabel metal2 73416 10024 73416 10024 0 _0184_
rlabel metal2 73640 9464 73640 9464 0 _0185_
rlabel metal2 71400 7952 71400 7952 0 _0186_
rlabel metal2 70504 11480 70504 11480 0 _0187_
rlabel metal3 70000 12040 70000 12040 0 _0188_
rlabel metal2 71344 12264 71344 12264 0 _0189_
rlabel metal2 71176 12208 71176 12208 0 _0190_
rlabel metal2 71176 8176 71176 8176 0 _0191_
rlabel metal3 72408 8232 72408 8232 0 _0192_
rlabel metal3 16800 29624 16800 29624 0 _0193_
rlabel metal3 75096 8232 75096 8232 0 _0194_
rlabel metal3 76048 8344 76048 8344 0 _0195_
rlabel metal2 77168 13608 77168 13608 0 _0196_
rlabel metal2 70392 15120 70392 15120 0 _0197_
rlabel metal2 70168 17640 70168 17640 0 _0198_
rlabel metal2 62104 18032 62104 18032 0 _0199_
rlabel metal2 60984 13776 60984 13776 0 _0200_
rlabel metal3 61096 17528 61096 17528 0 _0201_
rlabel metal3 60536 18424 60536 18424 0 _0202_
rlabel metal2 60088 20888 60088 20888 0 _0203_
rlabel metal2 19320 24416 19320 24416 0 _0204_
rlabel metal3 59192 20664 59192 20664 0 _0205_
rlabel metal3 59192 20888 59192 20888 0 _0206_
rlabel metal2 57960 21224 57960 21224 0 _0207_
rlabel metal2 60200 19320 60200 19320 0 _0208_
rlabel metal2 59864 20496 59864 20496 0 _0209_
rlabel metal2 61936 19208 61936 19208 0 _0210_
rlabel metal2 77784 18200 77784 18200 0 _0211_
rlabel metal3 76440 13160 76440 13160 0 _0212_
rlabel metal3 76440 13496 76440 13496 0 _0213_
rlabel metal2 8344 18592 8344 18592 0 _0214_
rlabel metal2 77616 14504 77616 14504 0 _0215_
rlabel metal2 73864 18424 73864 18424 0 _0216_
rlabel metal2 70448 8344 70448 8344 0 _0217_
rlabel metal3 72968 9016 72968 9016 0 _0218_
rlabel metal2 73584 17416 73584 17416 0 _0219_
rlabel metal2 75544 7840 75544 7840 0 _0220_
rlabel metal3 75880 9016 75880 9016 0 _0221_
rlabel metal2 76944 13384 76944 13384 0 _0222_
rlabel metal2 72128 4088 72128 4088 0 _0223_
rlabel metal2 72352 16072 72352 16072 0 _0224_
rlabel metal2 10696 22288 10696 22288 0 _0225_
rlabel metal2 68376 4816 68376 4816 0 _0226_
rlabel metal2 67760 3752 67760 3752 0 _0227_
rlabel metal2 68264 6608 68264 6608 0 _0228_
rlabel metal2 68040 18816 68040 18816 0 _0229_
rlabel metal2 63672 19656 63672 19656 0 _0230_
rlabel metal3 68488 19096 68488 19096 0 _0231_
rlabel metal2 71288 19600 71288 19600 0 _0232_
rlabel metal2 67704 6384 67704 6384 0 _0233_
rlabel metal2 66136 20832 66136 20832 0 _0234_
rlabel metal2 67592 21168 67592 21168 0 _0235_
rlabel metal2 20216 22904 20216 22904 0 _0236_
rlabel metal3 70280 20664 70280 20664 0 _0237_
rlabel metal2 72520 18032 72520 18032 0 _0238_
rlabel metal2 74088 16072 74088 16072 0 _0239_
rlabel metal2 71288 15008 71288 15008 0 _0240_
rlabel metal3 72632 13832 72632 13832 0 _0241_
rlabel metal2 67816 6104 67816 6104 0 _0242_
rlabel metal3 69216 13608 69216 13608 0 _0243_
rlabel metal2 67480 14000 67480 14000 0 _0244_
rlabel metal3 71008 14504 71008 14504 0 _0245_
rlabel metal3 72744 14616 72744 14616 0 _0246_
rlabel metal2 17640 30632 17640 30632 0 _0247_
rlabel metal2 73976 14868 73976 14868 0 _0248_
rlabel metal3 76552 16072 76552 16072 0 _0249_
rlabel metal3 76440 17640 76440 17640 0 _0250_
rlabel metal3 76272 17752 76272 17752 0 _0251_
rlabel metal3 71456 18424 71456 18424 0 _0252_
rlabel metal2 71512 17528 71512 17528 0 _0253_
rlabel metal2 71064 17752 71064 17752 0 _0254_
rlabel metal2 70056 19320 70056 19320 0 _0255_
rlabel metal2 61656 20720 61656 20720 0 _0256_
rlabel metal2 60704 21560 60704 21560 0 _0257_
rlabel metal2 16968 31472 16968 31472 0 _0258_
rlabel metal2 70056 17528 70056 17528 0 _0259_
rlabel metal2 68824 29232 68824 29232 0 _0260_
rlabel metal2 76720 19992 76720 19992 0 _0261_
rlabel metal2 74648 20048 74648 20048 0 _0262_
rlabel metal3 71904 13720 71904 13720 0 _0263_
rlabel metal2 73640 14448 73640 14448 0 _0264_
rlabel metal2 73024 13720 73024 13720 0 _0265_
rlabel metal2 73304 19824 73304 19824 0 _0266_
rlabel metal2 73752 16240 73752 16240 0 _0267_
rlabel metal2 17864 33152 17864 33152 0 _0268_
rlabel metal2 75208 20664 75208 20664 0 _0269_
rlabel metal3 70560 20328 70560 20328 0 _0270_
rlabel metal2 72184 21336 72184 21336 0 _0271_
rlabel metal4 65688 21784 65688 21784 0 _0272_
rlabel metal3 65352 18424 65352 18424 0 _0273_
rlabel metal2 70616 22736 70616 22736 0 _0274_
rlabel metal2 60648 23240 60648 23240 0 _0275_
rlabel metal3 59640 23016 59640 23016 0 _0276_
rlabel metal2 71176 22456 71176 22456 0 _0277_
rlabel metal3 72912 23128 72912 23128 0 _0278_
rlabel metal2 19488 29624 19488 29624 0 _0279_
rlabel metal2 67480 22568 67480 22568 0 _0280_
rlabel metal3 65912 22344 65912 22344 0 _0281_
rlabel metal2 66136 23408 66136 23408 0 _0282_
rlabel metal3 70896 22456 70896 22456 0 _0283_
rlabel metal2 76776 22008 76776 22008 0 _0284_
rlabel metal3 76496 22232 76496 22232 0 _0285_
rlabel metal2 66920 20664 66920 20664 0 _0286_
rlabel metal2 71176 20496 71176 20496 0 _0287_
rlabel metal3 70392 21000 70392 21000 0 _0288_
rlabel metal2 74648 22008 74648 22008 0 _0289_
rlabel metal2 18648 31556 18648 31556 0 _0290_
rlabel metal3 76552 20888 76552 20888 0 _0291_
rlabel metal2 74760 20272 74760 20272 0 _0292_
rlabel metal3 74872 19768 74872 19768 0 _0293_
rlabel metal2 74200 27440 74200 27440 0 _0294_
rlabel metal3 78344 26936 78344 26936 0 _0295_
rlabel metal3 75152 27944 75152 27944 0 _0296_
rlabel metal2 73752 18424 73752 18424 0 _0297_
rlabel metal2 77784 17640 77784 17640 0 _0298_
rlabel metal2 76440 27664 76440 27664 0 _0299_
rlabel metal2 70056 29064 70056 29064 0 _0300_
rlabel metal2 18872 32872 18872 32872 0 _0301_
rlabel metal3 64120 30184 64120 30184 0 _0302_
rlabel metal3 58632 21560 58632 21560 0 _0303_
rlabel metal2 52472 30240 52472 30240 0 _0304_
rlabel metal2 60648 29736 60648 29736 0 _0305_
rlabel metal2 51016 30744 51016 30744 0 _0306_
rlabel metal2 61880 20104 61880 20104 0 _0307_
rlabel metal2 62272 30744 62272 30744 0 _0308_
rlabel metal2 61824 31528 61824 31528 0 _0309_
rlabel metal2 61432 30632 61432 30632 0 _0310_
rlabel metal2 19768 32984 19768 32984 0 _0311_
rlabel metal3 68992 30072 68992 30072 0 _0312_
rlabel metal2 67144 30576 67144 30576 0 _0313_
rlabel metal2 62664 31248 62664 31248 0 _0314_
rlabel metal2 67592 31360 67592 31360 0 _0315_
rlabel metal3 70728 20552 70728 20552 0 _0316_
rlabel metal2 71064 21504 71064 21504 0 _0317_
rlabel metal2 75880 25312 75880 25312 0 _0318_
rlabel metal2 77112 21952 77112 21952 0 _0319_
rlabel metal2 76328 24640 76328 24640 0 _0320_
rlabel metal2 67312 22344 67312 22344 0 _0321_
rlabel metal2 66920 22680 66920 22680 0 _0322_
rlabel metal2 73528 24192 73528 24192 0 _0323_
rlabel metal2 71512 22456 71512 22456 0 _0324_
rlabel metal2 72184 23632 72184 23632 0 _0325_
rlabel metal3 57848 22904 57848 22904 0 _0326_
rlabel metal2 60312 22848 60312 22848 0 _0327_
rlabel metal2 61880 23632 61880 23632 0 _0328_
rlabel metal2 57848 24696 57848 24696 0 _0329_
rlabel metal3 56784 25704 56784 25704 0 _0330_
rlabel metal2 57960 24248 57960 24248 0 _0331_
rlabel metal3 15176 31192 15176 31192 0 _0332_
rlabel metal3 60088 23912 60088 23912 0 _0333_
rlabel metal3 69440 24808 69440 24808 0 _0334_
rlabel metal2 67704 25424 67704 25424 0 _0335_
rlabel metal2 66136 25648 66136 25648 0 _0336_
rlabel metal2 66808 25872 66808 25872 0 _0337_
rlabel metal3 69272 25368 69272 25368 0 _0338_
rlabel metal2 71904 24696 71904 24696 0 _0339_
rlabel metal2 73640 24080 73640 24080 0 _0340_
rlabel metal2 76440 23912 76440 23912 0 _0341_
rlabel metal2 76888 24864 76888 24864 0 _0342_
rlabel metal2 15848 30576 15848 30576 0 _0343_
rlabel metal2 77448 25928 77448 25928 0 _0344_
rlabel metal3 75824 20776 75824 20776 0 _0345_
rlabel metal3 74088 26600 74088 26600 0 _0346_
rlabel metal2 77672 28168 77672 28168 0 _0347_
rlabel metal2 76552 28112 76552 28112 0 _0348_
rlabel metal2 72744 29288 72744 29288 0 _0349_
rlabel metal2 66920 31136 66920 31136 0 _0350_
rlabel metal2 67368 31360 67368 31360 0 _0351_
rlabel metal2 65576 31248 65576 31248 0 _0352_
rlabel metal2 13776 31192 13776 31192 0 _0353_
rlabel metal2 72016 30968 72016 30968 0 _0354_
rlabel metal2 70728 30688 70728 30688 0 _0355_
rlabel metal3 74928 26264 74928 26264 0 _0356_
rlabel metal3 76832 25928 76832 25928 0 _0357_
rlabel metal2 67928 25816 67928 25816 0 _0358_
rlabel metal3 67424 26040 67424 26040 0 _0359_
rlabel metal3 70448 26264 70448 26264 0 _0360_
rlabel metal2 69272 24696 69272 24696 0 _0361_
rlabel metal2 69944 26320 69944 26320 0 _0362_
rlabel metal2 62776 25816 62776 25816 0 _0363_
rlabel metal2 54040 3864 54040 3864 0 _0364_
rlabel metal2 64904 27216 64904 27216 0 _0365_
rlabel metal2 67592 28280 67592 28280 0 _0366_
rlabel metal3 64400 26488 64400 26488 0 _0367_
rlabel metal2 62944 27272 62944 27272 0 _0368_
rlabel metal3 58800 24920 58800 24920 0 _0369_
rlabel metal2 61544 25928 61544 25928 0 _0370_
rlabel metal2 58520 28112 58520 28112 0 _0371_
rlabel via2 56840 29400 56840 29400 0 _0372_
rlabel metal2 57064 27552 57064 27552 0 _0373_
rlabel metal2 57288 26964 57288 26964 0 _0374_
rlabel metal3 9576 20664 9576 20664 0 _0375_
rlabel metal2 58296 27216 58296 27216 0 _0376_
rlabel metal3 60424 26936 60424 26936 0 _0377_
rlabel metal3 62552 26264 62552 26264 0 _0378_
rlabel metal3 68936 27048 68936 27048 0 _0379_
rlabel metal2 70392 26656 70392 26656 0 _0380_
rlabel metal2 70504 26768 70504 26768 0 _0381_
rlabel metal3 72240 27048 72240 27048 0 _0382_
rlabel metal2 72296 25088 72296 25088 0 _0383_
rlabel metal2 73304 25144 73304 25144 0 _0384_
rlabel metal2 72520 26264 72520 26264 0 _0385_
rlabel metal2 10136 27944 10136 27944 0 _0386_
rlabel metal2 73864 26656 73864 26656 0 _0387_
rlabel metal2 77840 27944 77840 27944 0 _0388_
rlabel metal3 77000 27272 77000 27272 0 _0389_
rlabel metal2 77896 29568 77896 29568 0 _0390_
rlabel metal3 76160 25704 76160 25704 0 _0391_
rlabel metal2 74312 29904 74312 29904 0 _0392_
rlabel metal2 74536 29568 74536 29568 0 _0393_
rlabel metal3 74928 30296 74928 30296 0 _0394_
rlabel metal2 72128 31640 72128 31640 0 _0395_
rlabel metal2 70280 31248 70280 31248 0 _0396_
rlabel metal2 11368 27328 11368 27328 0 _0397_
rlabel metal3 63000 26824 63000 26824 0 _0398_
rlabel metal3 63504 27048 63504 27048 0 _0399_
rlabel metal2 63952 27272 63952 27272 0 _0400_
rlabel metal3 58800 27608 58800 27608 0 _0401_
rlabel metal2 60200 28504 60200 28504 0 _0402_
rlabel metal3 59080 29400 59080 29400 0 _0403_
rlabel metal2 54824 30464 54824 30464 0 _0404_
rlabel metal3 57400 29288 57400 29288 0 _0405_
rlabel metal2 59752 28560 59752 28560 0 _0406_
rlabel metal2 10472 28224 10472 28224 0 _0407_
rlabel metal3 62832 27944 62832 27944 0 _0408_
rlabel metal2 65128 29008 65128 29008 0 _0409_
rlabel metal2 66696 28560 66696 28560 0 _0410_
rlabel metal3 68880 28504 68880 28504 0 _0411_
rlabel metal2 68936 26264 68936 26264 0 _0412_
rlabel metal2 69608 27104 69608 27104 0 _0413_
rlabel metal3 70560 28616 70560 28616 0 _0414_
rlabel metal2 71400 27608 71400 27608 0 _0415_
rlabel metal2 71512 28392 71512 28392 0 _0416_
rlabel metal2 72016 30184 72016 30184 0 _0417_
rlabel metal3 11200 30184 11200 30184 0 _0418_
rlabel metal3 77168 30072 77168 30072 0 _0419_
rlabel metal2 75488 30856 75488 30856 0 _0420_
rlabel metal2 74312 31892 74312 31892 0 _0421_
rlabel metal2 72296 31304 72296 31304 0 _0422_
rlabel metal3 72688 31192 72688 31192 0 _0423_
rlabel metal3 75488 31192 75488 31192 0 _0424_
rlabel metal2 73416 32256 73416 32256 0 _0425_
rlabel metal2 74760 32984 74760 32984 0 _0426_
rlabel metal2 71680 29624 71680 29624 0 _0427_
rlabel metal2 21672 23184 21672 23184 0 _0428_
rlabel metal2 64288 29400 64288 29400 0 _0429_
rlabel metal2 63840 31528 63840 31528 0 _0430_
rlabel metal3 64568 31528 64568 31528 0 _0431_
rlabel metal2 54880 31640 54880 31640 0 _0432_
rlabel metal3 54768 31976 54768 31976 0 _0433_
rlabel metal2 55608 31080 55608 31080 0 _0434_
rlabel metal3 58296 31640 58296 31640 0 _0435_
rlabel metal2 57512 30688 57512 30688 0 _0436_
rlabel metal2 58408 30520 58408 30520 0 _0437_
rlabel metal3 59024 31752 59024 31752 0 _0438_
rlabel metal3 21224 24024 21224 24024 0 _0439_
rlabel metal3 58408 31976 58408 31976 0 _0440_
rlabel metal2 60424 32256 60424 32256 0 _0441_
rlabel metal3 60816 32536 60816 32536 0 _0442_
rlabel metal2 61992 28336 61992 28336 0 _0443_
rlabel metal2 61544 29792 61544 29792 0 _0444_
rlabel metal2 63280 31752 63280 31752 0 _0445_
rlabel metal2 63112 32984 63112 32984 0 _0446_
rlabel metal2 63112 33544 63112 33544 0 _0447_
rlabel metal2 63896 32536 63896 32536 0 _0448_
rlabel metal3 64848 33320 64848 33320 0 _0449_
rlabel metal2 12600 28504 12600 28504 0 _0450_
rlabel metal2 69440 28840 69440 28840 0 _0451_
rlabel metal2 70672 29176 70672 29176 0 _0452_
rlabel metal2 67144 33040 67144 33040 0 _0453_
rlabel metal2 70616 32816 70616 32816 0 _0454_
rlabel metal2 70560 33320 70560 33320 0 _0455_
rlabel metal3 70448 30968 70448 30968 0 _0456_
rlabel metal2 68264 31416 68264 31416 0 _0457_
rlabel metal3 77000 31864 77000 31864 0 _0458_
rlabel metal3 74368 31640 74368 31640 0 _0459_
rlabel metal2 70168 30688 70168 30688 0 _0460_
rlabel metal2 20664 22848 20664 22848 0 _0461_
rlabel metal3 70224 31192 70224 31192 0 _0462_
rlabel metal2 70280 32648 70280 32648 0 _0463_
rlabel metal2 71120 33432 71120 33432 0 _0464_
rlabel metal2 69720 34664 69720 34664 0 _0465_
rlabel metal3 61096 33096 61096 33096 0 _0466_
rlabel metal2 57960 34160 57960 34160 0 _0467_
rlabel metal2 59752 34608 59752 34608 0 _0468_
rlabel metal2 51464 31248 51464 31248 0 _0469_
rlabel metal2 54992 30968 54992 30968 0 _0470_
rlabel metal3 6832 15176 6832 15176 0 _0471_
rlabel metal2 54320 31192 54320 31192 0 _0472_
rlabel metal2 51464 32760 51464 32760 0 _0473_
rlabel metal2 53816 33040 53816 33040 0 _0474_
rlabel metal2 54936 33600 54936 33600 0 _0475_
rlabel metal2 59192 35168 59192 35168 0 _0476_
rlabel metal2 60648 35392 60648 35392 0 _0477_
rlabel metal3 64120 34104 64120 34104 0 _0478_
rlabel metal2 62776 34664 62776 34664 0 _0479_
rlabel metal3 63616 34776 63616 34776 0 _0480_
rlabel metal2 69496 34888 69496 34888 0 _0481_
rlabel metal2 30744 22176 30744 22176 0 _0482_
rlabel metal2 72296 34888 72296 34888 0 _0483_
rlabel metal2 71848 33936 71848 33936 0 _0484_
rlabel metal3 71960 34776 71960 34776 0 _0485_
rlabel metal2 70840 35168 70840 35168 0 _0486_
rlabel metal2 61880 35616 61880 35616 0 _0487_
rlabel metal2 55272 34440 55272 34440 0 _0488_
rlabel metal2 56112 32760 56112 32760 0 _0489_
rlabel metal2 53928 33544 53928 33544 0 _0490_
rlabel metal3 57176 33320 57176 33320 0 _0491_
rlabel metal2 20440 20664 20440 20664 0 _0492_
rlabel metal2 55720 34216 55720 34216 0 _0493_
rlabel metal2 56112 34888 56112 34888 0 _0494_
rlabel metal3 58240 35560 58240 35560 0 _0495_
rlabel metal2 57064 35224 57064 35224 0 _0496_
rlabel metal3 59752 35672 59752 35672 0 _0497_
rlabel metal2 65016 35168 65016 35168 0 _0498_
rlabel metal2 66696 35168 66696 35168 0 _0499_
rlabel metal2 65576 35280 65576 35280 0 _0500_
rlabel metal2 65016 34608 65016 34608 0 _0501_
rlabel metal3 65184 35560 65184 35560 0 _0502_
rlabel metal2 12152 27048 12152 27048 0 _0503_
rlabel metal2 66864 35672 66864 35672 0 _0504_
rlabel metal2 60200 34944 60200 34944 0 _0505_
rlabel metal2 59416 35056 59416 35056 0 _0506_
rlabel metal2 58016 32760 58016 32760 0 _0507_
rlabel metal2 58464 32760 58464 32760 0 _0508_
rlabel metal2 58296 34888 58296 34888 0 _0509_
rlabel metal2 60088 36120 60088 36120 0 _0510_
rlabel metal2 18984 35224 18984 35224 0 _0511_
rlabel metal2 10360 30240 10360 30240 0 _0512_
rlabel metal3 23352 28056 23352 28056 0 _0513_
rlabel metal2 23128 27384 23128 27384 0 _0514_
rlabel metal2 13888 30968 13888 30968 0 _0515_
rlabel metal3 13720 32424 13720 32424 0 _0516_
rlabel metal2 17752 35336 17752 35336 0 _0517_
rlabel metal2 12040 35728 12040 35728 0 _0518_
rlabel metal2 11704 35672 11704 35672 0 _0519_
rlabel metal3 12600 35672 12600 35672 0 _0520_
rlabel metal2 12712 35280 12712 35280 0 _0521_
rlabel metal3 17360 34328 17360 34328 0 _0522_
rlabel metal2 10864 25480 10864 25480 0 _0523_
rlabel metal2 8344 27384 8344 27384 0 _0524_
rlabel metal2 55384 3080 55384 3080 0 _0525_
rlabel metal3 7000 21560 7000 21560 0 _0526_
rlabel metal2 7672 27104 7672 27104 0 _0527_
rlabel metal3 9072 31752 9072 31752 0 _0528_
rlabel metal3 11592 29624 11592 29624 0 _0529_
rlabel metal2 8904 31472 8904 31472 0 _0530_
rlabel metal2 19936 22120 19936 22120 0 _0531_
rlabel metal3 21168 20888 21168 20888 0 _0532_
rlabel metal3 18312 22232 18312 22232 0 _0533_
rlabel metal2 17752 21112 17752 21112 0 _0534_
rlabel metal2 9240 15512 9240 15512 0 _0535_
rlabel metal3 16856 19208 16856 19208 0 _0536_
rlabel metal2 16408 22680 16408 22680 0 _0537_
rlabel metal2 14952 24640 14952 24640 0 _0538_
rlabel metal2 10360 25928 10360 25928 0 _0539_
rlabel metal2 11256 25032 11256 25032 0 _0540_
rlabel metal2 13664 23912 13664 23912 0 _0541_
rlabel metal3 14056 24696 14056 24696 0 _0542_
rlabel metal2 9912 30016 9912 30016 0 _0543_
rlabel metal3 11760 33320 11760 33320 0 _0544_
rlabel metal3 13160 31192 13160 31192 0 _0545_
rlabel metal2 13160 32816 13160 32816 0 _0546_
rlabel metal3 15400 34888 15400 34888 0 _0547_
rlabel metal2 17304 35728 17304 35728 0 _0548_
rlabel metal3 15624 35560 15624 35560 0 _0549_
rlabel metal2 16744 35952 16744 35952 0 _0550_
rlabel metal3 11368 26264 11368 26264 0 _0551_
rlabel metal2 5096 29008 5096 29008 0 _0552_
rlabel metal2 3192 8232 3192 8232 0 _0553_
rlabel metal2 4424 24864 4424 24864 0 _0554_
rlabel metal2 13832 26544 13832 26544 0 _0555_
rlabel metal2 3640 23128 3640 23128 0 _0556_
rlabel metal3 4760 27048 4760 27048 0 _0557_
rlabel metal2 4536 28280 4536 28280 0 _0558_
rlabel metal2 4200 31248 4200 31248 0 _0559_
rlabel metal2 7000 29848 7000 29848 0 _0560_
rlabel metal2 16520 23632 16520 23632 0 _0561_
rlabel metal3 7560 28616 7560 28616 0 _0562_
rlabel metal2 19544 19320 19544 19320 0 _0563_
rlabel metal2 18144 19320 18144 19320 0 _0564_
rlabel metal3 7616 23128 7616 23128 0 _0565_
rlabel metal2 17528 18032 17528 18032 0 _0566_
rlabel metal3 44072 13216 44072 13216 0 _0567_
rlabel metal2 68264 12768 68264 12768 0 _0568_
rlabel metal3 18872 17864 18872 17864 0 _0569_
rlabel via2 7112 23016 7112 23016 0 _0570_
rlabel metal2 6664 24192 6664 24192 0 _0571_
rlabel metal2 7448 24248 7448 24248 0 _0572_
rlabel metal2 8120 24472 8120 24472 0 _0573_
rlabel metal3 10808 24024 10808 24024 0 _0574_
rlabel metal2 7672 24584 7672 24584 0 _0575_
rlabel metal2 6160 25592 6160 25592 0 _0576_
rlabel metal2 7056 28616 7056 28616 0 _0577_
rlabel metal2 6776 30016 6776 30016 0 _0578_
rlabel metal2 6776 29232 6776 29232 0 _0579_
rlabel metal3 5768 30968 5768 30968 0 _0580_
rlabel metal2 7280 24136 7280 24136 0 _0581_
rlabel metal3 6552 26264 6552 26264 0 _0582_
rlabel metal2 49672 7840 49672 7840 0 _0583_
rlabel metal3 2408 21672 2408 21672 0 _0584_
rlabel metal3 3416 23688 3416 23688 0 _0585_
rlabel metal3 4256 23016 4256 23016 0 _0586_
rlabel metal3 3416 23800 3416 23800 0 _0587_
rlabel metal3 4424 25592 4424 25592 0 _0588_
rlabel metal2 4088 26656 4088 26656 0 _0589_
rlabel metal2 4200 27496 4200 27496 0 _0590_
rlabel metal2 6552 24360 6552 24360 0 _0591_
rlabel metal3 4144 28392 4144 28392 0 _0592_
rlabel metal2 8344 19712 8344 19712 0 _0593_
rlabel metal2 9576 20356 9576 20356 0 _0594_
rlabel metal3 12096 17864 12096 17864 0 _0595_
rlabel metal3 12992 20552 12992 20552 0 _0596_
rlabel metal3 17752 18424 17752 18424 0 _0597_
rlabel metal2 13944 16128 13944 16128 0 _0598_
rlabel metal3 18480 19320 18480 19320 0 _0599_
rlabel metal2 15064 19712 15064 19712 0 _0600_
rlabel metal2 17696 16856 17696 16856 0 _0601_
rlabel metal2 19040 12152 19040 12152 0 _0602_
rlabel metal3 67536 13944 67536 13944 0 _0603_
rlabel metal2 19152 15512 19152 15512 0 _0604_
rlabel metal2 15176 19376 15176 19376 0 _0605_
rlabel metal2 13720 21112 13720 21112 0 _0606_
rlabel metal2 6664 27776 6664 27776 0 _0607_
rlabel metal2 4984 30968 4984 30968 0 _0608_
rlabel metal2 5992 31192 5992 31192 0 _0609_
rlabel metal2 7224 32816 7224 32816 0 _0610_
rlabel metal3 9688 30856 9688 30856 0 _0611_
rlabel metal2 9800 30576 9800 30576 0 _0612_
rlabel metal2 6776 33712 6776 33712 0 _0613_
rlabel metal2 8232 33712 8232 33712 0 _0614_
rlabel metal2 9912 32928 9912 32928 0 _0615_
rlabel metal2 7672 32928 7672 32928 0 _0616_
rlabel metal2 20216 33936 20216 33936 0 _0617_
rlabel metal2 14224 34216 14224 34216 0 _0618_
rlabel metal3 11592 33880 11592 33880 0 _0619_
rlabel metal2 21224 34160 21224 34160 0 _0620_
rlabel metal2 22456 34496 22456 34496 0 _0621_
rlabel metal2 21560 35392 21560 35392 0 _0622_
rlabel metal3 22904 35672 22904 35672 0 _0623_
rlabel metal3 19040 35672 19040 35672 0 _0624_
rlabel metal3 10192 34888 10192 34888 0 _0625_
rlabel metal3 12600 34216 12600 34216 0 _0626_
rlabel metal3 15904 35112 15904 35112 0 _0627_
rlabel metal2 23128 35336 23128 35336 0 _0628_
rlabel metal2 24304 35672 24304 35672 0 _0629_
rlabel metal2 4704 26264 4704 26264 0 _0630_
rlabel metal2 5544 26488 5544 26488 0 _0631_
rlabel metal2 27496 17752 27496 17752 0 _0632_
rlabel metal2 26824 28168 26824 28168 0 _0633_
rlabel metal3 25200 28728 25200 28728 0 _0634_
rlabel metal2 23912 29400 23912 29400 0 _0635_
rlabel metal2 5320 28112 5320 28112 0 _0636_
rlabel metal2 6160 27832 6160 27832 0 _0637_
rlabel metal2 5432 28952 5432 28952 0 _0638_
rlabel metal2 3864 22624 3864 22624 0 _0639_
rlabel metal2 4312 23632 4312 23632 0 _0640_
rlabel metal2 9352 22624 9352 22624 0 _0641_
rlabel metal2 10192 20552 10192 20552 0 _0642_
rlabel metal2 10192 18984 10192 18984 0 _0643_
rlabel metal3 9296 19208 9296 19208 0 _0644_
rlabel metal2 8120 22288 8120 22288 0 _0645_
rlabel metal2 4088 21896 4088 21896 0 _0646_
rlabel metal2 4648 21168 4648 21168 0 _0647_
rlabel metal3 6216 21672 6216 21672 0 _0648_
rlabel metal2 7672 22064 7672 22064 0 _0649_
rlabel metal3 9016 22456 9016 22456 0 _0650_
rlabel metal3 11816 23128 11816 23128 0 _0651_
rlabel metal2 14840 20496 14840 20496 0 _0652_
rlabel metal2 12824 22624 12824 22624 0 _0653_
rlabel metal2 10136 18368 10136 18368 0 _0654_
rlabel metal2 13608 18088 13608 18088 0 _0655_
rlabel metal2 21000 18032 21000 18032 0 _0656_
rlabel metal2 18256 15624 18256 15624 0 _0657_
rlabel metal2 17976 16464 17976 16464 0 _0658_
rlabel metal3 19936 16856 19936 16856 0 _0659_
rlabel metal2 17640 14280 17640 14280 0 _0660_
rlabel metal3 21896 12824 21896 12824 0 _0661_
rlabel metal3 19544 12824 19544 12824 0 _0662_
rlabel metal2 22232 16912 22232 16912 0 _0663_
rlabel metal2 22176 18312 22176 18312 0 _0664_
rlabel metal2 15064 22176 15064 22176 0 _0665_
rlabel metal2 15064 28672 15064 28672 0 _0666_
rlabel metal2 22960 30856 22960 30856 0 _0667_
rlabel metal2 24696 31304 24696 31304 0 _0668_
rlabel metal2 6328 31472 6328 31472 0 _0669_
rlabel metal2 5656 31808 5656 31808 0 _0670_
rlabel metal2 24584 31584 24584 31584 0 _0671_
rlabel metal2 25256 34888 25256 34888 0 _0672_
rlabel metal3 25088 34104 25088 34104 0 _0673_
rlabel metal2 26488 33992 26488 33992 0 _0674_
rlabel metal2 26264 34608 26264 34608 0 _0675_
rlabel metal3 29176 35672 29176 35672 0 _0676_
rlabel metal3 24640 35560 24640 35560 0 _0677_
rlabel metal3 24864 36344 24864 36344 0 _0678_
rlabel metal3 27888 36232 27888 36232 0 _0679_
rlabel metal2 28840 35280 28840 35280 0 _0680_
rlabel metal2 26488 35728 26488 35728 0 _0681_
rlabel metal3 27160 35896 27160 35896 0 _0682_
rlabel metal3 30212 35896 30212 35896 0 _0683_
rlabel metal3 27776 33096 27776 33096 0 _0684_
rlabel metal2 23576 29568 23576 29568 0 _0685_
rlabel metal2 24080 30296 24080 30296 0 _0686_
rlabel metal2 9016 22232 9016 22232 0 _0687_
rlabel metal2 10136 21784 10136 21784 0 _0688_
rlabel metal2 27384 29176 27384 29176 0 _0689_
rlabel via2 27944 26824 27944 26824 0 _0690_
rlabel metal2 28840 20496 28840 20496 0 _0691_
rlabel metal2 28280 24192 28280 24192 0 _0692_
rlabel metal3 28280 27944 28280 27944 0 _0693_
rlabel metal3 29344 28504 29344 28504 0 _0694_
rlabel metal3 28728 27272 28728 27272 0 _0695_
rlabel metal2 28168 29400 28168 29400 0 _0696_
rlabel metal2 27496 30240 27496 30240 0 _0697_
rlabel metal3 13328 22344 13328 22344 0 _0698_
rlabel metal2 14560 22344 14560 22344 0 _0699_
rlabel metal2 25256 29120 25256 29120 0 _0700_
rlabel metal2 3528 18032 3528 18032 0 _0701_
rlabel metal2 3752 20552 3752 20552 0 _0702_
rlabel metal2 4872 19600 4872 19600 0 _0703_
rlabel metal2 9576 16072 9576 16072 0 _0704_
rlabel metal2 9800 17360 9800 17360 0 _0705_
rlabel metal2 6552 18480 6552 18480 0 _0706_
rlabel metal2 3192 15064 3192 15064 0 _0707_
rlabel metal3 3360 16856 3360 16856 0 _0708_
rlabel metal2 3864 17976 3864 17976 0 _0709_
rlabel metal2 4984 18088 4984 18088 0 _0710_
rlabel metal2 5824 19320 5824 19320 0 _0711_
rlabel metal2 6776 19544 6776 19544 0 _0712_
rlabel metal2 22288 17640 22288 17640 0 _0713_
rlabel metal2 24136 19152 24136 19152 0 _0714_
rlabel metal2 13272 16072 13272 16072 0 _0715_
rlabel metal3 11816 15176 11816 15176 0 _0716_
rlabel metal3 14812 15512 14812 15512 0 _0717_
rlabel metal3 20048 13720 20048 13720 0 _0718_
rlabel metal3 69664 20552 69664 20552 0 _0719_
rlabel metal2 18424 15148 18424 15148 0 _0720_
rlabel metal2 24024 14112 24024 14112 0 _0721_
rlabel metal2 20832 12936 20832 12936 0 _0722_
rlabel metal2 67424 7672 67424 7672 0 _0723_
rlabel metal2 64904 22848 64904 22848 0 _0724_
rlabel metal2 22568 13048 22568 13048 0 _0725_
rlabel metal2 23912 14112 23912 14112 0 _0726_
rlabel metal2 24808 16184 24808 16184 0 _0727_
rlabel metal2 24472 18144 24472 18144 0 _0728_
rlabel metal2 24976 29960 24976 29960 0 _0729_
rlabel metal2 26824 31080 26824 31080 0 _0730_
rlabel metal2 27608 32200 27608 32200 0 _0731_
rlabel metal3 29120 33320 29120 33320 0 _0732_
rlabel metal2 31304 34552 31304 34552 0 _0733_
rlabel metal2 24864 31752 24864 31752 0 _0734_
rlabel metal2 30296 34496 30296 34496 0 _0735_
rlabel metal2 31416 35336 31416 35336 0 _0736_
rlabel metal2 35000 36120 35000 36120 0 _0737_
rlabel metal3 33264 35672 33264 35672 0 _0738_
rlabel metal2 28784 29624 28784 29624 0 _0739_
rlabel metal2 26376 30576 26376 30576 0 _0740_
rlabel metal2 27720 31360 27720 31360 0 _0741_
rlabel metal3 5488 19432 5488 19432 0 _0742_
rlabel metal2 5936 17864 5936 17864 0 _0743_
rlabel metal2 6608 18200 6608 18200 0 _0744_
rlabel metal2 29624 27104 29624 27104 0 _0745_
rlabel metal3 69384 7560 69384 7560 0 _0746_
rlabel metal3 29400 22120 29400 22120 0 _0747_
rlabel metal2 27552 25704 27552 25704 0 _0748_
rlabel metal2 28280 22008 28280 22008 0 _0749_
rlabel metal2 27776 24920 27776 24920 0 _0750_
rlabel metal2 27720 25760 27720 25760 0 _0751_
rlabel metal2 27496 26544 27496 26544 0 _0752_
rlabel metal2 28504 27496 28504 27496 0 _0753_
rlabel metal2 31528 30240 31528 30240 0 _0754_
rlabel metal2 31248 31752 31248 31752 0 _0755_
rlabel metal2 24360 19040 24360 19040 0 _0756_
rlabel metal3 25536 19432 25536 19432 0 _0757_
rlabel metal3 26992 29960 26992 29960 0 _0758_
rlabel metal2 4424 16520 4424 16520 0 _0759_
rlabel metal2 4760 16632 4760 16632 0 _0760_
rlabel metal3 4200 16744 4200 16744 0 _0761_
rlabel metal2 7000 16800 7000 16800 0 _0762_
rlabel metal3 12152 15848 12152 15848 0 _0763_
rlabel metal2 11592 15792 11592 15792 0 _0764_
rlabel metal2 7784 16016 7784 16016 0 _0765_
rlabel metal2 3416 13440 3416 13440 0 _0766_
rlabel metal2 2856 11144 2856 11144 0 _0767_
rlabel metal2 3640 13328 3640 13328 0 _0768_
rlabel metal3 5152 16184 5152 16184 0 _0769_
rlabel metal2 6888 16856 6888 16856 0 _0770_
rlabel metal2 25424 15848 25424 15848 0 _0771_
rlabel metal2 24304 15848 24304 15848 0 _0772_
rlabel metal2 25816 16800 25816 16800 0 _0773_
rlabel metal3 13272 15848 13272 15848 0 _0774_
rlabel metal2 13832 13328 13832 13328 0 _0775_
rlabel metal2 24696 14728 24696 14728 0 _0776_
rlabel metal3 19768 11928 19768 11928 0 _0777_
rlabel metal2 20272 16184 20272 16184 0 _0778_
rlabel metal2 25032 12824 25032 12824 0 _0779_
rlabel metal2 18536 11480 18536 11480 0 _0780_
rlabel metal2 45304 9016 45304 9016 0 _0781_
rlabel metal2 67368 24304 67368 24304 0 _0782_
rlabel metal3 19880 10024 19880 10024 0 _0783_
rlabel metal2 25256 12600 25256 12600 0 _0784_
rlabel metal2 26264 14000 26264 14000 0 _0785_
rlabel metal2 27272 16464 27272 16464 0 _0786_
rlabel metal2 29344 29288 29344 29288 0 _0787_
rlabel metal2 30968 31108 30968 31108 0 _0788_
rlabel metal2 33880 32928 33880 32928 0 _0789_
rlabel metal2 35224 33712 35224 33712 0 _0790_
rlabel metal2 29512 33040 29512 33040 0 _0791_
rlabel metal2 28392 34160 28392 34160 0 _0792_
rlabel metal2 37464 35392 37464 35392 0 _0793_
rlabel metal2 36792 34328 36792 34328 0 _0794_
rlabel metal2 36232 34720 36232 34720 0 _0795_
rlabel metal3 37296 36456 37296 36456 0 _0796_
rlabel metal2 39480 35280 39480 35280 0 _0797_
rlabel metal2 46200 35224 46200 35224 0 _0798_
rlabel metal2 37688 33992 37688 33992 0 _0799_
rlabel metal3 37128 34776 37128 34776 0 _0800_
rlabel metal3 38164 34664 38164 34664 0 _0801_
rlabel via2 47208 35672 47208 35672 0 _0802_
rlabel metal2 41496 34440 41496 34440 0 _0803_
rlabel metal2 33768 32984 33768 32984 0 _0804_
rlabel metal2 34272 32760 34272 32760 0 _0805_
rlabel metal2 39760 34888 39760 34888 0 _0806_
rlabel metal2 31864 31640 31864 31640 0 _0807_
rlabel metal2 31752 31864 31752 31864 0 _0808_
rlabel metal3 37352 32424 37352 32424 0 _0809_
rlabel metal2 28840 29120 28840 29120 0 _0810_
rlabel metal2 7672 16296 7672 16296 0 _0811_
rlabel metal2 31080 26544 31080 26544 0 _0812_
rlabel metal3 64960 21784 64960 21784 0 _0813_
rlabel metal3 31304 27832 31304 27832 0 _0814_
rlabel metal2 31640 27720 31640 27720 0 _0815_
rlabel metal3 28896 25592 28896 25592 0 _0816_
rlabel metal3 30408 26264 30408 26264 0 _0817_
rlabel metal2 27832 22176 27832 22176 0 _0818_
rlabel metal2 29176 22904 29176 22904 0 _0819_
rlabel metal2 30520 26096 30520 26096 0 _0820_
rlabel metal2 31416 26712 31416 26712 0 _0821_
rlabel metal2 32424 28224 32424 28224 0 _0822_
rlabel metal2 32088 29008 32088 29008 0 _0823_
rlabel metal2 35560 29624 35560 29624 0 _0824_
rlabel metal2 26264 16800 26264 16800 0 _0825_
rlabel metal2 26824 16856 26824 16856 0 _0826_
rlabel metal2 33992 30296 33992 30296 0 _0827_
rlabel metal2 4144 12936 4144 12936 0 _0828_
rlabel metal3 5544 14392 5544 14392 0 _0829_
rlabel metal3 13328 14392 13328 14392 0 _0830_
rlabel metal2 12040 14000 12040 14000 0 _0831_
rlabel metal2 9912 14112 9912 14112 0 _0832_
rlabel metal2 4536 11760 4536 11760 0 _0833_
rlabel metal2 8176 12712 8176 12712 0 _0834_
rlabel metal3 6944 13608 6944 13608 0 _0835_
rlabel metal2 8680 14168 8680 14168 0 _0836_
rlabel metal3 20664 14392 20664 14392 0 _0837_
rlabel metal3 25312 13720 25312 13720 0 _0838_
rlabel metal2 28056 14056 28056 14056 0 _0839_
rlabel metal2 13776 11592 13776 11592 0 _0840_
rlabel metal2 14896 11144 14896 11144 0 _0841_
rlabel metal2 24920 11928 24920 11928 0 _0842_
rlabel metal2 22344 10864 22344 10864 0 _0843_
rlabel metal2 21672 13832 21672 13832 0 _0844_
rlabel metal3 23576 11368 23576 11368 0 _0845_
rlabel metal3 20496 9912 20496 9912 0 _0846_
rlabel metal2 48552 7616 48552 7616 0 _0847_
rlabel metal2 61880 27888 61880 27888 0 _0848_
rlabel metal2 23296 9576 23296 9576 0 _0849_
rlabel metal3 24696 11480 24696 11480 0 _0850_
rlabel metal2 25816 11704 25816 11704 0 _0851_
rlabel metal2 26712 12712 26712 12712 0 _0852_
rlabel metal2 33488 29960 33488 29960 0 _0853_
rlabel metal2 37128 31500 37128 31500 0 _0854_
rlabel metal2 40376 34552 40376 34552 0 _0855_
rlabel metal3 41720 34888 41720 34888 0 _0856_
rlabel metal2 45528 36176 45528 36176 0 _0857_
rlabel metal2 48776 35224 48776 35224 0 _0858_
rlabel metal3 44520 34216 44520 34216 0 _0859_
rlabel metal2 46088 35784 46088 35784 0 _0860_
rlabel metal2 42840 34552 42840 34552 0 _0861_
rlabel metal2 33824 28840 33824 28840 0 _0862_
rlabel metal3 33376 29512 33376 29512 0 _0863_
rlabel metal2 33992 29848 33992 29848 0 _0864_
rlabel metal3 35056 30184 35056 30184 0 _0865_
rlabel metal2 36176 30184 36176 30184 0 _0866_
rlabel metal2 39144 30576 39144 30576 0 _0867_
rlabel metal2 28056 15008 28056 15008 0 _0868_
rlabel metal2 28728 15008 28728 15008 0 _0869_
rlabel metal2 28672 20776 28672 20776 0 _0870_
rlabel metal2 4704 11368 4704 11368 0 _0871_
rlabel metal2 6104 10920 6104 10920 0 _0872_
rlabel metal3 4984 11368 4984 11368 0 _0873_
rlabel metal2 8848 12152 8848 12152 0 _0874_
rlabel metal3 13608 10808 13608 10808 0 _0875_
rlabel metal2 13944 11088 13944 11088 0 _0876_
rlabel metal3 11536 11368 11536 11368 0 _0877_
rlabel metal3 7056 10024 7056 10024 0 _0878_
rlabel metal2 7448 10360 7448 10360 0 _0879_
rlabel metal3 8288 10696 8288 10696 0 _0880_
rlabel metal3 9576 12152 9576 12152 0 _0881_
rlabel metal3 20328 10864 20328 10864 0 _0882_
rlabel metal2 26040 11088 26040 11088 0 _0883_
rlabel metal2 26824 11816 26824 11816 0 _0884_
rlabel metal2 14000 8344 14000 8344 0 _0885_
rlabel metal3 14056 7672 14056 7672 0 _0886_
rlabel metal2 18536 7728 18536 7728 0 _0887_
rlabel metal2 17528 8960 17528 8960 0 _0888_
rlabel metal2 18536 10136 18536 10136 0 _0889_
rlabel metal2 18312 8904 18312 8904 0 _0890_
rlabel metal3 20608 5880 20608 5880 0 _0891_
rlabel metal2 48832 4312 48832 4312 0 _0892_
rlabel metal2 51240 3472 51240 3472 0 _0893_
rlabel metal2 19544 6664 19544 6664 0 _0894_
rlabel metal2 18928 8232 18928 8232 0 _0895_
rlabel metal3 19656 8120 19656 8120 0 _0896_
rlabel metal2 19208 8176 19208 8176 0 _0897_
rlabel metal2 35168 27720 35168 27720 0 _0898_
rlabel metal2 37912 28168 37912 28168 0 _0899_
rlabel metal2 31864 26712 31864 26712 0 _0900_
rlabel metal3 34216 26152 34216 26152 0 _0901_
rlabel metal3 8400 14280 8400 14280 0 _0902_
rlabel metal2 9968 13496 9968 13496 0 _0903_
rlabel metal2 33824 26152 33824 26152 0 _0904_
rlabel metal2 67816 21168 67816 21168 0 _0905_
rlabel metal2 53480 29904 53480 29904 0 _0906_
rlabel metal2 39816 25928 39816 25928 0 _0907_
rlabel metal3 39480 27272 39480 27272 0 _0908_
rlabel metal2 39144 26768 39144 26768 0 _0909_
rlabel metal2 34328 25760 34328 25760 0 _0910_
rlabel metal2 27048 23576 27048 23576 0 _0911_
rlabel metal2 26600 21952 26600 21952 0 _0912_
rlabel metal3 26656 24024 26656 24024 0 _0913_
rlabel metal3 28672 23688 28672 23688 0 _0914_
rlabel metal2 27440 21448 27440 21448 0 _0915_
rlabel metal3 29344 20216 29344 20216 0 _0916_
rlabel metal3 30016 23800 30016 23800 0 _0917_
rlabel metal2 30968 25088 30968 25088 0 _0918_
rlabel metal2 34944 26152 34944 26152 0 _0919_
rlabel metal2 35560 26376 35560 26376 0 _0920_
rlabel metal2 37128 28280 37128 28280 0 _0921_
rlabel metal2 37912 30128 37912 30128 0 _0922_
rlabel metal2 41832 32144 41832 32144 0 _0923_
rlabel metal2 42560 34328 42560 34328 0 _0924_
rlabel metal2 38136 32032 38136 32032 0 _0925_
rlabel metal2 37688 32480 37688 32480 0 _0926_
rlabel metal3 40488 33880 40488 33880 0 _0927_
rlabel metal2 48216 35168 48216 35168 0 _0928_
rlabel metal2 44184 36008 44184 36008 0 _0929_
rlabel metal3 44968 33320 44968 33320 0 _0930_
rlabel metal3 40936 30968 40936 30968 0 _0931_
rlabel metal2 41216 30968 41216 30968 0 _0932_
rlabel metal3 42840 31080 42840 31080 0 _0933_
rlabel metal3 35448 26488 35448 26488 0 _0934_
rlabel metal2 39928 27440 39928 27440 0 _0935_
rlabel metal3 41216 29400 41216 29400 0 _0936_
rlabel metal3 37184 28616 37184 28616 0 _0937_
rlabel metal2 38024 28896 38024 28896 0 _0938_
rlabel metal2 30632 24360 30632 24360 0 _0939_
rlabel metal2 32872 25032 32872 25032 0 _0940_
rlabel metal3 33208 24696 33208 24696 0 _0941_
rlabel metal2 8680 10360 8680 10360 0 _0942_
rlabel metal3 33152 23688 33152 23688 0 _0943_
rlabel metal2 68936 15456 68936 15456 0 _0944_
rlabel metal3 39928 23128 39928 23128 0 _0945_
rlabel metal2 40936 22736 40936 22736 0 _0946_
rlabel metal2 40824 22680 40824 22680 0 _0947_
rlabel metal2 40152 22960 40152 22960 0 _0948_
rlabel metal2 33880 22736 33880 22736 0 _0949_
rlabel metal2 30296 19376 30296 19376 0 _0950_
rlabel metal2 26040 21168 26040 21168 0 _0951_
rlabel metal2 32760 21112 32760 21112 0 _0952_
rlabel metal2 30352 19992 30352 19992 0 _0953_
rlabel metal2 31752 19376 31752 19376 0 _0954_
rlabel metal2 31976 22008 31976 22008 0 _0955_
rlabel metal2 34160 22344 34160 22344 0 _0956_
rlabel metal3 34328 23912 34328 23912 0 _0957_
rlabel metal3 34944 24696 34944 24696 0 _0958_
rlabel metal2 37128 24640 37128 24640 0 _0959_
rlabel metal3 28784 11368 28784 11368 0 _0960_
rlabel metal2 30016 11256 30016 11256 0 _0961_
rlabel metal2 35560 12320 35560 12320 0 _0962_
rlabel metal2 8400 7448 8400 7448 0 _0963_
rlabel metal3 6440 9912 6440 9912 0 _0964_
rlabel metal2 10472 10192 10472 10192 0 _0965_
rlabel metal2 16296 5824 16296 5824 0 _0966_
rlabel metal2 13832 8120 13832 8120 0 _0967_
rlabel metal3 12824 9128 12824 9128 0 _0968_
rlabel metal3 4928 9016 4928 9016 0 _0969_
rlabel metal3 9016 6664 9016 6664 0 _0970_
rlabel metal3 6272 8232 6272 8232 0 _0971_
rlabel metal2 10472 8736 10472 8736 0 _0972_
rlabel metal2 11368 9520 11368 9520 0 _0973_
rlabel metal2 25032 9520 25032 9520 0 _0974_
rlabel metal2 19544 8624 19544 8624 0 _0975_
rlabel metal2 23576 8736 23576 8736 0 _0976_
rlabel metal2 12936 6720 12936 6720 0 _0977_
rlabel metal2 15288 4200 15288 4200 0 _0978_
rlabel metal2 22008 5824 22008 5824 0 _0979_
rlabel metal2 23912 5488 23912 5488 0 _0980_
rlabel metal2 23240 6048 23240 6048 0 _0981_
rlabel metal2 22568 5432 22568 5432 0 _0982_
rlabel metal2 24584 4816 24584 4816 0 _0983_
rlabel metal2 51352 5712 51352 5712 0 _0984_
rlabel metal2 40376 3640 40376 3640 0 _0985_
rlabel metal3 23744 5208 23744 5208 0 _0986_
rlabel metal2 22232 5600 22232 5600 0 _0987_
rlabel metal2 23800 8176 23800 8176 0 _0988_
rlabel metal3 25368 9128 25368 9128 0 _0989_
rlabel metal2 26824 10136 26824 10136 0 _0990_
rlabel metal2 38192 23016 38192 23016 0 _0991_
rlabel metal2 38584 28728 38584 28728 0 _0992_
rlabel metal2 43848 31360 43848 31360 0 _0993_
rlabel metal2 43960 32648 43960 32648 0 _0994_
rlabel metal2 51016 33208 51016 33208 0 _0995_
rlabel metal3 49224 34776 49224 34776 0 _0996_
rlabel metal2 43176 34048 43176 34048 0 _0997_
rlabel metal2 50008 34776 50008 34776 0 _0998_
rlabel metal2 52024 35112 52024 35112 0 _0999_
rlabel metal3 52472 35784 52472 35784 0 _1000_
rlabel metal2 51576 33320 51576 33320 0 _1001_
rlabel metal3 52360 34104 52360 34104 0 _1002_
rlabel metal2 51296 34216 51296 34216 0 _1003_
rlabel metal2 45416 30800 45416 30800 0 _1004_
rlabel metal2 46424 32088 46424 32088 0 _1005_
rlabel metal2 39928 29400 39928 29400 0 _1006_
rlabel metal2 40656 28840 40656 28840 0 _1007_
rlabel metal2 44632 29792 44632 29792 0 _1008_
rlabel metal2 69608 20832 69608 20832 0 _1009_
rlabel metal2 43848 25760 43848 25760 0 _1010_
rlabel metal3 35280 23688 35280 23688 0 _1011_
rlabel metal2 35448 24192 35448 24192 0 _1012_
rlabel metal2 35784 24080 35784 24080 0 _1013_
rlabel metal2 41720 23520 41720 23520 0 _1014_
rlabel metal2 40768 24136 40768 24136 0 _1015_
rlabel metal3 41944 23800 41944 23800 0 _1016_
rlabel metal2 43512 25144 43512 25144 0 _1017_
rlabel metal2 4536 22400 4536 22400 0 _1018_
rlabel metal3 40936 26376 40936 26376 0 _1019_
rlabel metal3 37352 23688 37352 23688 0 _1020_
rlabel metal2 38920 24248 38920 24248 0 _1021_
rlabel metal2 32368 21560 32368 21560 0 _1022_
rlabel metal2 33040 21784 33040 21784 0 _1023_
rlabel metal3 34888 21672 34888 21672 0 _1024_
rlabel metal2 10976 10808 10976 10808 0 _1025_
rlabel metal2 11928 8792 11928 8792 0 _1026_
rlabel metal2 31248 17976 31248 17976 0 _1027_
rlabel metal2 40376 20440 40376 20440 0 _1028_
rlabel metal2 9912 24472 9912 24472 0 _1029_
rlabel metal3 41552 18424 41552 18424 0 _1030_
rlabel metal2 42168 20328 42168 20328 0 _1031_
rlabel metal3 40600 20888 40600 20888 0 _1032_
rlabel metal2 41160 21000 41160 21000 0 _1033_
rlabel metal2 35672 18928 35672 18928 0 _1034_
rlabel metal2 29960 15624 29960 15624 0 _1035_
rlabel metal2 30800 19432 30800 19432 0 _1036_
rlabel metal2 30968 19544 30968 19544 0 _1037_
rlabel metal3 29120 18424 29120 18424 0 _1038_
rlabel metal2 31304 18424 31304 18424 0 _1039_
rlabel metal3 16632 18648 16632 18648 0 _1040_
rlabel metal2 33880 18928 33880 18928 0 _1041_
rlabel metal2 35952 18648 35952 18648 0 _1042_
rlabel metal2 35280 19320 35280 19320 0 _1043_
rlabel metal2 36120 21224 36120 21224 0 _1044_
rlabel metal3 37184 21560 37184 21560 0 _1045_
rlabel metal3 24976 9240 24976 9240 0 _1046_
rlabel metal2 29736 9408 29736 9408 0 _1047_
rlabel metal3 20468 6440 20468 6440 0 _1048_
rlabel metal2 4200 7504 4200 7504 0 _1049_
rlabel metal2 18872 5208 18872 5208 0 _1050_
rlabel metal2 18088 15232 18088 15232 0 _1051_
rlabel metal2 13776 5320 13776 5320 0 _1052_
rlabel metal2 6104 6384 6104 6384 0 _1053_
rlabel metal3 7672 5320 7672 5320 0 _1054_
rlabel metal2 8680 6160 8680 6160 0 _1055_
rlabel metal2 4424 6272 4424 6272 0 _1056_
rlabel metal3 5152 7448 5152 7448 0 _1057_
rlabel metal2 21672 7784 21672 7784 0 _1058_
rlabel metal2 21952 4088 21952 4088 0 _1059_
rlabel metal2 22792 7504 22792 7504 0 _1060_
rlabel metal3 26320 1624 26320 1624 0 _1061_
rlabel metal3 21112 26936 21112 26936 0 _1062_
rlabel metal2 16296 4648 16296 4648 0 _1063_
rlabel metal2 20104 4704 20104 4704 0 _1064_
rlabel metal2 45416 7280 45416 7280 0 _1065_
rlabel metal2 44184 4816 44184 4816 0 _1066_
rlabel metal3 26712 4312 26712 4312 0 _1067_
rlabel metal2 21336 4312 21336 4312 0 _1068_
rlabel metal2 39760 5320 39760 5320 0 _1069_
rlabel metal2 49784 6104 49784 6104 0 _1070_
rlabel metal2 29176 4704 29176 4704 0 _1071_
rlabel metal3 24976 3192 24976 3192 0 _1072_
rlabel metal2 18872 28224 18872 28224 0 _1073_
rlabel metal2 20104 3864 20104 3864 0 _1074_
rlabel metal3 21392 7336 21392 7336 0 _1075_
rlabel metal3 23072 8232 23072 8232 0 _1076_
rlabel metal2 29624 9016 29624 9016 0 _1077_
rlabel metal3 36904 22120 36904 22120 0 _1078_
rlabel metal2 38584 23128 38584 23128 0 _1079_
rlabel metal2 39480 25480 39480 25480 0 _1080_
rlabel metal2 44408 28896 44408 28896 0 _1081_
rlabel metal2 47656 32144 47656 32144 0 _1082_
rlabel metal2 50792 33040 50792 33040 0 _1083_
rlabel metal2 46872 4200 46872 4200 0 _1084_
rlabel metal2 51408 33992 51408 33992 0 _1085_
rlabel metal2 42056 24640 42056 24640 0 _1086_
rlabel metal3 70112 20776 70112 20776 0 _1087_
rlabel metal2 44632 25144 44632 25144 0 _1088_
rlabel metal2 45864 26180 45864 26180 0 _1089_
rlabel metal2 39200 23912 39200 23912 0 _1090_
rlabel metal3 43288 26264 43288 26264 0 _1091_
rlabel metal3 35840 21000 35840 21000 0 _1092_
rlabel metal2 36680 21896 36680 21896 0 _1093_
rlabel metal3 16856 18536 16856 18536 0 _1094_
rlabel metal2 42000 19880 42000 19880 0 _1095_
rlabel metal3 44128 22344 44128 22344 0 _1096_
rlabel metal3 44912 23128 44912 23128 0 _1097_
rlabel metal2 36400 22120 36400 22120 0 _1098_
rlabel metal2 44296 22008 44296 22008 0 _1099_
rlabel metal2 34496 18536 34496 18536 0 _1100_
rlabel metal2 35056 18424 35056 18424 0 _1101_
rlabel metal3 33768 13720 33768 13720 0 _1102_
rlabel metal2 5936 7672 5936 7672 0 _1103_
rlabel metal2 4760 7056 4760 7056 0 _1104_
rlabel metal3 22008 21672 22008 21672 0 _1105_
rlabel metal2 5544 7448 5544 7448 0 _1106_
rlabel metal2 40600 18704 40600 18704 0 _1107_
rlabel metal3 43064 18312 43064 18312 0 _1108_
rlabel metal2 42392 18648 42392 18648 0 _1109_
rlabel metal2 35672 16856 35672 16856 0 _1110_
rlabel metal2 31192 17304 31192 17304 0 _1111_
rlabel metal2 32592 17640 32592 17640 0 _1112_
rlabel metal2 31864 16184 31864 16184 0 _1113_
rlabel metal2 31976 16576 31976 16576 0 _1114_
rlabel metal2 31864 16912 31864 16912 0 _1115_
rlabel metal2 21504 27720 21504 27720 0 _1116_
rlabel metal2 32144 16184 32144 16184 0 _1117_
rlabel metal3 33096 15960 33096 15960 0 _1118_
rlabel metal2 33992 13664 33992 13664 0 _1119_
rlabel metal2 34216 12488 34216 12488 0 _1120_
rlabel metal3 22960 7672 22960 7672 0 _1121_
rlabel metal2 22568 7952 22568 7952 0 _1122_
rlabel metal2 56616 2296 56616 2296 0 _1123_
rlabel metal3 9520 5768 9520 5768 0 _1124_
rlabel via2 10360 5096 10360 5096 0 _1125_
rlabel metal3 14000 3416 14000 3416 0 _1126_
rlabel metal3 26712 27048 26712 27048 0 _1127_
rlabel metal2 15512 4256 15512 4256 0 _1128_
rlabel metal2 15288 3304 15288 3304 0 _1129_
rlabel metal2 27608 6272 27608 6272 0 _1130_
rlabel metal3 29456 8120 29456 8120 0 _1131_
rlabel metal2 26712 5600 26712 5600 0 _1132_
rlabel metal2 10584 4816 10584 4816 0 _1133_
rlabel metal3 20440 2408 20440 2408 0 _1134_
rlabel metal2 21112 4816 21112 4816 0 _1135_
rlabel metal2 31248 4536 31248 4536 0 _1136_
rlabel metal2 54376 3248 54376 3248 0 _1137_
rlabel metal2 22680 27440 22680 27440 0 _1138_
rlabel metal3 37296 5992 37296 5992 0 _1139_
rlabel metal2 36792 4648 36792 4648 0 _1140_
rlabel metal2 47656 5208 47656 5208 0 _1141_
rlabel metal2 41888 4536 41888 4536 0 _1142_
rlabel metal2 39480 4592 39480 4592 0 _1143_
rlabel metal2 47544 3696 47544 3696 0 _1144_
rlabel metal3 49952 5096 49952 5096 0 _1145_
rlabel metal2 49224 6160 49224 6160 0 _1146_
rlabel metal2 39256 4536 39256 4536 0 _1147_
rlabel metal3 35336 4200 35336 4200 0 _1148_
rlabel metal2 18648 29064 18648 29064 0 _1149_
rlabel metal3 33208 4312 33208 4312 0 _1150_
rlabel metal2 33208 9072 33208 9072 0 _1151_
rlabel metal2 34440 11704 34440 11704 0 _1152_
rlabel metal2 43848 20832 43848 20832 0 _1153_
rlabel metal2 44520 23240 44520 23240 0 _1154_
rlabel metal2 44744 25032 44744 25032 0 _1155_
rlabel metal3 45976 27832 45976 27832 0 _1156_
rlabel metal2 46648 28672 46648 28672 0 _1157_
rlabel metal3 47488 30072 47488 30072 0 _1158_
rlabel metal2 44744 30240 44744 30240 0 _1159_
rlabel metal2 45864 5376 45864 5376 0 _1160_
rlabel metal2 46368 28728 46368 28728 0 _1161_
rlabel metal2 51352 29344 51352 29344 0 _1162_
rlabel metal2 51464 29008 51464 29008 0 _1163_
rlabel metal3 50792 29624 50792 29624 0 _1164_
rlabel metal2 50120 32984 50120 32984 0 _1165_
rlabel metal2 46592 31192 46592 31192 0 _1166_
rlabel metal3 47096 31640 47096 31640 0 _1167_
rlabel metal2 46536 32200 46536 32200 0 _1168_
rlabel metal2 49784 31416 49784 31416 0 _1169_
rlabel metal2 49896 34384 49896 34384 0 _1170_
rlabel metal2 17752 27496 17752 27496 0 _1171_
rlabel metal3 49672 31752 49672 31752 0 _1172_
rlabel metal2 50568 30912 50568 30912 0 _1173_
rlabel metal3 49280 30296 49280 30296 0 _1174_
rlabel metal3 45584 27048 45584 27048 0 _1175_
rlabel metal2 48776 27496 48776 27496 0 _1176_
rlabel metal2 48104 24080 48104 24080 0 _1177_
rlabel metal2 44576 21784 44576 21784 0 _1178_
rlabel metal3 46704 23240 46704 23240 0 _1179_
rlabel metal3 35840 13720 35840 13720 0 _1180_
rlabel metal2 27384 27776 27384 27776 0 _1181_
rlabel metal2 34776 14000 34776 14000 0 _1182_
rlabel metal2 34776 18368 34776 18368 0 _1183_
rlabel metal2 43848 18648 43848 18648 0 _1184_
rlabel metal3 43176 19320 43176 19320 0 _1185_
rlabel metal3 45192 19992 45192 19992 0 _1186_
rlabel metal2 48328 21168 48328 21168 0 _1187_
rlabel metal3 45640 20104 45640 20104 0 _1188_
rlabel metal2 45416 20496 45416 20496 0 _1189_
rlabel metal2 33544 10584 33544 10584 0 _1190_
rlabel metal2 41944 12096 41944 12096 0 _1191_
rlabel metal2 27048 27440 27048 27440 0 _1192_
rlabel metal2 34216 15848 34216 15848 0 _1193_
rlabel metal2 34776 15568 34776 15568 0 _1194_
rlabel metal2 34328 15624 34328 15624 0 _1195_
rlabel metal3 10864 3528 10864 3528 0 _1196_
rlabel metal2 11872 3416 11872 3416 0 _1197_
rlabel metal2 11816 2072 11816 2072 0 _1198_
rlabel metal3 51520 31528 51520 31528 0 _1199_
rlabel metal3 39144 17640 39144 17640 0 _1200_
rlabel metal3 44464 16968 44464 16968 0 _1201_
rlabel metal3 40712 17752 40712 17752 0 _1202_
rlabel metal2 20216 28504 20216 28504 0 _1203_
rlabel metal2 39704 16464 39704 16464 0 _1204_
rlabel metal2 31752 15680 31752 15680 0 _1205_
rlabel metal2 37632 15848 37632 15848 0 _1206_
rlabel metal3 37352 17640 37352 17640 0 _1207_
rlabel metal2 35112 16408 35112 16408 0 _1208_
rlabel metal3 36848 16856 36848 16856 0 _1209_
rlabel metal2 38584 16856 38584 16856 0 _1210_
rlabel metal2 39144 15624 39144 15624 0 _1211_
rlabel metal2 38024 14224 38024 14224 0 _1212_
rlabel metal2 39144 14000 39144 14000 0 _1213_
rlabel metal2 21336 29120 21336 29120 0 _1214_
rlabel metal3 40152 13720 40152 13720 0 _1215_
rlabel metal3 33880 3752 33880 3752 0 _1216_
rlabel metal2 39144 10696 39144 10696 0 _1217_
rlabel metal2 28560 7672 28560 7672 0 _1218_
rlabel metal2 27776 6776 27776 6776 0 _1219_
rlabel metal3 29624 6552 29624 6552 0 _1220_
rlabel metal3 35672 6552 35672 6552 0 _1221_
rlabel metal2 35392 6104 35392 6104 0 _1222_
rlabel metal3 33712 6664 33712 6664 0 _1223_
rlabel metal2 32312 9016 32312 9016 0 _1224_
rlabel metal2 24304 25368 24304 25368 0 _1225_
rlabel metal2 42728 9128 42728 9128 0 _1226_
rlabel metal3 30128 8232 30128 8232 0 _1227_
rlabel metal2 31528 7112 31528 7112 0 _1228_
rlabel metal2 32536 6384 32536 6384 0 _1229_
rlabel metal3 39144 5880 39144 5880 0 _1230_
rlabel metal2 38192 4536 38192 4536 0 _1231_
rlabel metal2 40376 5936 40376 5936 0 _1232_
rlabel metal3 35784 7336 35784 7336 0 _1233_
rlabel metal2 42056 8344 42056 8344 0 _1234_
rlabel metal2 44520 7392 44520 7392 0 _1235_
rlabel metal2 51352 3696 51352 3696 0 _1236_
rlabel metal2 44688 6440 44688 6440 0 _1237_
rlabel metal2 45192 3976 45192 3976 0 _1238_
rlabel metal3 45304 4984 45304 4984 0 _1239_
rlabel metal2 48496 4536 48496 4536 0 _1240_
rlabel metal2 51688 6160 51688 6160 0 _1241_
rlabel metal2 45752 5096 45752 5096 0 _1242_
rlabel metal2 44240 7448 44240 7448 0 _1243_
rlabel metal3 40544 6664 40544 6664 0 _1244_
rlabel metal2 39928 7168 39928 7168 0 _1245_
rlabel metal3 21896 29288 21896 29288 0 _1246_
rlabel metal2 39200 5992 39200 5992 0 _1247_
rlabel metal2 39928 12880 39928 12880 0 _1248_
rlabel metal3 41664 12936 41664 12936 0 _1249_
rlabel metal2 45416 17864 45416 17864 0 _1250_
rlabel metal3 47152 21560 47152 21560 0 _1251_
rlabel metal2 45976 27440 45976 27440 0 _1252_
rlabel metal2 52920 27776 52920 27776 0 _1253_
rlabel metal2 50456 28896 50456 28896 0 _1254_
rlabel metal3 48272 29400 48272 29400 0 _1255_
rlabel metal3 23408 29400 23408 29400 0 _1256_
rlabel metal2 44520 18536 44520 18536 0 _1257_
rlabel metal2 48664 19992 48664 19992 0 _1258_
rlabel metal2 37744 13944 37744 13944 0 _1259_
rlabel metal3 40152 14392 40152 14392 0 _1260_
rlabel metal2 39816 14840 39816 14840 0 _1261_
rlabel metal2 46984 18032 46984 18032 0 _1262_
rlabel metal2 40040 11872 40040 11872 0 _1263_
rlabel metal2 45976 14336 45976 14336 0 _1264_
rlabel metal2 42504 14504 42504 14504 0 _1265_
rlabel metal2 31192 7056 31192 7056 0 _1266_
rlabel metal2 32032 7448 32032 7448 0 _1267_
rlabel metal2 41608 13888 41608 13888 0 _1268_
rlabel metal2 36680 17696 36680 17696 0 _1269_
rlabel metal2 37912 16688 37912 16688 0 _1270_
rlabel metal2 51688 17136 51688 17136 0 _1271_
rlabel metal2 50568 17248 50568 17248 0 _1272_
rlabel metal2 51576 17304 51576 17304 0 _1273_
rlabel metal3 52304 16744 52304 16744 0 _1274_
rlabel metal3 47096 16800 47096 16800 0 _1275_
rlabel metal2 44184 16072 44184 16072 0 _1276_
rlabel metal2 20888 30520 20888 30520 0 _1277_
rlabel metal2 44968 13328 44968 13328 0 _1278_
rlabel metal2 41048 7056 41048 7056 0 _1279_
rlabel metal2 40152 7672 40152 7672 0 _1280_
rlabel metal2 31472 9240 31472 9240 0 _1281_
rlabel metal2 40600 10920 40600 10920 0 _1282_
rlabel metal2 41608 8232 41608 8232 0 _1283_
rlabel metal3 37296 8232 37296 8232 0 _1284_
rlabel metal2 38304 10584 38304 10584 0 _1285_
rlabel metal2 35896 10864 35896 10864 0 _1286_
rlabel metal3 56168 10808 56168 10808 0 _1287_
rlabel metal2 13832 17136 13832 17136 0 _1288_
rlabel metal3 33936 10584 33936 10584 0 _1289_
rlabel metal2 38584 10136 38584 10136 0 _1290_
rlabel metal2 40096 9800 40096 9800 0 _1291_
rlabel metal3 44576 10584 44576 10584 0 _1292_
rlabel metal2 45360 5096 45360 5096 0 _1293_
rlabel metal2 44408 8036 44408 8036 0 _1294_
rlabel metal3 41272 9016 41272 9016 0 _1295_
rlabel metal2 50680 7952 50680 7952 0 _1296_
rlabel metal3 46984 8120 46984 8120 0 _1297_
rlabel metal2 49784 5656 49784 5656 0 _1298_
rlabel metal2 13272 26376 13272 26376 0 _1299_
rlabel metal3 47152 5768 47152 5768 0 _1300_
rlabel metal2 48328 7504 48328 7504 0 _1301_
rlabel metal2 50120 7112 50120 7112 0 _1302_
rlabel metal2 53592 5880 53592 5880 0 _1303_
rlabel metal2 48440 7336 48440 7336 0 _1304_
rlabel metal3 47096 8232 47096 8232 0 _1305_
rlabel metal2 45808 8344 45808 8344 0 _1306_
rlabel metal2 45528 10192 45528 10192 0 _1307_
rlabel metal2 44184 11704 44184 11704 0 _1308_
rlabel metal2 44520 12768 44520 12768 0 _1309_
rlabel metal3 19376 30968 19376 30968 0 _1310_
rlabel metal2 46200 14224 46200 14224 0 _1311_
rlabel metal2 46760 14924 46760 14924 0 _1312_
rlabel metal2 48440 20160 48440 20160 0 _1313_
rlabel metal2 49896 21168 49896 21168 0 _1314_
rlabel metal2 48104 22736 48104 22736 0 _1315_
rlabel metal2 48104 22064 48104 22064 0 _1316_
rlabel metal2 52360 23800 52360 23800 0 _1317_
rlabel metal3 53648 25480 53648 25480 0 _1318_
rlabel metal2 48440 25032 48440 25032 0 _1319_
rlabel metal2 48832 26488 48832 26488 0 _1320_
rlabel metal2 17752 29008 17752 29008 0 _1321_
rlabel metal2 49560 27048 49560 27048 0 _1322_
rlabel metal3 47432 27048 47432 27048 0 _1323_
rlabel metal2 53704 27888 53704 27888 0 _1324_
rlabel metal2 53592 28000 53592 28000 0 _1325_
rlabel metal3 53536 27944 53536 27944 0 _1326_
rlabel metal2 54936 27440 54936 27440 0 _1327_
rlabel metal2 54600 27328 54600 27328 0 _1328_
rlabel metal2 53480 26040 53480 26040 0 _1329_
rlabel metal2 48552 20216 48552 20216 0 _1330_
rlabel metal2 19096 28280 19096 28280 0 _1331_
rlabel metal2 49168 21560 49168 21560 0 _1332_
rlabel metal2 50008 21952 50008 21952 0 _1333_
rlabel metal2 48216 18928 48216 18928 0 _1334_
rlabel metal3 46928 15736 46928 15736 0 _1335_
rlabel metal2 47936 19320 47936 19320 0 _1336_
rlabel metal2 43176 14560 43176 14560 0 _1337_
rlabel metal2 43848 14504 43848 14504 0 _1338_
rlabel metal2 48776 14280 48776 14280 0 _1339_
rlabel metal2 44296 12152 44296 12152 0 _1340_
rlabel metal2 48664 13720 48664 13720 0 _1341_
rlabel metal2 18984 29008 18984 29008 0 _1342_
rlabel metal2 46200 17080 46200 17080 0 _1343_
rlabel metal2 46200 15680 46200 15680 0 _1344_
rlabel metal2 46592 15960 46592 15960 0 _1345_
rlabel metal3 50512 14504 50512 14504 0 _1346_
rlabel metal2 39928 9968 39928 9968 0 _1347_
rlabel metal2 39200 9800 39200 9800 0 _1348_
rlabel metal2 52696 12600 52696 12600 0 _1349_
rlabel metal3 56672 15848 56672 15848 0 _1350_
rlabel metal3 50064 14616 50064 14616 0 _1351_
rlabel via2 54824 15960 54824 15960 0 _1352_
rlabel metal2 18424 26600 18424 26600 0 _1353_
rlabel metal2 54040 14784 54040 14784 0 _1354_
rlabel metal2 52808 17304 52808 17304 0 _1355_
rlabel metal2 54096 13720 54096 13720 0 _1356_
rlabel metal2 54376 13160 54376 13160 0 _1357_
rlabel metal2 54488 12600 54488 12600 0 _1358_
rlabel metal2 50904 12488 50904 12488 0 _1359_
rlabel metal2 44632 10304 44632 10304 0 _1360_
rlabel metal3 47040 12264 47040 12264 0 _1361_
rlabel metal2 43960 9520 43960 9520 0 _1362_
rlabel metal2 43176 10304 43176 10304 0 _1363_
rlabel metal2 17976 25816 17976 25816 0 _1364_
rlabel metal2 35784 10136 35784 10136 0 _1365_
rlabel metal2 51016 10752 51016 10752 0 _1366_
rlabel metal3 49112 9128 49112 9128 0 _1367_
rlabel metal2 41776 9016 41776 9016 0 _1368_
rlabel metal2 54264 10640 54264 10640 0 _1369_
rlabel metal3 57680 11368 57680 11368 0 _1370_
rlabel metal2 68992 8792 68992 8792 0 _1371_
rlabel metal3 57624 11480 57624 11480 0 _1372_
rlabel metal2 54376 10920 54376 10920 0 _1373_
rlabel metal2 53032 11032 53032 11032 0 _1374_
rlabel metal3 7728 21672 7728 21672 0 _1375_
rlabel metal3 50232 11368 50232 11368 0 _1376_
rlabel metal2 48104 7952 48104 7952 0 _1377_
rlabel metal2 48664 10248 48664 10248 0 _1378_
rlabel metal2 51240 9296 51240 9296 0 _1379_
rlabel metal2 49224 9128 49224 9128 0 _1380_
rlabel metal2 54824 8960 54824 8960 0 _1381_
rlabel metal2 51576 7728 51576 7728 0 _1382_
rlabel metal3 54656 30072 54656 30072 0 _1383_
rlabel metal3 51688 31640 51688 31640 0 _1384_
rlabel metal3 51912 6664 51912 6664 0 _1385_
rlabel metal2 37688 19656 37688 19656 0 _1386_
rlabel metal2 2744 2142 2744 2142 0 clk
rlabel metal3 10472 4312 10472 4312 0 dba[0]
rlabel metal2 32536 1526 32536 1526 0 dba[10]
rlabel metal2 34776 2184 34776 2184 0 dba[11]
rlabel metal3 36568 3528 36568 3528 0 dba[12]
rlabel metal2 39144 4032 39144 4032 0 dba[13]
rlabel metal2 41160 3416 41160 3416 0 dba[14]
rlabel metal2 43344 4424 43344 4424 0 dba[15]
rlabel metal2 13608 3640 13608 3640 0 dba[1]
rlabel metal2 15512 854 15512 854 0 dba[2]
rlabel metal2 17976 4592 17976 4592 0 dba[3]
rlabel metal3 18424 3528 18424 3528 0 dba[4]
rlabel metal3 21560 3528 21560 3528 0 dba[5]
rlabel metal2 24024 854 24024 854 0 dba[6]
rlabel metal3 24976 3416 24976 3416 0 dba[7]
rlabel metal3 28784 3528 28784 3528 0 dba[8]
rlabel metal2 30520 2184 30520 2184 0 dba[9]
rlabel metal3 46648 3416 46648 3416 0 dbb[0]
rlabel metal3 70504 4984 70504 4984 0 dbb[10]
rlabel metal2 70280 3528 70280 3528 0 dbb[11]
rlabel metal3 74592 3416 74592 3416 0 dbb[12]
rlabel metal2 73416 4368 73416 4368 0 dbb[13]
rlabel metal2 74424 2520 74424 2520 0 dbb[14]
rlabel metal2 76776 3696 76776 3696 0 dbb[15]
rlabel metal2 51016 3472 51016 3472 0 dbb[1]
rlabel metal3 51520 4424 51520 4424 0 dbb[2]
rlabel metal2 52752 3528 52752 3528 0 dbb[3]
rlabel metal2 53816 1806 53816 1806 0 dbb[4]
rlabel metal2 56056 4312 56056 4312 0 dbb[5]
rlabel metal3 62328 3416 62328 3416 0 dbb[6]
rlabel metal2 63000 3472 63000 3472 0 dbb[7]
rlabel metal3 62944 4424 62944 4424 0 dbb[8]
rlabel metal2 64792 4760 64792 4760 0 dbb[9]
rlabel metal3 9744 3416 9744 3416 0 done
rlabel metal3 7504 3416 7504 3416 0 enable
rlabel metal3 2408 21784 2408 21784 0 net1
rlabel metal3 7728 20776 7728 20776 0 net10
rlabel metal2 27608 18704 27608 18704 0 net11
rlabel metal2 2576 12712 2576 12712 0 net12
rlabel metal2 29176 17360 29176 17360 0 net13
rlabel metal2 26712 3332 26712 3332 0 net14
rlabel metal3 29008 3304 29008 3304 0 net15
rlabel metal2 68488 7952 68488 7952 0 net16
rlabel metal2 47376 3640 47376 3640 0 net17
rlabel metal3 68656 6104 68656 6104 0 net18
rlabel metal2 68040 7616 68040 7616 0 net19
rlabel metal3 54432 4984 54432 4984 0 net2
rlabel metal2 68936 6216 68936 6216 0 net20
rlabel metal2 73192 4592 73192 4592 0 net21
rlabel metal2 74088 5376 74088 5376 0 net22
rlabel metal2 76328 3864 76328 3864 0 net23
rlabel metal2 46312 3304 46312 3304 0 net24
rlabel metal2 44408 5768 44408 5768 0 net25
rlabel metal2 48328 6272 48328 6272 0 net26
rlabel metal2 46536 5992 46536 5992 0 net27
rlabel metal2 50120 6160 50120 6160 0 net28
rlabel metal2 57736 4648 57736 4648 0 net29
rlabel metal2 69328 5208 69328 5208 0 net3
rlabel metal3 60088 3304 60088 3304 0 net30
rlabel metal2 62552 5488 62552 5488 0 net31
rlabel metal2 43960 4480 43960 4480 0 net32
rlabel metal3 5880 3472 5880 3472 0 net33
rlabel metal3 27384 25424 27384 25424 0 net34
rlabel metal2 27832 36512 27832 36512 0 net35
rlabel metal2 30520 36400 30520 36400 0 net36
rlabel metal2 51240 34552 51240 34552 0 net37
rlabel metal2 74200 36064 74200 36064 0 net38
rlabel metal2 53144 35952 53144 35952 0 net39
rlabel metal2 70280 6328 70280 6328 0 net4
rlabel metal2 52192 34776 52192 34776 0 net40
rlabel metal2 1624 17808 1624 17808 0 net41
rlabel metal2 1512 17416 1512 17416 0 net42
rlabel metal3 2072 7560 2072 7560 0 net43
rlabel metal2 2352 7672 2352 7672 0 net44
rlabel metal2 23800 27496 23800 27496 0 net45
rlabel metal3 2576 18536 2576 18536 0 net46
rlabel metal2 2464 26040 2464 26040 0 net47
rlabel metal2 2240 17640 2240 17640 0 net48
rlabel metal2 3976 19264 3976 19264 0 net49
rlabel metal2 50232 5152 50232 5152 0 net5
rlabel metal2 3192 30016 3192 30016 0 net50
rlabel metal3 4704 31640 4704 31640 0 net51
rlabel metal2 3696 32760 3696 32760 0 net52
rlabel metal2 3640 28784 3640 28784 0 net53
rlabel metal2 3192 33376 3192 33376 0 net54
rlabel metal3 5768 35000 5768 35000 0 net55
rlabel metal2 24024 29456 24024 29456 0 net56
rlabel metal2 4872 35280 4872 35280 0 net57
rlabel metal2 5320 36120 5320 36120 0 net58
rlabel metal3 75600 30968 75600 30968 0 net59
rlabel metal2 50904 3976 50904 3976 0 net6
rlabel metal3 21000 32984 21000 32984 0 net60
rlabel metal2 73584 34328 73584 34328 0 net61
rlabel metal2 77112 35784 77112 35784 0 net62
rlabel metal2 20440 35728 20440 35728 0 net63
rlabel metal2 24920 36848 24920 36848 0 net64
rlabel metal3 29904 34776 29904 34776 0 net65
rlabel metal3 7336 3640 7336 3640 0 net66
rlabel metal3 76608 3528 76608 3528 0 net67
rlabel metal2 78120 27664 78120 27664 0 net68
rlabel metal2 75264 29400 75264 29400 0 net69
rlabel metal2 54544 3528 54544 3528 0 net7
rlabel metal2 76216 32424 76216 32424 0 net70
rlabel metal2 74480 35784 74480 35784 0 net71
rlabel metal3 73920 36232 73920 36232 0 net72
rlabel metal3 74704 35784 74704 35784 0 net73
rlabel metal2 76496 4312 76496 4312 0 net74
rlabel metal2 76104 6720 76104 6720 0 net75
rlabel metal2 76384 28280 76384 28280 0 net76
rlabel metal3 77896 31752 77896 31752 0 net77
rlabel metal2 74816 14616 74816 14616 0 net78
rlabel metal3 77840 34216 77840 34216 0 net79
rlabel metal2 5656 20496 5656 20496 0 net8
rlabel metal2 77280 19320 77280 19320 0 net80
rlabel metal2 73696 34664 73696 34664 0 net81
rlabel metal2 77504 27048 77504 27048 0 net82
rlabel metal2 2968 4816 2968 4816 0 net83
rlabel metal2 2744 26264 2744 26264 0 net84
rlabel metal2 2856 28952 2856 28952 0 net85
rlabel metal2 2912 33096 2912 33096 0 net86
rlabel metal2 3080 34384 3080 34384 0 net87
rlabel metal2 3080 35728 3080 35728 0 net88
rlabel metal2 3080 35112 3080 35112 0 net89
rlabel metal3 2912 19992 2912 19992 0 net9
rlabel metal2 3080 4592 3080 4592 0 net90
rlabel metal2 3080 7112 3080 7112 0 net91
rlabel metal2 2800 9576 2800 9576 0 net92
rlabel metal2 2856 17080 2856 17080 0 net93
rlabel metal2 2856 14952 2856 14952 0 net94
rlabel metal2 2072 17136 2072 17136 0 net95
rlabel metal3 3360 19096 3360 19096 0 net96
rlabel metal2 3080 21056 3080 21056 0 net97
rlabel metal2 2744 29288 2744 29288 0 net98
rlabel metal2 74872 2576 74872 2576 0 yA[0]
rlabel metal3 77378 26152 77378 26152 0 yA[10]
rlabel metal2 76104 28952 76104 28952 0 yA[11]
rlabel metal2 75544 31472 75544 31472 0 yA[12]
rlabel metal2 76104 33824 76104 33824 0 yA[13]
rlabel metal2 76104 35840 76104 35840 0 yA[14]
rlabel metal2 77896 37128 77896 37128 0 yA[15]
rlabel metal2 75544 4088 75544 4088 0 yA[1]
rlabel metal2 75096 6496 75096 6496 0 yA[2]
rlabel metal3 77378 8904 77378 8904 0 yA[3]
rlabel metal2 75544 11760 75544 11760 0 yA[4]
rlabel metal2 76104 14112 76104 14112 0 yA[5]
rlabel metal3 76104 16800 76104 16800 0 yA[6]
rlabel metal2 75544 19152 75544 19152 0 yA[7]
rlabel metal2 76104 21336 76104 21336 0 yA[8]
rlabel metal2 75544 23856 75544 23856 0 yA[9]
rlabel metal3 1302 1512 1302 1512 0 yB[0]
rlabel metal3 1358 26152 1358 26152 0 yB[10]
rlabel metal3 1358 28616 1358 28616 0 yB[11]
rlabel metal3 1358 31080 1358 31080 0 yB[12]
rlabel metal3 1358 33544 1358 33544 0 yB[13]
rlabel metal3 1358 36008 1358 36008 0 yB[14]
rlabel metal3 1470 38472 1470 38472 0 yB[15]
rlabel metal3 1358 3976 1358 3976 0 yB[1]
rlabel metal3 1358 6440 1358 6440 0 yB[2]
rlabel metal3 1358 8904 1358 8904 0 yB[3]
rlabel metal3 1358 11368 1358 11368 0 yB[4]
rlabel metal3 1358 13832 1358 13832 0 yB[5]
rlabel metal3 1638 16296 1638 16296 0 yB[6]
rlabel metal3 1358 18760 1358 18760 0 yB[7]
rlabel metal3 1358 21224 1358 21224 0 yB[8]
rlabel metal3 1358 23688 1358 23688 0 yB[9]
<< properties >>
string FIXED_BBOX 0 0 80000 40000
<< end >>
