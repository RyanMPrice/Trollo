// This is the unpowered netlist.
module BinMultiplier (clk,
    done,
    enable,
    rst,
    Y,
    dba,
    dbb,
    yA,
    yB);
 input clk;
 output done;
 input enable;
 input rst;
 output [31:0] Y;
 input [15:0] dba;
 input [15:0] dbb;
 output [15:0] yA;
 output [15:0] yB;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;

 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1387_ (.I(net9),
    .Z(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1388_ (.I(_1018_),
    .Z(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1389_ (.I(net17),
    .Z(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1390_ (.I(_1040_),
    .Z(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1391_ (.I(_1051_),
    .Z(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1392_ (.A1(_1029_),
    .A2(_1062_),
    .ZN(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1393_ (.I(net24),
    .Z(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1394_ (.I(_1084_),
    .Z(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1395_ (.I(_1094_),
    .Z(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1396_ (.I(_1105_),
    .Z(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1397_ (.I(net8),
    .Z(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1398_ (.I(_1127_),
    .Z(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1399_ (.A1(_1116_),
    .A2(_1138_),
    .ZN(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1400_ (.I(net25),
    .Z(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1401_ (.I(_1160_),
    .Z(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1402_ (.I(net1),
    .Z(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1403_ (.I(_1181_),
    .Z(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1404_ (.A1(_1171_),
    .A2(_1192_),
    .Z(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _1405_ (.A1(_1073_),
    .A2(_1149_),
    .A3(_1203_),
    .ZN(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1406_ (.A1(_1062_),
    .A2(_1192_),
    .Z(_1225_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1407_ (.I(_1225_),
    .Z(net34));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1408_ (.A1(_1116_),
    .A2(_1138_),
    .A3(net34),
    .ZN(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1409_ (.A1(_1214_),
    .A2(_1246_),
    .Z(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1410_ (.I(_1256_),
    .Z(net56));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1411_ (.A1(_1214_),
    .A2(_1246_),
    .ZN(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1412_ (.I(net26),
    .Z(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1413_ (.I(_1288_),
    .Z(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1414_ (.A1(_1181_),
    .A2(_1299_),
    .ZN(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1415_ (.A1(_1073_),
    .A2(_1149_),
    .ZN(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1416_ (.A1(_1073_),
    .A2(_1149_),
    .ZN(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1417_ (.A1(_1321_),
    .A2(_1203_),
    .B(_1331_),
    .ZN(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1418_ (.A1(_1029_),
    .A2(_1116_),
    .ZN(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1419_ (.A1(_1138_),
    .A2(_1171_),
    .ZN(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1420_ (.I(net10),
    .Z(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1421_ (.I(_1375_),
    .Z(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1422_ (.A1(_1062_),
    .A2(_1386_),
    .ZN(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _1423_ (.A1(_1353_),
    .A2(_1364_),
    .A3(_0010_),
    .Z(_0020_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1424_ (.A1(_1342_),
    .A2(_0020_),
    .ZN(_0031_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1425_ (.A1(_1310_),
    .A2(_0031_),
    .Z(_0042_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1426_ (.A1(_1277_),
    .A2(_0042_),
    .Z(_0053_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1427_ (.I(_0053_),
    .Z(net59));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1428_ (.A1(_1277_),
    .A2(_0042_),
    .Z(_0074_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1429_ (.A1(_1138_),
    .A2(_1299_),
    .ZN(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1430_ (.I(net27),
    .Z(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1431_ (.I(_0095_),
    .Z(_0106_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1432_ (.A1(_1181_),
    .A2(_0106_),
    .ZN(_0117_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1433_ (.A1(_0085_),
    .A2(_0117_),
    .ZN(_0128_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1434_ (.A1(_1127_),
    .A2(_0106_),
    .ZN(_0139_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1435_ (.A1(_1310_),
    .A2(_0139_),
    .Z(_0150_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1436_ (.A1(_0128_),
    .A2(_0150_),
    .ZN(_0160_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1437_ (.A1(_1116_),
    .A2(_1386_),
    .ZN(_0171_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1438_ (.A1(_1029_),
    .A2(_1116_),
    .B1(_1386_),
    .B2(_1062_),
    .ZN(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _1439_ (.A1(_1073_),
    .A2(_0171_),
    .B1(_0182_),
    .B2(_1364_),
    .ZN(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1440_ (.A1(_1029_),
    .A2(_1171_),
    .ZN(_0204_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1441_ (.I(net11),
    .Z(_0214_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1442_ (.I(_0214_),
    .Z(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1443_ (.A1(_1051_),
    .A2(_0225_),
    .ZN(_0236_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _1444_ (.A1(_0171_),
    .A2(_0204_),
    .A3(_0236_),
    .ZN(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1445_ (.A1(_0193_),
    .A2(_0247_),
    .ZN(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1446_ (.A1(_0160_),
    .A2(_0258_),
    .Z(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1447_ (.A1(_1342_),
    .A2(_0020_),
    .Z(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1448_ (.A1(_1310_),
    .A2(_0031_),
    .B(_0279_),
    .ZN(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1449_ (.A1(_0268_),
    .A2(_0290_),
    .Z(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1450_ (.A1(_0074_),
    .A2(_0301_),
    .Z(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1451_ (.I(_0311_),
    .Z(net60));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1452_ (.A1(_0193_),
    .A2(_0247_),
    .ZN(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1453_ (.A1(_0193_),
    .A2(_0247_),
    .ZN(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1454_ (.A1(_0160_),
    .A2(_0332_),
    .B(_0343_),
    .ZN(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1455_ (.I(net28),
    .Z(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1456_ (.I(_0364_),
    .Z(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1457_ (.A1(net1),
    .A2(_0375_),
    .ZN(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1458_ (.A1(_1029_),
    .A2(_1299_),
    .ZN(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1459_ (.A1(_0139_),
    .A2(_0397_),
    .ZN(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1460_ (.A1(_0386_),
    .A2(_0407_),
    .ZN(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1461_ (.A1(_1105_),
    .A2(_0214_),
    .ZN(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1462_ (.A1(_1116_),
    .A2(_1386_),
    .B1(_0225_),
    .B2(_1062_),
    .ZN(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1463_ (.A1(_0010_),
    .A2(_0428_),
    .B1(_0439_),
    .B2(_0204_),
    .ZN(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1464_ (.A1(_1171_),
    .A2(_1375_),
    .ZN(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1465_ (.I(net12),
    .Z(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1466_ (.I(_0471_),
    .Z(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1467_ (.A1(_1051_),
    .A2(_0482_),
    .ZN(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _1468_ (.A1(_0428_),
    .A2(_0461_),
    .A3(_0492_),
    .ZN(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1469_ (.A1(_0450_),
    .A2(_0503_),
    .ZN(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1470_ (.A1(_0418_),
    .A2(_0512_),
    .Z(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1471_ (.A1(_0353_),
    .A2(_0515_),
    .ZN(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1472_ (.A1(_0150_),
    .A2(_0516_),
    .ZN(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1473_ (.A1(_0268_),
    .A2(_0290_),
    .ZN(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1474_ (.A1(_0074_),
    .A2(_0301_),
    .ZN(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1475_ (.A1(_0518_),
    .A2(_0519_),
    .ZN(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1476_ (.A1(_0517_),
    .A2(_0520_),
    .ZN(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1477_ (.I(_0521_),
    .Z(net61));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1478_ (.A1(_0518_),
    .A2(_0517_),
    .ZN(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1479_ (.A1(_1018_),
    .A2(_0106_),
    .ZN(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1480_ (.A1(_0085_),
    .A2(_0523_),
    .B1(_0407_),
    .B2(_0386_),
    .ZN(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1481_ (.I(net29),
    .Z(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1482_ (.I(_0525_),
    .Z(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1483_ (.A1(net1),
    .A2(_0526_),
    .ZN(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1484_ (.A1(_0524_),
    .A2(_0527_),
    .Z(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1485_ (.A1(_0450_),
    .A2(_0503_),
    .ZN(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1486_ (.A1(_0418_),
    .A2(_0512_),
    .B(_0529_),
    .ZN(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1487_ (.A1(_1094_),
    .A2(_0471_),
    .ZN(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1488_ (.A1(_1105_),
    .A2(_0225_),
    .B1(_0482_),
    .B2(_1051_),
    .ZN(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1489_ (.A1(_0236_),
    .A2(_0531_),
    .B1(_0532_),
    .B2(_0461_),
    .ZN(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1490_ (.A1(_1171_),
    .A2(_0214_),
    .ZN(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1491_ (.I(net13),
    .Z(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1492_ (.A1(_1040_),
    .A2(_0535_),
    .ZN(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _1493_ (.A1(_0531_),
    .A2(_0534_),
    .A3(_0536_),
    .ZN(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1494_ (.A1(_0533_),
    .A2(_0537_),
    .ZN(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1495_ (.A1(_1375_),
    .A2(_1299_),
    .ZN(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1496_ (.A1(_0523_),
    .A2(_0539_),
    .Z(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1497_ (.A1(_1127_),
    .A2(_0375_),
    .ZN(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1498_ (.A1(_0540_),
    .A2(_0541_),
    .Z(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1499_ (.A1(_0538_),
    .A2(_0542_),
    .Z(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _1500_ (.A1(_0528_),
    .A2(_0530_),
    .A3(_0543_),
    .ZN(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1501_ (.A1(_0353_),
    .A2(_0515_),
    .ZN(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1502_ (.A1(_0150_),
    .A2(_0516_),
    .B(_0545_),
    .ZN(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1503_ (.A1(_0544_),
    .A2(_0546_),
    .ZN(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1504_ (.A1(_0522_),
    .A2(_0547_),
    .Z(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1505_ (.A1(_0519_),
    .A2(_0517_),
    .ZN(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1506_ (.A1(_0548_),
    .A2(_0549_),
    .ZN(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1507_ (.I(_0550_),
    .Z(net62));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1508_ (.A1(_1138_),
    .A2(_0375_),
    .A3(_0540_),
    .ZN(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1509_ (.A1(_0523_),
    .A2(_0539_),
    .B(_0551_),
    .ZN(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1510_ (.I(net30),
    .Z(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1511_ (.I(_0553_),
    .Z(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1512_ (.A1(_1138_),
    .A2(_0526_),
    .B1(_0554_),
    .B2(_1181_),
    .ZN(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1513_ (.A1(net8),
    .A2(_0554_),
    .ZN(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1514_ (.A1(_0527_),
    .A2(_0556_),
    .ZN(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1515_ (.A1(_0555_),
    .A2(_0557_),
    .ZN(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1516_ (.A1(_0552_),
    .A2(_0558_),
    .ZN(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1517_ (.A1(_0552_),
    .A2(_0558_),
    .Z(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1518_ (.A1(_0533_),
    .A2(_0537_),
    .ZN(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1519_ (.A1(_0538_),
    .A2(_0542_),
    .B(_0561_),
    .ZN(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1520_ (.A1(_1094_),
    .A2(net13),
    .ZN(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1521_ (.A1(_1105_),
    .A2(_0482_),
    .B1(_0535_),
    .B2(_1051_),
    .ZN(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1522_ (.A1(_0492_),
    .A2(_0563_),
    .B1(_0564_),
    .B2(_0534_),
    .ZN(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1523_ (.A1(_1160_),
    .A2(_0471_),
    .ZN(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1524_ (.I(net14),
    .Z(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1525_ (.I(_0567_),
    .Z(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1526_ (.A1(_1040_),
    .A2(_0568_),
    .ZN(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _1527_ (.A1(_0563_),
    .A2(_0566_),
    .A3(_0569_),
    .ZN(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1528_ (.A1(_0565_),
    .A2(_0570_),
    .ZN(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1529_ (.A1(_1029_),
    .A2(_0375_),
    .ZN(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _1530_ (.A1(_1375_),
    .A2(_1299_),
    .A3(_0225_),
    .A4(_0106_),
    .Z(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1531_ (.A1(_1299_),
    .A2(_0225_),
    .B1(_0106_),
    .B2(_1386_),
    .ZN(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1532_ (.A1(_0573_),
    .A2(_0574_),
    .ZN(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1533_ (.A1(_0572_),
    .A2(_0575_),
    .Z(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1534_ (.A1(_0571_),
    .A2(_0576_),
    .Z(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1535_ (.A1(_0562_),
    .A2(_0577_),
    .Z(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1536_ (.A1(_0562_),
    .A2(_0577_),
    .Z(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1537_ (.A1(_0560_),
    .A2(_0578_),
    .B(_0579_),
    .ZN(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1538_ (.A1(_0572_),
    .A2(_0573_),
    .A3(_0574_),
    .ZN(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1539_ (.A1(_0573_),
    .A2(_0581_),
    .ZN(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1540_ (.I(net31),
    .Z(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1541_ (.I(_0583_),
    .Z(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1542_ (.A1(net1),
    .A2(_0584_),
    .ZN(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1543_ (.A1(net9),
    .A2(_0525_),
    .ZN(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1544_ (.A1(_0556_),
    .A2(_0586_),
    .ZN(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1545_ (.A1(_0585_),
    .A2(_0587_),
    .ZN(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1546_ (.A1(_0582_),
    .A2(_0588_),
    .ZN(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1547_ (.A1(_0557_),
    .A2(_0589_),
    .Z(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1548_ (.A1(_0565_),
    .A2(_0570_),
    .ZN(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1549_ (.A1(_0571_),
    .A2(_0576_),
    .B(_0591_),
    .ZN(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1550_ (.A1(_0214_),
    .A2(_0095_),
    .ZN(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1551_ (.A1(_1375_),
    .A2(_0375_),
    .ZN(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1552_ (.A1(_1288_),
    .A2(_0471_),
    .ZN(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _1553_ (.A1(_0593_),
    .A2(_0594_),
    .A3(_0595_),
    .Z(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1554_ (.A1(_1094_),
    .A2(_0568_),
    .ZN(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1555_ (.I(_0535_),
    .Z(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1556_ (.A1(_1116_),
    .A2(_0598_),
    .B1(_0568_),
    .B2(_1062_),
    .ZN(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1557_ (.A1(_0536_),
    .A2(_0597_),
    .B1(_0599_),
    .B2(_0566_),
    .ZN(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1558_ (.A1(_1171_),
    .A2(_0535_),
    .ZN(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1559_ (.I(net15),
    .Z(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1560_ (.I(_0602_),
    .Z(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1561_ (.A1(_1051_),
    .A2(_0603_),
    .ZN(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _1562_ (.A1(_0597_),
    .A2(_0601_),
    .A3(_0604_),
    .ZN(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1563_ (.A1(_0600_),
    .A2(_0605_),
    .ZN(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1564_ (.A1(_0596_),
    .A2(_0606_),
    .Z(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _1565_ (.A1(_0590_),
    .A2(_0592_),
    .A3(_0607_),
    .Z(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _1566_ (.A1(_0559_),
    .A2(_0580_),
    .A3(_0608_),
    .ZN(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1567_ (.A1(_1192_),
    .A2(_0526_),
    .A3(_0524_),
    .ZN(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1568_ (.A1(_0530_),
    .A2(_0543_),
    .ZN(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1569_ (.A1(_0530_),
    .A2(_0543_),
    .ZN(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1570_ (.A1(_0528_),
    .A2(_0611_),
    .B(_0612_),
    .ZN(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1571_ (.A1(_0560_),
    .A2(_0578_),
    .Z(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1572_ (.A1(_0613_),
    .A2(_0614_),
    .ZN(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1573_ (.A1(_0613_),
    .A2(_0614_),
    .ZN(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1574_ (.A1(_0610_),
    .A2(_0615_),
    .B(_0616_),
    .ZN(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1575_ (.A1(_0544_),
    .A2(_0546_),
    .ZN(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _1576_ (.A1(_0610_),
    .A2(_0613_),
    .A3(_0614_),
    .Z(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1577_ (.A1(_0618_),
    .A2(_0619_),
    .ZN(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _1578_ (.A1(_0609_),
    .A2(_0617_),
    .A3(_0620_),
    .ZN(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _1579_ (.A1(_0518_),
    .A2(_0517_),
    .A3(_0547_),
    .A4(_0619_),
    .Z(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1580_ (.A1(_0621_),
    .A2(_0622_),
    .Z(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1581_ (.A1(_0519_),
    .A2(_0517_),
    .A3(_0548_),
    .ZN(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _1582_ (.A1(_0610_),
    .A2(_0613_),
    .A3(_0614_),
    .ZN(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1583_ (.A1(_0518_),
    .A2(_0517_),
    .A3(_0547_),
    .B(_0618_),
    .ZN(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1584_ (.A1(_0625_),
    .A2(_0626_),
    .Z(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1585_ (.A1(_0624_),
    .A2(_0627_),
    .Z(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1586_ (.A1(_0623_),
    .A2(_0628_),
    .Z(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1587_ (.I(_0629_),
    .Z(net64));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _1588_ (.A1(_0527_),
    .A2(_0556_),
    .A3(_0589_),
    .Z(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1589_ (.A1(_0582_),
    .A2(_0588_),
    .B(_0630_),
    .ZN(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1590_ (.I(net32),
    .Z(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1591_ (.I(_0632_),
    .Z(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1592_ (.A1(_1192_),
    .A2(_0633_),
    .ZN(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1593_ (.A1(_0631_),
    .A2(_0634_),
    .ZN(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1594_ (.A1(_0592_),
    .A2(_0607_),
    .ZN(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1595_ (.A1(_0592_),
    .A2(_0607_),
    .ZN(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1596_ (.A1(_0590_),
    .A2(_0636_),
    .B(_0637_),
    .ZN(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1597_ (.A1(_0556_),
    .A2(_0586_),
    .ZN(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1598_ (.A1(_0585_),
    .A2(_0587_),
    .ZN(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1599_ (.A1(_0639_),
    .A2(_0640_),
    .ZN(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1600_ (.A1(_1299_),
    .A2(_0225_),
    .ZN(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1601_ (.A1(_0095_),
    .A2(_0471_),
    .ZN(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1602_ (.A1(_0593_),
    .A2(_0595_),
    .Z(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1603_ (.A1(_0642_),
    .A2(_0643_),
    .B1(_0644_),
    .B2(_0594_),
    .ZN(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1604_ (.A1(_1018_),
    .A2(_0554_),
    .ZN(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1605_ (.A1(net8),
    .A2(_0584_),
    .ZN(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1606_ (.A1(_1375_),
    .A2(_0526_),
    .ZN(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _1607_ (.A1(_0646_),
    .A2(_0647_),
    .A3(_0648_),
    .Z(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1608_ (.A1(_0645_),
    .A2(_0649_),
    .Z(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1609_ (.A1(_0641_),
    .A2(_0650_),
    .ZN(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1610_ (.A1(_0600_),
    .A2(_0605_),
    .ZN(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1611_ (.A1(_0596_),
    .A2(_0606_),
    .B(_0652_),
    .ZN(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1612_ (.A1(_0214_),
    .A2(_0375_),
    .ZN(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1613_ (.A1(_1288_),
    .A2(net13),
    .ZN(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _1614_ (.A1(_0643_),
    .A2(_0654_),
    .A3(_0655_),
    .Z(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1615_ (.A1(_1084_),
    .A2(_0602_),
    .ZN(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1616_ (.A1(_1040_),
    .A2(_0603_),
    .B1(_0568_),
    .B2(_1105_),
    .ZN(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1617_ (.A1(_0569_),
    .A2(_0657_),
    .B1(_0658_),
    .B2(_0601_),
    .ZN(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1618_ (.A1(_1160_),
    .A2(_0567_),
    .ZN(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1619_ (.I(net16),
    .Z(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1620_ (.A1(_1040_),
    .A2(_0661_),
    .ZN(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _1621_ (.A1(_0657_),
    .A2(_0660_),
    .A3(_0662_),
    .ZN(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1622_ (.A1(_0659_),
    .A2(_0663_),
    .ZN(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1623_ (.A1(_0656_),
    .A2(_0664_),
    .Z(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _1624_ (.A1(_0651_),
    .A2(_0653_),
    .A3(_0665_),
    .ZN(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1625_ (.A1(_0638_),
    .A2(_0666_),
    .Z(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1626_ (.A1(_0635_),
    .A2(_0667_),
    .Z(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1627_ (.A1(_0580_),
    .A2(_0608_),
    .Z(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1628_ (.A1(_0580_),
    .A2(_0608_),
    .Z(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1629_ (.A1(_0559_),
    .A2(_0669_),
    .B(_0670_),
    .ZN(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1630_ (.A1(_0668_),
    .A2(_0671_),
    .Z(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1631_ (.A1(_0609_),
    .A2(_0617_),
    .Z(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1632_ (.A1(_0609_),
    .A2(_0617_),
    .Z(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1633_ (.A1(_0673_),
    .A2(_0620_),
    .B(_0674_),
    .ZN(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1634_ (.A1(_0672_),
    .A2(_0675_),
    .Z(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1635_ (.A1(_0621_),
    .A2(_0622_),
    .Z(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1636_ (.A1(_0623_),
    .A2(_0628_),
    .ZN(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1637_ (.A1(_0677_),
    .A2(_0678_),
    .ZN(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1638_ (.A1(_0676_),
    .A2(_0679_),
    .ZN(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1639_ (.I(_0680_),
    .Z(net65));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1640_ (.A1(_0673_),
    .A2(_0620_),
    .A3(_0672_),
    .ZN(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1641_ (.A1(_0677_),
    .A2(_0681_),
    .Z(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _1642_ (.A1(_0681_),
    .A2(_0676_),
    .B1(_0682_),
    .B2(_0678_),
    .ZN(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1643_ (.A1(_1192_),
    .A2(_0633_),
    .A3(_0631_),
    .ZN(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1644_ (.A1(_0638_),
    .A2(_0666_),
    .Z(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1645_ (.A1(_0635_),
    .A2(_0667_),
    .B(_0685_),
    .ZN(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1646_ (.I(_0649_),
    .ZN(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1647_ (.A1(_0645_),
    .A2(_0687_),
    .ZN(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1648_ (.A1(_0641_),
    .A2(_0650_),
    .B(_0688_),
    .ZN(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1649_ (.A1(_1127_),
    .A2(_0633_),
    .ZN(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1650_ (.I(net18),
    .Z(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1651_ (.I(_0691_),
    .Z(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1652_ (.A1(_1181_),
    .A2(_0692_),
    .ZN(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _1653_ (.A1(_1138_),
    .A2(_1181_),
    .A3(_0633_),
    .A4(_0692_),
    .ZN(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1654_ (.I(_0694_),
    .ZN(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1655_ (.A1(_0690_),
    .A2(_0693_),
    .B(_0695_),
    .ZN(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1656_ (.A1(_0689_),
    .A2(_0696_),
    .Z(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1657_ (.A1(_0653_),
    .A2(_0665_),
    .ZN(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1658_ (.A1(_0653_),
    .A2(_0665_),
    .ZN(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1659_ (.A1(_0651_),
    .A2(_0698_),
    .B(_0699_),
    .ZN(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1660_ (.A1(net10),
    .A2(_0553_),
    .ZN(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1661_ (.A1(_0646_),
    .A2(_0648_),
    .Z(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1662_ (.A1(_0586_),
    .A2(_0701_),
    .B1(_0702_),
    .B2(_0647_),
    .ZN(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1663_ (.A1(_0095_),
    .A2(_0535_),
    .ZN(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1664_ (.A1(_0643_),
    .A2(_0655_),
    .Z(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1665_ (.A1(_0595_),
    .A2(_0704_),
    .B1(_0705_),
    .B2(_0654_),
    .ZN(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1666_ (.A1(net11),
    .A2(_0525_),
    .ZN(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1667_ (.A1(_0701_),
    .A2(_0707_),
    .ZN(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1668_ (.A1(_1018_),
    .A2(_0584_),
    .ZN(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1669_ (.A1(_0708_),
    .A2(_0709_),
    .ZN(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1670_ (.A1(_0706_),
    .A2(_0710_),
    .Z(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1671_ (.A1(_0703_),
    .A2(_0711_),
    .Z(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1672_ (.A1(_0659_),
    .A2(_0663_),
    .ZN(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1673_ (.A1(_0656_),
    .A2(_0664_),
    .B(_0713_),
    .ZN(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1674_ (.A1(_0482_),
    .A2(_0375_),
    .ZN(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1675_ (.A1(_1288_),
    .A2(_0568_),
    .ZN(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _1676_ (.A1(_0704_),
    .A2(_0715_),
    .A3(_0716_),
    .Z(_0717_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1677_ (.A1(_1094_),
    .A2(_0661_),
    .ZN(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1678_ (.I(_0661_),
    .Z(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1679_ (.A1(_1105_),
    .A2(_0603_),
    .B1(_0719_),
    .B2(_1051_),
    .ZN(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1680_ (.A1(_0604_),
    .A2(_0718_),
    .B1(_0720_),
    .B2(_0660_),
    .ZN(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1681_ (.A1(_1171_),
    .A2(_0602_),
    .ZN(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1682_ (.I(net2),
    .Z(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1683_ (.I(_0723_),
    .Z(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1684_ (.A1(_1040_),
    .A2(_0724_),
    .ZN(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _1685_ (.A1(_0718_),
    .A2(_0722_),
    .A3(_0725_),
    .ZN(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1686_ (.A1(_0721_),
    .A2(_0726_),
    .ZN(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1687_ (.A1(_0717_),
    .A2(_0727_),
    .Z(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _1688_ (.A1(_0712_),
    .A2(_0714_),
    .A3(_0728_),
    .ZN(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1689_ (.A1(_0700_),
    .A2(_0729_),
    .Z(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1690_ (.A1(_0697_),
    .A2(_0730_),
    .ZN(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1691_ (.A1(_0686_),
    .A2(_0731_),
    .ZN(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1692_ (.A1(_0684_),
    .A2(_0732_),
    .ZN(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1693_ (.A1(_0668_),
    .A2(_0671_),
    .ZN(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1694_ (.A1(_0674_),
    .A2(_0672_),
    .ZN(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1695_ (.A1(_0734_),
    .A2(_0735_),
    .ZN(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1696_ (.A1(_0733_),
    .A2(_0736_),
    .ZN(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1697_ (.A1(_0683_),
    .A2(_0737_),
    .Z(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1698_ (.I(_0738_),
    .Z(net35));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1699_ (.A1(_0689_),
    .A2(_0696_),
    .ZN(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1700_ (.A1(_0700_),
    .A2(_0729_),
    .Z(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1701_ (.A1(_0697_),
    .A2(_0730_),
    .B(_0740_),
    .ZN(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1702_ (.I(_0703_),
    .ZN(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1703_ (.I(_0710_),
    .ZN(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1704_ (.A1(_0706_),
    .A2(_0743_),
    .ZN(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1705_ (.A1(_0742_),
    .A2(_0711_),
    .B(_0744_),
    .ZN(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1706_ (.I(net19),
    .Z(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1707_ (.I(_0746_),
    .Z(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1708_ (.A1(net1),
    .A2(_0747_),
    .ZN(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1709_ (.A1(net9),
    .A2(_0691_),
    .ZN(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1710_ (.A1(_0690_),
    .A2(_0749_),
    .ZN(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1711_ (.A1(_1018_),
    .A2(_0633_),
    .B1(_0692_),
    .B2(net8),
    .ZN(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1712_ (.A1(_0750_),
    .A2(_0751_),
    .ZN(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1713_ (.A1(_0748_),
    .A2(_0752_),
    .Z(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1714_ (.A1(_0694_),
    .A2(_0753_),
    .Z(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1715_ (.A1(_0745_),
    .A2(_0754_),
    .Z(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1716_ (.A1(_0714_),
    .A2(_0728_),
    .ZN(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1717_ (.A1(_0714_),
    .A2(_0728_),
    .ZN(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1718_ (.A1(_0712_),
    .A2(_0756_),
    .B(_0757_),
    .ZN(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1719_ (.A1(net11),
    .A2(_0553_),
    .ZN(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1720_ (.A1(_0648_),
    .A2(_0759_),
    .ZN(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1721_ (.A1(_0708_),
    .A2(_0709_),
    .ZN(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1722_ (.A1(_0760_),
    .A2(_0761_),
    .ZN(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1723_ (.A1(_0106_),
    .A2(_0568_),
    .ZN(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1724_ (.A1(_0704_),
    .A2(_0716_),
    .Z(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1725_ (.A1(_0655_),
    .A2(_0763_),
    .B1(_0764_),
    .B2(_0715_),
    .ZN(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1726_ (.A1(net10),
    .A2(_0584_),
    .ZN(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1727_ (.A1(net12),
    .A2(_0525_),
    .ZN(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1728_ (.A1(_0759_),
    .A2(_0767_),
    .ZN(_0768_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1729_ (.A1(_0766_),
    .A2(_0768_),
    .Z(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1730_ (.A1(_0765_),
    .A2(_0769_),
    .ZN(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1731_ (.A1(_0762_),
    .A2(_0770_),
    .ZN(_0771_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1732_ (.A1(_0721_),
    .A2(_0726_),
    .ZN(_0772_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1733_ (.A1(_0717_),
    .A2(_0727_),
    .B(_0772_),
    .ZN(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1734_ (.A1(_0375_),
    .A2(_0598_),
    .ZN(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1735_ (.A1(_1288_),
    .A2(_0603_),
    .ZN(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _1736_ (.A1(_0763_),
    .A2(_0774_),
    .A3(_0775_),
    .Z(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1737_ (.A1(_1094_),
    .A2(_0724_),
    .ZN(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1738_ (.A1(_1105_),
    .A2(_0719_),
    .B1(_0724_),
    .B2(_1062_),
    .ZN(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1739_ (.A1(_0662_),
    .A2(_0777_),
    .B1(_0778_),
    .B2(_0722_),
    .ZN(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1740_ (.A1(_1171_),
    .A2(_0719_),
    .ZN(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1741_ (.I(net3),
    .Z(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1742_ (.I(_0781_),
    .Z(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1743_ (.A1(_1040_),
    .A2(_0782_),
    .ZN(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _1744_ (.A1(_0777_),
    .A2(_0780_),
    .A3(_0783_),
    .ZN(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1745_ (.A1(_0779_),
    .A2(_0784_),
    .ZN(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1746_ (.A1(_0776_),
    .A2(_0785_),
    .Z(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _1747_ (.A1(_0771_),
    .A2(_0773_),
    .A3(_0786_),
    .ZN(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1748_ (.A1(_0758_),
    .A2(_0787_),
    .Z(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1749_ (.A1(_0755_),
    .A2(_0788_),
    .ZN(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _1750_ (.A1(_0739_),
    .A2(_0741_),
    .A3(_0789_),
    .ZN(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1751_ (.A1(_0686_),
    .A2(_0731_),
    .Z(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1752_ (.A1(_0684_),
    .A2(_0732_),
    .B(_0791_),
    .ZN(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1753_ (.A1(_0790_),
    .A2(_0792_),
    .Z(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1754_ (.A1(_0734_),
    .A2(_0733_),
    .ZN(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1755_ (.A1(_0735_),
    .A2(_0733_),
    .ZN(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1756_ (.A1(_0683_),
    .A2(_0737_),
    .B(_0795_),
    .ZN(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _1757_ (.A1(_0793_),
    .A2(_0794_),
    .A3(_0796_),
    .ZN(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1758_ (.I(_0797_),
    .Z(net36));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1759_ (.A1(_0683_),
    .A2(_0737_),
    .A3(_0793_),
    .Z(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1760_ (.A1(_0793_),
    .A2(_0794_),
    .ZN(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1761_ (.A1(_0793_),
    .A2(_0794_),
    .B(_0795_),
    .ZN(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1762_ (.A1(_0799_),
    .A2(_0800_),
    .ZN(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1763_ (.A1(_0798_),
    .A2(_0801_),
    .ZN(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1764_ (.A1(_0790_),
    .A2(_0792_),
    .Z(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1765_ (.A1(_0741_),
    .A2(_0789_),
    .Z(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1766_ (.A1(_0741_),
    .A2(_0789_),
    .Z(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1767_ (.A1(_0739_),
    .A2(_0804_),
    .B(_0805_),
    .ZN(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1768_ (.A1(_0745_),
    .A2(_0754_),
    .ZN(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1769_ (.A1(_0758_),
    .A2(_0787_),
    .Z(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1770_ (.A1(_0755_),
    .A2(_0788_),
    .B(_0808_),
    .ZN(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1771_ (.A1(_0694_),
    .A2(_0753_),
    .ZN(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1772_ (.A1(_0765_),
    .A2(_0769_),
    .ZN(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1773_ (.A1(_0762_),
    .A2(_0770_),
    .B(_0811_),
    .ZN(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1774_ (.I(net20),
    .Z(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1775_ (.I(_0813_),
    .Z(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1776_ (.A1(_1181_),
    .A2(_0814_),
    .ZN(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1777_ (.A1(_0690_),
    .A2(_0749_),
    .B1(_0751_),
    .B2(_0748_),
    .ZN(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1778_ (.I(_0816_),
    .ZN(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1779_ (.A1(net8),
    .A2(_0746_),
    .ZN(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1780_ (.A1(_1375_),
    .A2(_0632_),
    .ZN(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _1781_ (.A1(_0749_),
    .A2(_0818_),
    .A3(_0819_),
    .Z(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1782_ (.A1(_0817_),
    .A2(_0820_),
    .Z(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1783_ (.A1(_0815_),
    .A2(_0821_),
    .ZN(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1784_ (.A1(_0812_),
    .A2(_0822_),
    .Z(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1785_ (.A1(_0810_),
    .A2(_0823_),
    .ZN(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1786_ (.A1(_0773_),
    .A2(_0786_),
    .ZN(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1787_ (.A1(_0773_),
    .A2(_0786_),
    .ZN(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1788_ (.A1(_0771_),
    .A2(_0825_),
    .B(_0826_),
    .ZN(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1789_ (.A1(_0471_),
    .A2(_0554_),
    .ZN(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1790_ (.A1(_0707_),
    .A2(_0828_),
    .B1(_0768_),
    .B2(_0766_),
    .ZN(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1791_ (.A1(_0106_),
    .A2(_0603_),
    .ZN(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1792_ (.A1(_0763_),
    .A2(_0775_),
    .Z(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1793_ (.A1(_0716_),
    .A2(_0830_),
    .B1(_0831_),
    .B2(_0774_),
    .ZN(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1794_ (.A1(net11),
    .A2(_0584_),
    .Z(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1795_ (.A1(_0535_),
    .A2(_0526_),
    .ZN(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _1796_ (.A1(_0828_),
    .A2(_0833_),
    .A3(_0834_),
    .Z(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1797_ (.A1(_0832_),
    .A2(_0835_),
    .ZN(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1798_ (.A1(_0829_),
    .A2(_0836_),
    .Z(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1799_ (.A1(_0779_),
    .A2(_0784_),
    .ZN(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1800_ (.A1(_0776_),
    .A2(_0785_),
    .B(_0838_),
    .ZN(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1801_ (.A1(_0364_),
    .A2(_0568_),
    .ZN(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1802_ (.A1(_1288_),
    .A2(_0719_),
    .ZN(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _1803_ (.A1(_0830_),
    .A2(_0840_),
    .A3(_0841_),
    .Z(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1804_ (.A1(_1094_),
    .A2(_0781_),
    .ZN(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1805_ (.A1(_1105_),
    .A2(_0724_),
    .B1(_0782_),
    .B2(_1051_),
    .ZN(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1806_ (.A1(_0725_),
    .A2(_0843_),
    .B1(_0844_),
    .B2(_0780_),
    .ZN(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1807_ (.A1(_1160_),
    .A2(_0723_),
    .ZN(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1808_ (.I(net4),
    .Z(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1809_ (.I(_0847_),
    .Z(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1810_ (.A1(net17),
    .A2(_0848_),
    .ZN(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _1811_ (.A1(_0843_),
    .A2(_0846_),
    .A3(_0849_),
    .ZN(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1812_ (.A1(_0845_),
    .A2(_0850_),
    .ZN(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1813_ (.A1(_0842_),
    .A2(_0851_),
    .Z(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _1814_ (.A1(_0837_),
    .A2(_0839_),
    .A3(_0852_),
    .ZN(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _1815_ (.A1(_0824_),
    .A2(_0827_),
    .A3(_0853_),
    .Z(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _1816_ (.A1(_0807_),
    .A2(_0809_),
    .A3(_0854_),
    .ZN(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1817_ (.A1(_0806_),
    .A2(_0855_),
    .Z(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1818_ (.A1(_0803_),
    .A2(_0856_),
    .ZN(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1819_ (.A1(_0802_),
    .A2(_0857_),
    .Z(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1820_ (.I(_0858_),
    .Z(net37));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1821_ (.A1(_0803_),
    .A2(_0856_),
    .ZN(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1822_ (.A1(_0802_),
    .A2(_0857_),
    .B(_0859_),
    .ZN(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1823_ (.A1(_0806_),
    .A2(_0855_),
    .ZN(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1824_ (.A1(_0812_),
    .A2(_0822_),
    .ZN(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1825_ (.A1(_0810_),
    .A2(_0823_),
    .ZN(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1826_ (.A1(_0862_),
    .A2(_0863_),
    .ZN(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1827_ (.A1(_0827_),
    .A2(_0853_),
    .ZN(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1828_ (.A1(_0827_),
    .A2(_0853_),
    .ZN(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1829_ (.A1(_0824_),
    .A2(_0865_),
    .B(_0866_),
    .ZN(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1830_ (.A1(_0839_),
    .A2(_0852_),
    .ZN(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1831_ (.A1(_0839_),
    .A2(_0852_),
    .ZN(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1832_ (.A1(_0837_),
    .A2(_0868_),
    .B(_0869_),
    .ZN(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1833_ (.A1(_0828_),
    .A2(_0834_),
    .ZN(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1834_ (.A1(net13),
    .A2(_0554_),
    .ZN(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1835_ (.A1(_0767_),
    .A2(_0872_),
    .ZN(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1836_ (.A1(_0833_),
    .A2(_0871_),
    .B(_0873_),
    .ZN(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1837_ (.A1(_0095_),
    .A2(_0661_),
    .ZN(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1838_ (.A1(_0095_),
    .A2(_0603_),
    .B1(_0719_),
    .B2(_1288_),
    .ZN(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1839_ (.A1(_0775_),
    .A2(_0875_),
    .B1(_0876_),
    .B2(_0840_),
    .ZN(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1840_ (.A1(net12),
    .A2(_0583_),
    .ZN(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1841_ (.A1(_0526_),
    .A2(_0567_),
    .ZN(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _1842_ (.A1(_0872_),
    .A2(_0878_),
    .A3(_0879_),
    .ZN(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1843_ (.A1(_0877_),
    .A2(_0880_),
    .ZN(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1844_ (.A1(_0874_),
    .A2(_0881_),
    .ZN(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1845_ (.A1(_0845_),
    .A2(_0850_),
    .ZN(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1846_ (.A1(_0842_),
    .A2(_0851_),
    .B(_0883_),
    .ZN(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1847_ (.A1(_0364_),
    .A2(_0603_),
    .ZN(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1848_ (.A1(_1288_),
    .A2(_0723_),
    .ZN(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _1849_ (.A1(_0875_),
    .A2(_0885_),
    .A3(_0886_),
    .Z(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1850_ (.A1(_1084_),
    .A2(_0847_),
    .ZN(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1851_ (.A1(_1094_),
    .A2(_0782_),
    .B1(_0848_),
    .B2(_1040_),
    .ZN(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1852_ (.A1(_0783_),
    .A2(_0888_),
    .B1(_0889_),
    .B2(_0846_),
    .ZN(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1853_ (.A1(_1160_),
    .A2(net3),
    .ZN(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1854_ (.I(net5),
    .Z(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1855_ (.I(_0892_),
    .Z(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1856_ (.A1(net17),
    .A2(_0893_),
    .ZN(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _1857_ (.A1(_0888_),
    .A2(_0891_),
    .A3(_0894_),
    .ZN(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1858_ (.A1(_0890_),
    .A2(_0895_),
    .ZN(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1859_ (.A1(_0887_),
    .A2(_0896_),
    .Z(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _1860_ (.A1(_0882_),
    .A2(_0884_),
    .A3(_0897_),
    .ZN(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1861_ (.A1(_0870_),
    .A2(_0898_),
    .ZN(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1862_ (.A1(_1181_),
    .A2(_0814_),
    .A3(_0821_),
    .ZN(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1863_ (.A1(_0817_),
    .A2(_0820_),
    .B(_0900_),
    .ZN(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1864_ (.I(_0829_),
    .ZN(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1865_ (.A1(_0832_),
    .A2(_0835_),
    .ZN(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1866_ (.A1(_0902_),
    .A2(_0836_),
    .B(_0903_),
    .ZN(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1867_ (.I(net21),
    .Z(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1868_ (.I(_0905_),
    .Z(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1869_ (.A1(_1127_),
    .A2(_0814_),
    .B1(_0906_),
    .B2(net1),
    .ZN(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _1870_ (.A1(_1127_),
    .A2(net1),
    .A3(_0814_),
    .A4(_0906_),
    .ZN(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1871_ (.I(_0908_),
    .ZN(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1872_ (.A1(_0907_),
    .A2(_0909_),
    .ZN(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1873_ (.A1(_1029_),
    .A2(_0633_),
    .ZN(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1874_ (.A1(net10),
    .A2(_0691_),
    .ZN(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1875_ (.A1(_1386_),
    .A2(_0633_),
    .B1(_0692_),
    .B2(_1018_),
    .ZN(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1876_ (.A1(_0911_),
    .A2(_0912_),
    .B1(_0913_),
    .B2(_0818_),
    .ZN(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1877_ (.A1(_1018_),
    .A2(_0747_),
    .ZN(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1878_ (.A1(net11),
    .A2(_0632_),
    .ZN(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _1879_ (.A1(_0912_),
    .A2(_0915_),
    .A3(_0916_),
    .ZN(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1880_ (.A1(_0914_),
    .A2(_0917_),
    .Z(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1881_ (.A1(_0910_),
    .A2(_0918_),
    .Z(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1882_ (.A1(_0904_),
    .A2(_0919_),
    .Z(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1883_ (.A1(_0901_),
    .A2(_0920_),
    .ZN(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1884_ (.A1(_0899_),
    .A2(_0921_),
    .Z(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _1885_ (.A1(_0864_),
    .A2(_0867_),
    .A3(_0922_),
    .ZN(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1886_ (.I(_0923_),
    .ZN(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1887_ (.A1(_0809_),
    .A2(_0854_),
    .Z(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1888_ (.A1(_0809_),
    .A2(_0854_),
    .Z(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1889_ (.A1(_0807_),
    .A2(_0925_),
    .B(_0926_),
    .ZN(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _1890_ (.A1(_0861_),
    .A2(_0924_),
    .A3(_0927_),
    .Z(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1891_ (.A1(_0860_),
    .A2(_0928_),
    .ZN(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1892_ (.I(_0929_),
    .Z(net38));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1893_ (.A1(_0924_),
    .A2(_0927_),
    .Z(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1894_ (.A1(_0867_),
    .A2(_0922_),
    .Z(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1895_ (.A1(_0867_),
    .A2(_0922_),
    .Z(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1896_ (.A1(_0864_),
    .A2(_0931_),
    .B(_0932_),
    .ZN(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1897_ (.A1(_0901_),
    .A2(_0920_),
    .Z(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1898_ (.A1(_0904_),
    .A2(_0919_),
    .B(_0934_),
    .ZN(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1899_ (.A1(_0908_),
    .A2(_0935_),
    .Z(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1900_ (.A1(_0870_),
    .A2(_0898_),
    .ZN(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1901_ (.A1(_0899_),
    .A2(_0921_),
    .B(_0937_),
    .ZN(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1902_ (.A1(_0914_),
    .A2(_0917_),
    .ZN(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1903_ (.A1(_0910_),
    .A2(_0918_),
    .ZN(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1904_ (.A1(_0939_),
    .A2(_0940_),
    .ZN(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1905_ (.A1(_0877_),
    .A2(_0880_),
    .ZN(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1906_ (.A1(_0874_),
    .A2(_0881_),
    .B(_0942_),
    .ZN(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1907_ (.I(net22),
    .Z(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1908_ (.A1(net1),
    .A2(_0944_),
    .ZN(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1909_ (.A1(net8),
    .A2(_0905_),
    .ZN(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1910_ (.A1(net9),
    .A2(net20),
    .ZN(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1911_ (.A1(_0946_),
    .A2(_0947_),
    .ZN(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1912_ (.A1(_0945_),
    .A2(_0948_),
    .ZN(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1913_ (.A1(net11),
    .A2(_0691_),
    .ZN(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1914_ (.A1(_0214_),
    .A2(_0633_),
    .B1(_0692_),
    .B2(_1375_),
    .ZN(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1915_ (.A1(_0819_),
    .A2(_0950_),
    .B1(_0951_),
    .B2(_0915_),
    .ZN(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1916_ (.A1(net10),
    .A2(_0746_),
    .ZN(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1917_ (.A1(_0471_),
    .A2(_0632_),
    .ZN(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _1918_ (.A1(_0950_),
    .A2(_0953_),
    .A3(_0954_),
    .Z(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1919_ (.A1(_0952_),
    .A2(_0955_),
    .Z(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1920_ (.A1(_0949_),
    .A2(_0956_),
    .Z(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1921_ (.A1(_0943_),
    .A2(_0957_),
    .Z(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1922_ (.A1(_0941_),
    .A2(_0958_),
    .ZN(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1923_ (.A1(_0884_),
    .A2(_0897_),
    .ZN(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1924_ (.A1(_0884_),
    .A2(_0897_),
    .ZN(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1925_ (.A1(_0882_),
    .A2(_0960_),
    .B(_0961_),
    .ZN(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1926_ (.A1(net14),
    .A2(_0553_),
    .ZN(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1927_ (.A1(_0872_),
    .A2(_0879_),
    .Z(_0964_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1928_ (.A1(_0834_),
    .A2(_0963_),
    .B1(_0964_),
    .B2(_0878_),
    .ZN(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1929_ (.A1(net27),
    .A2(_0723_),
    .ZN(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1930_ (.A1(_0875_),
    .A2(_0886_),
    .Z(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1931_ (.A1(_0841_),
    .A2(_0966_),
    .B1(_0967_),
    .B2(_0885_),
    .ZN(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1932_ (.A1(net13),
    .A2(_0584_),
    .ZN(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1933_ (.A1(_0525_),
    .A2(_0602_),
    .ZN(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1934_ (.A1(_0963_),
    .A2(_0970_),
    .ZN(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1935_ (.A1(_0969_),
    .A2(_0971_),
    .Z(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1936_ (.A1(_0968_),
    .A2(_0972_),
    .ZN(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1937_ (.A1(_0965_),
    .A2(_0973_),
    .Z(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1938_ (.A1(_0890_),
    .A2(_0895_),
    .ZN(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1939_ (.A1(_0887_),
    .A2(_0896_),
    .B(_0975_),
    .ZN(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1940_ (.A1(_0364_),
    .A2(_0661_),
    .ZN(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1941_ (.A1(net26),
    .A2(_0781_),
    .ZN(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _1942_ (.A1(_0966_),
    .A2(_0977_),
    .A3(_0978_),
    .Z(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1943_ (.A1(_1084_),
    .A2(_0892_),
    .ZN(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1944_ (.A1(_1084_),
    .A2(_0847_),
    .B1(_0893_),
    .B2(net17),
    .ZN(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1945_ (.A1(_0849_),
    .A2(_0980_),
    .B1(_0981_),
    .B2(_0891_),
    .ZN(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1946_ (.A1(_1160_),
    .A2(net4),
    .ZN(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1947_ (.I(net6),
    .Z(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1948_ (.A1(net17),
    .A2(_0984_),
    .ZN(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _1949_ (.A1(_0980_),
    .A2(_0983_),
    .A3(_0985_),
    .ZN(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1950_ (.A1(_0982_),
    .A2(_0986_),
    .ZN(_0987_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1951_ (.A1(_0979_),
    .A2(_0987_),
    .Z(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1952_ (.A1(_0976_),
    .A2(_0988_),
    .ZN(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1953_ (.A1(_0974_),
    .A2(_0989_),
    .Z(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1954_ (.A1(_0962_),
    .A2(_0990_),
    .ZN(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1955_ (.A1(_0959_),
    .A2(_0991_),
    .Z(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _1956_ (.A1(_0936_),
    .A2(_0938_),
    .A3(_0992_),
    .ZN(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1957_ (.A1(_0933_),
    .A2(_0993_),
    .Z(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1958_ (.A1(_0930_),
    .A2(_0994_),
    .Z(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1959_ (.A1(_0802_),
    .A2(_0857_),
    .A3(_0928_),
    .ZN(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1960_ (.A1(_0924_),
    .A2(_0927_),
    .ZN(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1961_ (.A1(_0861_),
    .A2(_0859_),
    .B(_0930_),
    .C(_0997_),
    .ZN(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1962_ (.A1(_0996_),
    .A2(_0998_),
    .Z(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1963_ (.A1(_0995_),
    .A2(_0999_),
    .Z(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1964_ (.I(_1000_),
    .Z(net39));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1965_ (.A1(_0930_),
    .A2(_0994_),
    .ZN(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1966_ (.A1(_0995_),
    .A2(_0999_),
    .ZN(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1967_ (.A1(_1001_),
    .A2(_1002_),
    .ZN(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1968_ (.A1(_0908_),
    .A2(_0935_),
    .Z(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1969_ (.A1(_0933_),
    .A2(_0993_),
    .Z(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1970_ (.A1(_0938_),
    .A2(_0992_),
    .Z(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1971_ (.A1(_0938_),
    .A2(_0992_),
    .Z(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1972_ (.A1(_0936_),
    .A2(_1006_),
    .B(_1007_),
    .ZN(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1973_ (.I(net23),
    .Z(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1974_ (.A1(_1192_),
    .A2(_1009_),
    .ZN(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1975_ (.A1(_0943_),
    .A2(_0957_),
    .ZN(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1976_ (.A1(_0941_),
    .A2(_0958_),
    .ZN(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1977_ (.A1(_1011_),
    .A2(_1012_),
    .ZN(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1978_ (.A1(_0946_),
    .A2(_0947_),
    .ZN(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1979_ (.A1(_0945_),
    .A2(_0948_),
    .ZN(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1980_ (.A1(_1014_),
    .A2(_1015_),
    .ZN(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1981_ (.A1(_1013_),
    .A2(_1016_),
    .ZN(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1982_ (.A1(_1010_),
    .A2(_1017_),
    .Z(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1983_ (.A1(_0962_),
    .A2(_0990_),
    .ZN(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1984_ (.A1(_0959_),
    .A2(_0991_),
    .B(_1020_),
    .ZN(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1985_ (.I(_0955_),
    .ZN(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1986_ (.A1(_0952_),
    .A2(_1022_),
    .ZN(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1987_ (.A1(_0949_),
    .A2(_0956_),
    .B(_1023_),
    .ZN(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1988_ (.I(_0965_),
    .ZN(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1989_ (.A1(_0968_),
    .A2(_0972_),
    .ZN(_1026_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1990_ (.A1(_1025_),
    .A2(_0973_),
    .B(_1026_),
    .ZN(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1991_ (.A1(_1127_),
    .A2(_0944_),
    .ZN(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1992_ (.A1(net10),
    .A2(net21),
    .ZN(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1993_ (.A1(_0947_),
    .A2(_1030_),
    .ZN(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1994_ (.A1(net10),
    .A2(_0813_),
    .B1(_0905_),
    .B2(_1018_),
    .ZN(_1032_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1995_ (.A1(_1031_),
    .A2(_1032_),
    .Z(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1996_ (.A1(_1028_),
    .A2(_1033_),
    .ZN(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1997_ (.A1(net12),
    .A2(_0691_),
    .ZN(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1998_ (.A1(_0950_),
    .A2(_0954_),
    .Z(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1999_ (.A1(_0916_),
    .A2(_1035_),
    .B1(_1036_),
    .B2(_0953_),
    .ZN(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2000_ (.A1(net11),
    .A2(_0746_),
    .ZN(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2001_ (.A1(net13),
    .A2(_0632_),
    .ZN(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2002_ (.A1(_1035_),
    .A2(_1038_),
    .A3(_1039_),
    .Z(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2003_ (.A1(_1037_),
    .A2(_1041_),
    .Z(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2004_ (.A1(_1034_),
    .A2(_1042_),
    .Z(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2005_ (.A1(_1027_),
    .A2(_1043_),
    .Z(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2006_ (.A1(_1024_),
    .A2(_1044_),
    .ZN(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2007_ (.A1(_0976_),
    .A2(_0988_),
    .ZN(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2008_ (.A1(_0974_),
    .A2(_0989_),
    .B(_1046_),
    .ZN(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2009_ (.A1(_0602_),
    .A2(_0553_),
    .ZN(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2010_ (.A1(_0879_),
    .A2(_1048_),
    .B1(_0971_),
    .B2(_0969_),
    .ZN(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2011_ (.A1(net27),
    .A2(net3),
    .ZN(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2012_ (.A1(_0966_),
    .A2(_0978_),
    .Z(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2013_ (.A1(_0886_),
    .A2(_1050_),
    .B1(_1052_),
    .B2(_0977_),
    .ZN(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2014_ (.A1(net14),
    .A2(_0583_),
    .ZN(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2015_ (.A1(_0525_),
    .A2(_0661_),
    .ZN(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _2016_ (.A1(_1048_),
    .A2(_1054_),
    .A3(_1055_),
    .ZN(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2017_ (.A1(_1053_),
    .A2(_1056_),
    .ZN(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2018_ (.A1(_1049_),
    .A2(_1057_),
    .Z(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2019_ (.A1(_0982_),
    .A2(_0986_),
    .ZN(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2020_ (.A1(_0979_),
    .A2(_0987_),
    .B(_1059_),
    .ZN(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2021_ (.A1(net28),
    .A2(net2),
    .ZN(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2022_ (.A1(net26),
    .A2(_0847_),
    .ZN(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2023_ (.A1(_1050_),
    .A2(_1061_),
    .A3(_1063_),
    .Z(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2024_ (.A1(net24),
    .A2(net6),
    .ZN(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2025_ (.I(_0984_),
    .Z(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2026_ (.A1(_1084_),
    .A2(_0892_),
    .B1(_1066_),
    .B2(net17),
    .ZN(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2027_ (.A1(_0894_),
    .A2(_1065_),
    .B1(_1067_),
    .B2(_0983_),
    .ZN(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2028_ (.A1(net25),
    .A2(net5),
    .ZN(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2029_ (.I(net7),
    .Z(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2030_ (.A1(net17),
    .A2(_1070_),
    .ZN(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _2031_ (.A1(_1065_),
    .A2(_1069_),
    .A3(_1071_),
    .ZN(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2032_ (.A1(_1068_),
    .A2(_1072_),
    .ZN(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2033_ (.A1(_1064_),
    .A2(_1074_),
    .Z(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2034_ (.A1(_1060_),
    .A2(_1075_),
    .ZN(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2035_ (.A1(_1058_),
    .A2(_1076_),
    .Z(_1077_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2036_ (.A1(_1047_),
    .A2(_1077_),
    .ZN(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2037_ (.A1(_1045_),
    .A2(_1078_),
    .Z(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2038_ (.A1(_1021_),
    .A2(_1079_),
    .ZN(_1080_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2039_ (.A1(_1019_),
    .A2(_1080_),
    .ZN(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2040_ (.A1(_1008_),
    .A2(_1081_),
    .Z(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2041_ (.A1(_1004_),
    .A2(_1005_),
    .A3(_1082_),
    .Z(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2042_ (.A1(_1003_),
    .A2(_1083_),
    .Z(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2043_ (.I(_1085_),
    .Z(net40));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2044_ (.A1(_1014_),
    .A2(_1015_),
    .B(_1013_),
    .ZN(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2045_ (.I(_1009_),
    .Z(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2046_ (.A1(_1192_),
    .A2(_1087_),
    .A3(_1017_),
    .ZN(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2047_ (.A1(_1086_),
    .A2(_1088_),
    .ZN(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2048_ (.A1(_1021_),
    .A2(_1079_),
    .ZN(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2049_ (.A1(_1019_),
    .A2(_1080_),
    .B(_1090_),
    .ZN(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2050_ (.A1(_1027_),
    .A2(_1043_),
    .Z(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2051_ (.A1(_1024_),
    .A2(_1044_),
    .B(_1092_),
    .ZN(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2052_ (.A1(_1028_),
    .A2(_1033_),
    .ZN(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2053_ (.A1(_1031_),
    .A2(_1095_),
    .ZN(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2054_ (.A1(_1093_),
    .A2(_1096_),
    .ZN(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2055_ (.A1(_1047_),
    .A2(_1077_),
    .ZN(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2056_ (.A1(_1045_),
    .A2(_1078_),
    .B(_1098_),
    .ZN(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2057_ (.I(_1041_),
    .ZN(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2058_ (.A1(_1037_),
    .A2(_1100_),
    .ZN(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2059_ (.A1(_1034_),
    .A2(_1042_),
    .B(_1101_),
    .ZN(_1102_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2060_ (.I(_1049_),
    .ZN(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2061_ (.A1(_1053_),
    .A2(_1056_),
    .ZN(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2062_ (.A1(_1103_),
    .A2(_1057_),
    .B(_1104_),
    .ZN(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2063_ (.A1(_1127_),
    .A2(net23),
    .ZN(_1107_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2064_ (.A1(net9),
    .A2(net22),
    .ZN(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2065_ (.A1(_1030_),
    .A2(_1108_),
    .ZN(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2066_ (.A1(_1107_),
    .A2(_1109_),
    .ZN(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2067_ (.A1(net13),
    .A2(_0691_),
    .ZN(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2068_ (.A1(_1035_),
    .A2(_1039_),
    .Z(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _2069_ (.A1(_0954_),
    .A2(_1111_),
    .B1(_1112_),
    .B2(_1038_),
    .ZN(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2070_ (.A1(_0214_),
    .A2(_0813_),
    .ZN(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2071_ (.A1(net12),
    .A2(_0746_),
    .ZN(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2072_ (.A1(_1111_),
    .A2(_1115_),
    .ZN(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2073_ (.A1(_1114_),
    .A2(_1117_),
    .Z(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _2074_ (.A1(_1110_),
    .A2(_1113_),
    .A3(_1118_),
    .ZN(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _2075_ (.A1(_1102_),
    .A2(_1106_),
    .A3(_1119_),
    .ZN(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2076_ (.A1(_1060_),
    .A2(_1075_),
    .ZN(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2077_ (.A1(_1058_),
    .A2(_1076_),
    .B(_1121_),
    .ZN(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2078_ (.A1(net30),
    .A2(net16),
    .ZN(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2079_ (.A1(_1048_),
    .A2(_1055_),
    .Z(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2080_ (.A1(_0970_),
    .A2(_1123_),
    .B1(_1124_),
    .B2(_1054_),
    .ZN(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2081_ (.A1(net27),
    .A2(net4),
    .ZN(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2082_ (.A1(_1050_),
    .A2(_1063_),
    .Z(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2083_ (.A1(_0978_),
    .A2(_1126_),
    .B1(_1128_),
    .B2(_1061_),
    .ZN(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2084_ (.A1(net14),
    .A2(net32),
    .ZN(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2085_ (.A1(_0602_),
    .A2(_0583_),
    .ZN(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _2086_ (.A1(_1123_),
    .A2(_1130_),
    .A3(_1131_),
    .ZN(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2087_ (.A1(_1129_),
    .A2(_1132_),
    .ZN(_1133_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2088_ (.A1(_1125_),
    .A2(_1133_),
    .Z(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2089_ (.A1(_1068_),
    .A2(_1072_),
    .ZN(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2090_ (.A1(_1064_),
    .A2(_1074_),
    .B(_1135_),
    .ZN(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2091_ (.A1(net29),
    .A2(net2),
    .ZN(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2092_ (.A1(net28),
    .A2(_0781_),
    .ZN(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2093_ (.A1(_1126_),
    .A2(_1137_),
    .A3(_1139_),
    .Z(_1140_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2094_ (.A1(net24),
    .A2(net7),
    .ZN(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2095_ (.A1(_1084_),
    .A2(_0984_),
    .B1(_1070_),
    .B2(net17),
    .ZN(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2096_ (.A1(_0985_),
    .A2(_1141_),
    .B1(_1142_),
    .B2(_1069_),
    .ZN(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2097_ (.A1(net26),
    .A2(net5),
    .ZN(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2098_ (.A1(net25),
    .A2(net6),
    .ZN(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _2099_ (.A1(_1141_),
    .A2(_1144_),
    .A3(_1145_),
    .ZN(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2100_ (.A1(_1143_),
    .A2(_1146_),
    .ZN(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2101_ (.A1(_1140_),
    .A2(_1147_),
    .Z(_1148_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2102_ (.A1(_1136_),
    .A2(_1148_),
    .ZN(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2103_ (.A1(_1134_),
    .A2(_1150_),
    .Z(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2104_ (.A1(_1122_),
    .A2(_1151_),
    .ZN(_1152_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2105_ (.A1(_1120_),
    .A2(_1152_),
    .Z(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2106_ (.A1(_1099_),
    .A2(_1153_),
    .ZN(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2107_ (.A1(_1097_),
    .A2(_1154_),
    .Z(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2108_ (.A1(_1091_),
    .A2(_1155_),
    .Z(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2109_ (.A1(_1089_),
    .A2(_1156_),
    .ZN(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2110_ (.I(_1004_),
    .ZN(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2111_ (.A1(_1008_),
    .A2(_1081_),
    .ZN(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2112_ (.A1(_1158_),
    .A2(_1082_),
    .B(_1159_),
    .ZN(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2113_ (.A1(_1157_),
    .A2(_1161_),
    .Z(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2114_ (.A1(_1157_),
    .A2(_1161_),
    .ZN(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2115_ (.A1(_1162_),
    .A2(_1163_),
    .ZN(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2116_ (.A1(_0995_),
    .A2(_1083_),
    .Z(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2117_ (.A1(_1004_),
    .A2(_1082_),
    .Z(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2118_ (.A1(_1004_),
    .A2(_1082_),
    .ZN(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2119_ (.A1(_1005_),
    .A2(_1001_),
    .B1(_1166_),
    .B2(_1167_),
    .ZN(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2120_ (.A1(_0998_),
    .A2(_1165_),
    .B(_1168_),
    .ZN(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2121_ (.A1(_0857_),
    .A2(_0928_),
    .ZN(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _2122_ (.A1(_0798_),
    .A2(_0801_),
    .B(_1170_),
    .C(_1165_),
    .ZN(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2123_ (.A1(_1169_),
    .A2(_1172_),
    .Z(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2124_ (.A1(_1164_),
    .A2(_1173_),
    .Z(_1174_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2125_ (.I(_1174_),
    .Z(net41));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2126_ (.A1(_1091_),
    .A2(_1155_),
    .Z(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2127_ (.A1(_1089_),
    .A2(_1156_),
    .B(_1175_),
    .ZN(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2128_ (.A1(_1093_),
    .A2(_1096_),
    .ZN(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2129_ (.A1(_1099_),
    .A2(_1153_),
    .ZN(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2130_ (.A1(_1097_),
    .A2(_1154_),
    .B(_1178_),
    .ZN(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2131_ (.A1(_1106_),
    .A2(_1119_),
    .Z(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2132_ (.A1(_1106_),
    .A2(_1119_),
    .Z(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2133_ (.A1(_1102_),
    .A2(_1180_),
    .B(_1182_),
    .ZN(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2134_ (.A1(_1030_),
    .A2(_1108_),
    .ZN(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2135_ (.A1(_1107_),
    .A2(_1109_),
    .ZN(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2136_ (.A1(_1184_),
    .A2(_1185_),
    .ZN(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2137_ (.A1(_1183_),
    .A2(_1186_),
    .Z(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2138_ (.A1(_1183_),
    .A2(_1186_),
    .ZN(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2139_ (.A1(_1187_),
    .A2(_1188_),
    .ZN(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2140_ (.A1(_1122_),
    .A2(_1151_),
    .ZN(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2141_ (.A1(_1120_),
    .A2(_1152_),
    .B(_1190_),
    .ZN(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2142_ (.A1(_1113_),
    .A2(_1118_),
    .ZN(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2143_ (.A1(_1113_),
    .A2(_1118_),
    .ZN(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2144_ (.A1(_1110_),
    .A2(_1193_),
    .B(_1194_),
    .ZN(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2145_ (.I(_1125_),
    .ZN(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2146_ (.A1(_1129_),
    .A2(_1132_),
    .ZN(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2147_ (.A1(_1196_),
    .A2(_1133_),
    .B(_1197_),
    .ZN(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2148_ (.I(_0944_),
    .Z(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2149_ (.A1(_1386_),
    .A2(_1199_),
    .B1(net23),
    .B2(_1029_),
    .ZN(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2150_ (.A1(_1386_),
    .A2(net23),
    .ZN(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2151_ (.A1(_1108_),
    .A2(_1201_),
    .ZN(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2152_ (.A1(_1200_),
    .A2(_1202_),
    .ZN(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2153_ (.A1(net13),
    .A2(_0746_),
    .ZN(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2154_ (.A1(_1035_),
    .A2(_1205_),
    .B1(_1117_),
    .B2(_1114_),
    .ZN(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2155_ (.A1(_0214_),
    .A2(_0905_),
    .ZN(_1207_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2156_ (.A1(net12),
    .A2(net20),
    .ZN(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2157_ (.A1(_1205_),
    .A2(_1208_),
    .ZN(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2158_ (.A1(_1207_),
    .A2(_1209_),
    .Z(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2159_ (.A1(_1206_),
    .A2(_1210_),
    .Z(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2160_ (.A1(_1204_),
    .A2(_1211_),
    .Z(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2161_ (.A1(_1198_),
    .A2(_1212_),
    .Z(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2162_ (.A1(_1195_),
    .A2(_1213_),
    .ZN(_1215_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2163_ (.A1(_1136_),
    .A2(_1148_),
    .ZN(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2164_ (.A1(_1134_),
    .A2(_1150_),
    .B(_1216_),
    .ZN(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2165_ (.A1(_0583_),
    .A2(_0661_),
    .ZN(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2166_ (.A1(_1123_),
    .A2(_1131_),
    .Z(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2167_ (.A1(_1048_),
    .A2(_1218_),
    .B1(_1219_),
    .B2(_1130_),
    .ZN(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2168_ (.A1(_0364_),
    .A2(_0847_),
    .ZN(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2169_ (.A1(_1126_),
    .A2(_1139_),
    .Z(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2170_ (.A1(_1050_),
    .A2(_1221_),
    .B1(_1222_),
    .B2(_1137_),
    .ZN(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2171_ (.A1(_0567_),
    .A2(_0691_),
    .ZN(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2172_ (.A1(_0602_),
    .A2(net32),
    .ZN(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2173_ (.A1(_1218_),
    .A2(_1226_),
    .ZN(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2174_ (.A1(_1224_),
    .A2(_1227_),
    .Z(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2175_ (.A1(_1223_),
    .A2(_1228_),
    .ZN(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2176_ (.A1(_1220_),
    .A2(_1229_),
    .Z(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2177_ (.A1(_1143_),
    .A2(_1146_),
    .ZN(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2178_ (.A1(_1140_),
    .A2(_1147_),
    .B(_1231_),
    .ZN(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2179_ (.A1(_0554_),
    .A2(_0723_),
    .ZN(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2180_ (.A1(_0526_),
    .A2(_0782_),
    .ZN(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2181_ (.A1(_1221_),
    .A2(_1233_),
    .A3(_1234_),
    .Z(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2182_ (.A1(net25),
    .A2(_1070_),
    .ZN(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2183_ (.I(_1070_),
    .Z(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2184_ (.A1(_1160_),
    .A2(_1066_),
    .B1(_1237_),
    .B2(_1084_),
    .ZN(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2185_ (.A1(_1065_),
    .A2(_1236_),
    .B1(_1238_),
    .B2(_1144_),
    .ZN(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2186_ (.A1(net27),
    .A2(_0892_),
    .ZN(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2187_ (.A1(net26),
    .A2(_0984_),
    .ZN(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _2188_ (.A1(_1236_),
    .A2(_1240_),
    .A3(_1241_),
    .ZN(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2189_ (.A1(_1239_),
    .A2(_1242_),
    .ZN(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2190_ (.A1(_1235_),
    .A2(_1243_),
    .Z(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2191_ (.A1(_1232_),
    .A2(_1244_),
    .ZN(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2192_ (.A1(_1230_),
    .A2(_1245_),
    .Z(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2193_ (.A1(_1217_),
    .A2(_1247_),
    .ZN(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2194_ (.A1(_1215_),
    .A2(_1248_),
    .Z(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2195_ (.A1(_1191_),
    .A2(_1249_),
    .ZN(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2196_ (.A1(_1189_),
    .A2(_1250_),
    .Z(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2197_ (.A1(_1177_),
    .A2(_1179_),
    .A3(_1251_),
    .Z(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2198_ (.A1(_1176_),
    .A2(_1252_),
    .ZN(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2199_ (.A1(_1164_),
    .A2(_1173_),
    .B(_1162_),
    .ZN(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2200_ (.A1(_1253_),
    .A2(_1254_),
    .Z(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2201_ (.I(_1255_),
    .Z(net42));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2202_ (.A1(_1191_),
    .A2(_1249_),
    .ZN(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2203_ (.A1(_1189_),
    .A2(_1250_),
    .B(_1257_),
    .ZN(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2204_ (.A1(_1198_),
    .A2(_1212_),
    .ZN(_1259_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2205_ (.A1(_1195_),
    .A2(_1213_),
    .ZN(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2206_ (.A1(_1259_),
    .A2(_1260_),
    .ZN(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2207_ (.A1(_1202_),
    .A2(_1261_),
    .ZN(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2208_ (.A1(_1217_),
    .A2(_1247_),
    .ZN(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2209_ (.A1(_1215_),
    .A2(_1248_),
    .B(_1263_),
    .ZN(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2210_ (.A1(_1206_),
    .A2(_1210_),
    .B1(_1211_),
    .B2(_1204_),
    .ZN(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2211_ (.I(_1220_),
    .ZN(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2212_ (.A1(_1223_),
    .A2(_1228_),
    .ZN(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2213_ (.A1(_1266_),
    .A2(_1229_),
    .B(_1267_),
    .ZN(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2214_ (.A1(_0598_),
    .A2(_0814_),
    .ZN(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _2215_ (.A1(_1115_),
    .A2(_1269_),
    .B1(_1209_),
    .B2(_1207_),
    .ZN(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2216_ (.A1(_0225_),
    .A2(_1199_),
    .ZN(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2217_ (.A1(_0482_),
    .A2(_0535_),
    .A3(_0813_),
    .A4(_0905_),
    .Z(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2218_ (.A1(_0598_),
    .A2(_0813_),
    .B1(_0906_),
    .B2(_0482_),
    .ZN(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2219_ (.A1(_1272_),
    .A2(_1273_),
    .Z(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2220_ (.A1(_1271_),
    .A2(_1274_),
    .ZN(_1275_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2221_ (.A1(_1201_),
    .A2(_1270_),
    .A3(_1275_),
    .Z(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2222_ (.A1(_1265_),
    .A2(_1268_),
    .A3(_1276_),
    .Z(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2223_ (.A1(_1232_),
    .A2(_1244_),
    .ZN(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2224_ (.A1(_1230_),
    .A2(_1245_),
    .B(_1279_),
    .ZN(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2225_ (.A1(_0661_),
    .A2(net32),
    .ZN(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2226_ (.A1(_1131_),
    .A2(_1281_),
    .B1(_1227_),
    .B2(_1224_),
    .ZN(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2227_ (.A1(_0526_),
    .A2(_0847_),
    .ZN(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2228_ (.A1(_1221_),
    .A2(_1234_),
    .Z(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2229_ (.A1(_1139_),
    .A2(_1283_),
    .B1(_1284_),
    .B2(_1233_),
    .ZN(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2230_ (.A1(_0567_),
    .A2(_0747_),
    .ZN(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2231_ (.A1(_0602_),
    .A2(_0691_),
    .ZN(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2232_ (.A1(_1281_),
    .A2(_1287_),
    .ZN(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2233_ (.A1(_1286_),
    .A2(_1289_),
    .Z(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2234_ (.A1(_1285_),
    .A2(_1290_),
    .ZN(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2235_ (.A1(_1282_),
    .A2(_1291_),
    .Z(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2236_ (.A1(_1239_),
    .A2(_1242_),
    .ZN(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2237_ (.A1(_1235_),
    .A2(_1243_),
    .B(_1293_),
    .ZN(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2238_ (.A1(_0584_),
    .A2(_0723_),
    .ZN(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2239_ (.A1(_0554_),
    .A2(_0781_),
    .ZN(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2240_ (.A1(_1283_),
    .A2(_1295_),
    .A3(_1296_),
    .Z(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2241_ (.A1(net26),
    .A2(_1070_),
    .ZN(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2242_ (.A1(net26),
    .A2(_1066_),
    .B1(_1237_),
    .B2(_1160_),
    .ZN(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2243_ (.A1(_1145_),
    .A2(_1298_),
    .B1(_1300_),
    .B2(_1240_),
    .ZN(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2244_ (.A1(net28),
    .A2(_0892_),
    .ZN(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2245_ (.A1(net27),
    .A2(_0984_),
    .ZN(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _2246_ (.A1(_1298_),
    .A2(_1302_),
    .A3(_1303_),
    .ZN(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2247_ (.A1(_1301_),
    .A2(_1304_),
    .ZN(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2248_ (.A1(_1297_),
    .A2(_1305_),
    .Z(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2249_ (.A1(_1294_),
    .A2(_1306_),
    .ZN(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2250_ (.A1(_1292_),
    .A2(_1307_),
    .Z(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2251_ (.A1(_1280_),
    .A2(_1308_),
    .ZN(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2252_ (.A1(_1278_),
    .A2(_1309_),
    .Z(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2253_ (.A1(_1264_),
    .A2(_1311_),
    .ZN(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2254_ (.A1(_1262_),
    .A2(_1312_),
    .Z(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _2255_ (.A1(_1187_),
    .A2(_1258_),
    .A3(_1313_),
    .ZN(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2256_ (.A1(_1179_),
    .A2(_1251_),
    .ZN(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2257_ (.A1(_1179_),
    .A2(_1251_),
    .ZN(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _2258_ (.A1(_1093_),
    .A2(_1096_),
    .A3(_1315_),
    .B(_1316_),
    .ZN(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2259_ (.A1(_1314_),
    .A2(_1317_),
    .ZN(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2260_ (.A1(_1179_),
    .A2(_1251_),
    .Z(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2261_ (.A1(_1177_),
    .A2(_1319_),
    .Z(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2262_ (.A1(_1177_),
    .A2(_1319_),
    .ZN(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2263_ (.A1(_1089_),
    .A2(_1156_),
    .B(_1252_),
    .C(_1175_),
    .ZN(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__oai33_1 _2264_ (.A1(_1176_),
    .A2(_1320_),
    .A3(_1322_),
    .B1(_1323_),
    .B2(_1157_),
    .B3(_1161_),
    .ZN(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2265_ (.A1(_1157_),
    .A2(_1161_),
    .Z(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2266_ (.I(_1173_),
    .ZN(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2267_ (.A1(_1325_),
    .A2(_1326_),
    .A3(_1253_),
    .Z(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2268_ (.A1(_1324_),
    .A2(_1327_),
    .ZN(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2269_ (.A1(_1318_),
    .A2(_1328_),
    .Z(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2270_ (.I(_1329_),
    .Z(net43));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2271_ (.A1(_1258_),
    .A2(_1313_),
    .ZN(_1330_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2272_ (.A1(_1258_),
    .A2(_1313_),
    .ZN(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2273_ (.A1(_1187_),
    .A2(_1330_),
    .B(_1332_),
    .ZN(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2274_ (.A1(_1202_),
    .A2(_1261_),
    .ZN(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2275_ (.A1(_1264_),
    .A2(_1311_),
    .ZN(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2276_ (.A1(_1262_),
    .A2(_1312_),
    .B(_1335_),
    .ZN(_1336_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2277_ (.A1(_1268_),
    .A2(_1276_),
    .ZN(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2278_ (.A1(_1268_),
    .A2(_1276_),
    .ZN(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2279_ (.A1(_1265_),
    .A2(_1337_),
    .B(_1338_),
    .ZN(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2280_ (.A1(_1280_),
    .A2(_1308_),
    .ZN(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2281_ (.A1(_1278_),
    .A2(_1309_),
    .B(_1340_),
    .ZN(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2282_ (.I(_1275_),
    .ZN(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2283_ (.A1(_1270_),
    .A2(_1343_),
    .ZN(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2284_ (.A1(_1270_),
    .A2(_1343_),
    .ZN(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2285_ (.A1(_1201_),
    .A2(_1344_),
    .B(_1345_),
    .ZN(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2286_ (.I(_1282_),
    .ZN(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2287_ (.A1(_1285_),
    .A2(_1290_),
    .ZN(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2288_ (.A1(_1347_),
    .A2(_1291_),
    .B(_1348_),
    .ZN(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2289_ (.A1(_0535_),
    .A2(_0905_),
    .ZN(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2290_ (.A1(_0471_),
    .A2(_0944_),
    .ZN(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2291_ (.A1(_0225_),
    .A2(net23),
    .Z(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _2292_ (.A1(_1350_),
    .A2(_1351_),
    .A3(_1352_),
    .ZN(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2293_ (.A1(_1271_),
    .A2(_1274_),
    .ZN(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2294_ (.A1(_1272_),
    .A2(_1355_),
    .ZN(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2295_ (.A1(_1354_),
    .A2(_1356_),
    .Z(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2296_ (.A1(_1349_),
    .A2(_1357_),
    .ZN(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2297_ (.A1(_1346_),
    .A2(_1358_),
    .Z(_1359_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2298_ (.A1(_1294_),
    .A2(_1306_),
    .ZN(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2299_ (.A1(_1292_),
    .A2(_1307_),
    .B(_1360_),
    .ZN(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2300_ (.A1(net16),
    .A2(net18),
    .ZN(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2301_ (.A1(_1226_),
    .A2(_1362_),
    .ZN(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2302_ (.A1(_1286_),
    .A2(_1289_),
    .ZN(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2303_ (.A1(_1363_),
    .A2(_1365_),
    .ZN(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2304_ (.A1(_0554_),
    .A2(_0847_),
    .ZN(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2305_ (.A1(_1283_),
    .A2(_1296_),
    .Z(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2306_ (.A1(_1234_),
    .A2(_1367_),
    .B1(_1368_),
    .B2(_1295_),
    .ZN(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2307_ (.A1(_0567_),
    .A2(_0813_),
    .ZN(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2308_ (.A1(net15),
    .A2(net19),
    .ZN(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2309_ (.A1(_1362_),
    .A2(_1371_),
    .ZN(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2310_ (.A1(_1370_),
    .A2(_1372_),
    .Z(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2311_ (.A1(_1369_),
    .A2(_1373_),
    .ZN(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2312_ (.A1(_1366_),
    .A2(_1374_),
    .ZN(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2313_ (.A1(_1301_),
    .A2(_1304_),
    .ZN(_1377_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2314_ (.A1(_1297_),
    .A2(_1305_),
    .B(_1377_),
    .ZN(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2315_ (.A1(_0632_),
    .A2(_0723_),
    .ZN(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2316_ (.A1(_0584_),
    .A2(_0781_),
    .ZN(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2317_ (.A1(_1367_),
    .A2(_1379_),
    .A3(_1380_),
    .Z(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2318_ (.A1(_0095_),
    .A2(_1237_),
    .ZN(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2319_ (.I(_1066_),
    .Z(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2320_ (.I(_1237_),
    .Z(_1384_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2321_ (.A1(_0106_),
    .A2(_1383_),
    .B1(_1384_),
    .B2(_1299_),
    .ZN(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2322_ (.A1(_1241_),
    .A2(_1382_),
    .B1(_1385_),
    .B2(_1302_),
    .ZN(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2323_ (.A1(_0525_),
    .A2(_0893_),
    .ZN(_0001_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2324_ (.A1(_0364_),
    .A2(_1066_),
    .ZN(_0002_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _2325_ (.A1(_1382_),
    .A2(_0001_),
    .A3(_0002_),
    .ZN(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2326_ (.A1(_0000_),
    .A2(_0003_),
    .ZN(_0004_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2327_ (.A1(_1381_),
    .A2(_0004_),
    .Z(_0005_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _2328_ (.A1(_1376_),
    .A2(_1378_),
    .A3(_0005_),
    .ZN(_0006_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2329_ (.A1(_1361_),
    .A2(_0006_),
    .ZN(_0007_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2330_ (.A1(_1359_),
    .A2(_0007_),
    .Z(_0008_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2331_ (.A1(_1341_),
    .A2(_0008_),
    .Z(_0009_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2332_ (.A1(_1339_),
    .A2(_0009_),
    .Z(_0011_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _2333_ (.A1(_1334_),
    .A2(_1336_),
    .A3(_0011_),
    .ZN(_0012_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2334_ (.A1(_1333_),
    .A2(_0012_),
    .Z(_0013_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2335_ (.A1(_1314_),
    .A2(_1317_),
    .ZN(_0014_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2336_ (.A1(_1318_),
    .A2(_1328_),
    .B(_0014_),
    .ZN(_0015_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2337_ (.A1(_0013_),
    .A2(_0015_),
    .Z(_0016_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2338_ (.I(_0016_),
    .Z(net44));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2339_ (.A1(_1341_),
    .A2(_0008_),
    .ZN(_0017_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2340_ (.A1(_1339_),
    .A2(_0009_),
    .ZN(_0018_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2341_ (.A1(_0017_),
    .A2(_0018_),
    .ZN(_0019_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2342_ (.I(_1358_),
    .ZN(_0021_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2343_ (.A1(_1349_),
    .A2(_1357_),
    .Z(_0022_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2344_ (.A1(_1346_),
    .A2(_0021_),
    .B(_0022_),
    .ZN(_0023_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2345_ (.A1(_1361_),
    .A2(_0006_),
    .ZN(_0024_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2346_ (.A1(_1359_),
    .A2(_0007_),
    .B(_0024_),
    .ZN(_0025_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2347_ (.A1(_1354_),
    .A2(_1356_),
    .Z(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2348_ (.A1(_1369_),
    .A2(_1373_),
    .ZN(_0027_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2349_ (.A1(_1366_),
    .A2(_1374_),
    .B(_0027_),
    .ZN(_0028_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2350_ (.A1(_0598_),
    .A2(_0944_),
    .B1(_1009_),
    .B2(_0482_),
    .ZN(_0029_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2351_ (.A1(_0482_),
    .A2(_0598_),
    .A3(_0944_),
    .A4(net23),
    .Z(_0030_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2352_ (.A1(_0029_),
    .A2(_0030_),
    .Z(_0032_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2353_ (.A1(_1350_),
    .A2(_1351_),
    .ZN(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2354_ (.A1(_1350_),
    .A2(_1351_),
    .ZN(_0034_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2355_ (.A1(_0033_),
    .A2(_1352_),
    .B(_0034_),
    .ZN(_0035_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2356_ (.A1(_0032_),
    .A2(_0035_),
    .Z(_0036_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2357_ (.A1(_0028_),
    .A2(_0036_),
    .ZN(_0037_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2358_ (.A1(_0026_),
    .A2(_0037_),
    .Z(_0038_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2359_ (.A1(_1378_),
    .A2(_0005_),
    .ZN(_0039_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2360_ (.A1(_1378_),
    .A2(_0005_),
    .ZN(_0040_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2361_ (.A1(_1376_),
    .A2(_0039_),
    .B(_0040_),
    .ZN(_0041_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2362_ (.A1(net16),
    .A2(net19),
    .ZN(_0043_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2363_ (.A1(_1287_),
    .A2(_0043_),
    .ZN(_0044_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2364_ (.A1(_1370_),
    .A2(_1372_),
    .ZN(_0045_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2365_ (.A1(_0044_),
    .A2(_0045_),
    .ZN(_0046_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2366_ (.A1(_0583_),
    .A2(_0847_),
    .ZN(_0047_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2367_ (.A1(_1367_),
    .A2(_1380_),
    .Z(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2368_ (.A1(_1296_),
    .A2(_0047_),
    .B1(_0048_),
    .B2(_1379_),
    .ZN(_0049_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2369_ (.A1(_0567_),
    .A2(_0905_),
    .ZN(_0050_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2370_ (.A1(net15),
    .A2(net20),
    .ZN(_0051_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2371_ (.A1(_0043_),
    .A2(_0051_),
    .ZN(_0052_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2372_ (.A1(_0050_),
    .A2(_0052_),
    .Z(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2373_ (.A1(_0049_),
    .A2(_0054_),
    .ZN(_0055_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2374_ (.A1(_0046_),
    .A2(_0055_),
    .ZN(_0056_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2375_ (.A1(_0000_),
    .A2(_0003_),
    .ZN(_0057_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2376_ (.A1(_1381_),
    .A2(_0004_),
    .B(_0057_),
    .ZN(_0058_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2377_ (.A1(net28),
    .A2(_1070_),
    .ZN(_0059_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2378_ (.A1(_0364_),
    .A2(_1066_),
    .B1(_1237_),
    .B2(_0095_),
    .ZN(_0060_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2379_ (.A1(_1303_),
    .A2(_0059_),
    .B1(_0060_),
    .B2(_0001_),
    .ZN(_0061_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2380_ (.A1(_0553_),
    .A2(_0892_),
    .ZN(_0062_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2381_ (.A1(net29),
    .A2(_0984_),
    .ZN(_0063_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _2382_ (.A1(_0059_),
    .A2(_0062_),
    .A3(_0063_),
    .ZN(_0064_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2383_ (.A1(_0061_),
    .A2(_0064_),
    .ZN(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2384_ (.A1(_0724_),
    .A2(_0692_),
    .ZN(_0066_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2385_ (.A1(net32),
    .A2(_0781_),
    .ZN(_0067_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2386_ (.A1(_0047_),
    .A2(_0067_),
    .ZN(_0068_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2387_ (.A1(_0066_),
    .A2(_0068_),
    .ZN(_0069_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2388_ (.A1(_0065_),
    .A2(_0069_),
    .Z(_0070_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _2389_ (.A1(_0056_),
    .A2(_0058_),
    .A3(_0070_),
    .ZN(_0071_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2390_ (.A1(_0041_),
    .A2(_0071_),
    .Z(_0072_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2391_ (.A1(_0038_),
    .A2(_0072_),
    .Z(_0073_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2392_ (.A1(_0025_),
    .A2(_0073_),
    .ZN(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2393_ (.A1(_0023_),
    .A2(_0075_),
    .Z(_0076_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2394_ (.A1(_0019_),
    .A2(_0076_),
    .Z(_0077_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2395_ (.A1(_1336_),
    .A2(_0011_),
    .ZN(_0078_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2396_ (.A1(_1336_),
    .A2(_0011_),
    .ZN(_0079_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2397_ (.A1(_1334_),
    .A2(_0078_),
    .B(_0079_),
    .ZN(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2398_ (.A1(_0077_),
    .A2(_0080_),
    .ZN(_0081_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2399_ (.A1(_1314_),
    .A2(_1317_),
    .Z(_0082_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _2400_ (.A1(_1325_),
    .A2(_1253_),
    .A3(_0082_),
    .A4(_0013_),
    .ZN(_0083_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2401_ (.A1(_1173_),
    .A2(_0083_),
    .ZN(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2402_ (.A1(_0082_),
    .A2(_1324_),
    .A3(_0013_),
    .ZN(_0086_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2403_ (.A1(_1333_),
    .A2(_0012_),
    .ZN(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2404_ (.A1(_1333_),
    .A2(_0012_),
    .B(_1314_),
    .C(_1317_),
    .ZN(_0088_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2405_ (.A1(_0087_),
    .A2(_0088_),
    .Z(_0089_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2406_ (.A1(_0086_),
    .A2(_0089_),
    .ZN(_0090_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2407_ (.A1(_0084_),
    .A2(_0090_),
    .ZN(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2408_ (.A1(_0081_),
    .A2(_0091_),
    .Z(_0092_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2409_ (.I(_0092_),
    .Z(net46));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2410_ (.A1(_0077_),
    .A2(_0080_),
    .Z(_0093_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2411_ (.A1(_0081_),
    .A2(_0091_),
    .ZN(_0094_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2412_ (.A1(_0093_),
    .A2(_0094_),
    .ZN(_0096_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2413_ (.A1(_0019_),
    .A2(_0076_),
    .Z(_0097_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2414_ (.A1(_0025_),
    .A2(_0073_),
    .ZN(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2415_ (.A1(_0023_),
    .A2(_0075_),
    .Z(_0099_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2416_ (.A1(_0028_),
    .A2(_0036_),
    .ZN(_0100_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2417_ (.A1(_0026_),
    .A2(_0037_),
    .B(_0100_),
    .ZN(_0101_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2418_ (.A1(_0041_),
    .A2(_0071_),
    .Z(_0102_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2419_ (.A1(_0038_),
    .A2(_0072_),
    .B(_0102_),
    .ZN(_0103_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2420_ (.A1(_0032_),
    .A2(_0035_),
    .Z(_0104_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2421_ (.A1(_0049_),
    .A2(_0054_),
    .ZN(_0105_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2422_ (.A1(_0046_),
    .A2(_0055_),
    .B(_0105_),
    .ZN(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2423_ (.A1(_0598_),
    .A2(_1009_),
    .A3(_1351_),
    .ZN(_0108_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2424_ (.A1(_0107_),
    .A2(_0108_),
    .Z(_0109_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2425_ (.A1(_0104_),
    .A2(_0109_),
    .Z(_0110_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2426_ (.A1(_0058_),
    .A2(_0070_),
    .ZN(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2427_ (.A1(_0058_),
    .A2(_0070_),
    .ZN(_0112_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2428_ (.A1(_0056_),
    .A2(_0111_),
    .B(_0112_),
    .ZN(_0113_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2429_ (.A1(_0061_),
    .A2(_0064_),
    .ZN(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2430_ (.A1(_0065_),
    .A2(_0069_),
    .B(_0114_),
    .ZN(_0115_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2431_ (.A1(net29),
    .A2(net7),
    .ZN(_0116_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2432_ (.A1(_0525_),
    .A2(_1066_),
    .B1(_1237_),
    .B2(_0364_),
    .ZN(_0118_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2433_ (.A1(_0002_),
    .A2(_0116_),
    .B1(_0118_),
    .B2(_0062_),
    .ZN(_0119_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2434_ (.A1(net31),
    .A2(_0892_),
    .ZN(_0120_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2435_ (.A1(_0553_),
    .A2(_0984_),
    .ZN(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _2436_ (.A1(_0116_),
    .A2(_0120_),
    .A3(_0121_),
    .ZN(_0122_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2437_ (.A1(_0119_),
    .A2(_0122_),
    .ZN(_0123_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2438_ (.A1(_0723_),
    .A2(_0746_),
    .ZN(_0124_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2439_ (.A1(net32),
    .A2(net4),
    .ZN(_0125_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2440_ (.A1(net18),
    .A2(net3),
    .ZN(_0126_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2441_ (.A1(_0125_),
    .A2(_0126_),
    .ZN(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2442_ (.A1(_0124_),
    .A2(_0127_),
    .ZN(_0129_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2443_ (.A1(_0123_),
    .A2(_0129_),
    .Z(_0130_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2444_ (.A1(_0115_),
    .A2(_0130_),
    .Z(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2445_ (.A1(net16),
    .A2(net20),
    .ZN(_0132_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2446_ (.A1(_1371_),
    .A2(_0132_),
    .ZN(_0133_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2447_ (.A1(_0050_),
    .A2(_0052_),
    .ZN(_0134_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2448_ (.A1(_0133_),
    .A2(_0134_),
    .ZN(_0135_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2449_ (.A1(_1380_),
    .A2(_0125_),
    .B1(_0068_),
    .B2(_0066_),
    .ZN(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2450_ (.A1(_0568_),
    .A2(net22),
    .ZN(_0137_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2451_ (.A1(net15),
    .A2(net21),
    .ZN(_0138_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2452_ (.A1(_0132_),
    .A2(_0138_),
    .ZN(_0140_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2453_ (.A1(_0137_),
    .A2(_0140_),
    .ZN(_0141_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2454_ (.A1(_0136_),
    .A2(_0141_),
    .Z(_0142_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2455_ (.A1(_0135_),
    .A2(_0142_),
    .Z(_0143_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2456_ (.A1(_0131_),
    .A2(_0143_),
    .Z(_0144_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2457_ (.A1(_0113_),
    .A2(_0144_),
    .Z(_0145_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2458_ (.A1(_0110_),
    .A2(_0145_),
    .ZN(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2459_ (.A1(_0103_),
    .A2(_0146_),
    .Z(_0147_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2460_ (.A1(_0101_),
    .A2(_0147_),
    .ZN(_0148_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2461_ (.A1(_0098_),
    .A2(_0099_),
    .B(_0148_),
    .ZN(_0149_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2462_ (.A1(_0098_),
    .A2(_0099_),
    .A3(_0148_),
    .Z(_0151_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2463_ (.A1(_0149_),
    .A2(_0151_),
    .ZN(_0152_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2464_ (.A1(_0097_),
    .A2(_0152_),
    .ZN(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2465_ (.A1(_0096_),
    .A2(_0153_),
    .Z(_0154_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2466_ (.I(_0154_),
    .Z(net47));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2467_ (.A1(_0598_),
    .A2(_1087_),
    .A3(_1351_),
    .A4(_0107_),
    .ZN(_0155_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2468_ (.A1(_0104_),
    .A2(_0109_),
    .B(_0155_),
    .ZN(_0156_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2469_ (.A1(_0113_),
    .A2(_0144_),
    .Z(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2470_ (.A1(_0110_),
    .A2(_0145_),
    .B(_0157_),
    .ZN(_0158_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2471_ (.I(_0141_),
    .ZN(_0159_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2472_ (.A1(_0136_),
    .A2(_0159_),
    .ZN(_0161_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2473_ (.A1(_0135_),
    .A2(_0142_),
    .B(_0161_),
    .ZN(_0162_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2474_ (.A1(_0030_),
    .A2(_0162_),
    .Z(_0163_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2475_ (.A1(_0115_),
    .A2(_0130_),
    .Z(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2476_ (.A1(_0131_),
    .A2(_0143_),
    .B(_0164_),
    .ZN(_0165_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2477_ (.A1(_0119_),
    .A2(_0122_),
    .ZN(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2478_ (.A1(_0123_),
    .A2(_0129_),
    .B(_0166_),
    .ZN(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2479_ (.A1(net30),
    .A2(net7),
    .ZN(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2480_ (.A1(_0553_),
    .A2(_0984_),
    .B1(_1070_),
    .B2(net29),
    .ZN(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2481_ (.A1(_0063_),
    .A2(_0168_),
    .B1(_0169_),
    .B2(_0120_),
    .ZN(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2482_ (.A1(net32),
    .A2(net5),
    .ZN(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2483_ (.A1(_0583_),
    .A2(net6),
    .ZN(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _2484_ (.A1(_0168_),
    .A2(_0172_),
    .A3(_0173_),
    .ZN(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2485_ (.A1(_0170_),
    .A2(_0174_),
    .ZN(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2486_ (.A1(net18),
    .A2(net4),
    .ZN(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2487_ (.A1(net2),
    .A2(net20),
    .ZN(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2488_ (.A1(_0781_),
    .A2(_0746_),
    .ZN(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2489_ (.A1(_0176_),
    .A2(_0177_),
    .A3(_0178_),
    .Z(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2490_ (.A1(_0175_),
    .A2(_0179_),
    .Z(_0180_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2491_ (.A1(_0167_),
    .A2(_0180_),
    .Z(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2492_ (.A1(_0132_),
    .A2(_0138_),
    .ZN(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2493_ (.A1(_0137_),
    .A2(_0140_),
    .ZN(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2494_ (.A1(_0183_),
    .A2(_0184_),
    .ZN(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2495_ (.A1(_0067_),
    .A2(_0176_),
    .B1(_0127_),
    .B2(_0124_),
    .ZN(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2496_ (.A1(net16),
    .A2(net21),
    .ZN(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2497_ (.A1(net15),
    .A2(net22),
    .ZN(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2498_ (.A1(_0187_),
    .A2(_0188_),
    .ZN(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2499_ (.A1(_0567_),
    .A2(net23),
    .ZN(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2500_ (.A1(_0189_),
    .A2(_0190_),
    .ZN(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2501_ (.A1(_0186_),
    .A2(_0191_),
    .Z(_0192_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2502_ (.A1(_0185_),
    .A2(_0192_),
    .Z(_0194_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2503_ (.A1(_0181_),
    .A2(_0194_),
    .Z(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2504_ (.A1(_0165_),
    .A2(_0195_),
    .ZN(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2505_ (.A1(_0163_),
    .A2(_0196_),
    .ZN(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2506_ (.A1(_0158_),
    .A2(_0197_),
    .Z(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2507_ (.A1(_0156_),
    .A2(_0198_),
    .ZN(_0199_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2508_ (.A1(_0103_),
    .A2(_0146_),
    .ZN(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2509_ (.A1(_0101_),
    .A2(_0147_),
    .B(_0200_),
    .ZN(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2510_ (.A1(_0199_),
    .A2(_0201_),
    .ZN(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2511_ (.A1(_0149_),
    .A2(_0202_),
    .ZN(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2512_ (.A1(_0097_),
    .A2(_0093_),
    .B(_0152_),
    .ZN(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2513_ (.A1(_0081_),
    .A2(_0091_),
    .A3(_0153_),
    .B(_0205_),
    .ZN(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2514_ (.A1(_0203_),
    .A2(_0206_),
    .Z(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2515_ (.I(_0207_),
    .Z(net48));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2516_ (.A1(_0098_),
    .A2(_0099_),
    .B(_0148_),
    .C(_0202_),
    .ZN(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2517_ (.A1(_0203_),
    .A2(_0206_),
    .B(_0208_),
    .ZN(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2518_ (.A1(_0199_),
    .A2(_0201_),
    .ZN(_0210_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2519_ (.A1(_0030_),
    .A2(_0162_),
    .ZN(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2520_ (.I(_0165_),
    .ZN(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2521_ (.A1(_0212_),
    .A2(_0195_),
    .ZN(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2522_ (.A1(_0163_),
    .A2(_0196_),
    .ZN(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2523_ (.A1(_0213_),
    .A2(_0215_),
    .ZN(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2524_ (.I(_0191_),
    .ZN(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2525_ (.A1(_0186_),
    .A2(_0217_),
    .ZN(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2526_ (.A1(_0185_),
    .A2(_0192_),
    .B(_0218_),
    .ZN(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2527_ (.A1(_0167_),
    .A2(_0180_),
    .ZN(_0220_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2528_ (.A1(_0181_),
    .A2(_0194_),
    .ZN(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2529_ (.A1(_0220_),
    .A2(_0221_),
    .ZN(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2530_ (.A1(_0170_),
    .A2(_0174_),
    .ZN(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2531_ (.A1(_0175_),
    .A2(_0179_),
    .B(_0223_),
    .ZN(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2532_ (.A1(_0583_),
    .A2(_1070_),
    .ZN(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2533_ (.A1(_0168_),
    .A2(_0173_),
    .Z(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2534_ (.A1(_0121_),
    .A2(_0226_),
    .B1(_0227_),
    .B2(_0172_),
    .ZN(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2535_ (.A1(net18),
    .A2(_0892_),
    .ZN(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2536_ (.A1(_0632_),
    .A2(_1066_),
    .ZN(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _2537_ (.A1(_0226_),
    .A2(_0229_),
    .A3(_0230_),
    .ZN(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2538_ (.A1(_0228_),
    .A2(_0231_),
    .ZN(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2539_ (.A1(_0747_),
    .A2(_0848_),
    .ZN(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2540_ (.A1(_0724_),
    .A2(_0905_),
    .ZN(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2541_ (.A1(_0782_),
    .A2(_0813_),
    .ZN(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2542_ (.A1(_0233_),
    .A2(_0234_),
    .A3(_0235_),
    .Z(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2543_ (.A1(_0232_),
    .A2(_0237_),
    .Z(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2544_ (.A1(_0224_),
    .A2(_0238_),
    .ZN(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2545_ (.A1(_0719_),
    .A2(_0944_),
    .ZN(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2546_ (.A1(_0138_),
    .A2(_0240_),
    .B1(_0189_),
    .B2(_0190_),
    .ZN(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2547_ (.A1(_0176_),
    .A2(_0178_),
    .Z(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2548_ (.A1(_0126_),
    .A2(_0233_),
    .B1(_0242_),
    .B2(_0177_),
    .ZN(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2549_ (.A1(_0603_),
    .A2(net23),
    .ZN(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2550_ (.A1(_0240_),
    .A2(_0244_),
    .ZN(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2551_ (.A1(_0243_),
    .A2(_0245_),
    .Z(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2552_ (.A1(_0241_),
    .A2(_0246_),
    .Z(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2553_ (.A1(_0239_),
    .A2(_0248_),
    .Z(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2554_ (.A1(_0222_),
    .A2(_0249_),
    .Z(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2555_ (.A1(_0219_),
    .A2(_0250_),
    .Z(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _2556_ (.A1(_0211_),
    .A2(_0216_),
    .A3(_0251_),
    .ZN(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2557_ (.A1(_0158_),
    .A2(_0197_),
    .ZN(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2558_ (.A1(_0156_),
    .A2(_0198_),
    .B(_0253_),
    .ZN(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2559_ (.A1(_0252_),
    .A2(_0254_),
    .Z(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2560_ (.A1(_0210_),
    .A2(_0255_),
    .ZN(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2561_ (.A1(_0209_),
    .A2(_0256_),
    .ZN(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2562_ (.I(_0257_),
    .Z(net49));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2563_ (.A1(_0156_),
    .A2(_0198_),
    .Z(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2564_ (.A1(_0253_),
    .A2(_0259_),
    .B(_0252_),
    .ZN(_0260_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2565_ (.A1(_0222_),
    .A2(_0249_),
    .ZN(_0261_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2566_ (.A1(_0219_),
    .A2(_0250_),
    .ZN(_0262_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2567_ (.I(_0243_),
    .ZN(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2568_ (.I(_0246_),
    .ZN(_0264_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2569_ (.A1(_0241_),
    .A2(_0264_),
    .ZN(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2570_ (.A1(_0263_),
    .A2(_0245_),
    .B(_0265_),
    .ZN(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2571_ (.A1(_0224_),
    .A2(_0238_),
    .ZN(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2572_ (.A1(_0239_),
    .A2(_0248_),
    .B(_0267_),
    .ZN(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2573_ (.A1(_0228_),
    .A2(_0231_),
    .ZN(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2574_ (.A1(_0232_),
    .A2(_0237_),
    .B(_0270_),
    .ZN(_0271_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2575_ (.A1(_0632_),
    .A2(_1237_),
    .ZN(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2576_ (.A1(_0226_),
    .A2(_0230_),
    .Z(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2577_ (.A1(_0173_),
    .A2(_0272_),
    .B1(_0273_),
    .B2(_0229_),
    .ZN(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2578_ (.A1(_0747_),
    .A2(_0893_),
    .ZN(_0275_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2579_ (.A1(_0692_),
    .A2(_1383_),
    .ZN(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _2580_ (.A1(_0272_),
    .A2(_0275_),
    .A3(_0276_),
    .ZN(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2581_ (.A1(_0274_),
    .A2(_0277_),
    .ZN(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2582_ (.A1(_0848_),
    .A2(_0814_),
    .ZN(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2583_ (.A1(_0724_),
    .A2(_1199_),
    .ZN(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2584_ (.A1(_0782_),
    .A2(_0906_),
    .ZN(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2585_ (.A1(_0280_),
    .A2(_0281_),
    .A3(_0282_),
    .Z(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2586_ (.A1(_0278_),
    .A2(_0283_),
    .Z(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2587_ (.A1(_0271_),
    .A2(_0284_),
    .ZN(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2588_ (.A1(_0233_),
    .A2(_0235_),
    .Z(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2589_ (.A1(_0178_),
    .A2(_0280_),
    .B1(_0286_),
    .B2(_0234_),
    .ZN(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2590_ (.A1(_0719_),
    .A2(_1009_),
    .A3(_0188_),
    .ZN(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2591_ (.A1(_0287_),
    .A2(_0288_),
    .Z(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2592_ (.A1(_0285_),
    .A2(_0289_),
    .Z(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2593_ (.A1(_0269_),
    .A2(_0291_),
    .Z(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2594_ (.A1(_0266_),
    .A2(_0292_),
    .ZN(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2595_ (.A1(_0261_),
    .A2(_0262_),
    .B(_0293_),
    .ZN(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2596_ (.A1(_0261_),
    .A2(_0262_),
    .A3(_0293_),
    .Z(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2597_ (.A1(_0294_),
    .A2(_0295_),
    .ZN(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2598_ (.A1(_0216_),
    .A2(_0251_),
    .ZN(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2599_ (.A1(_0216_),
    .A2(_0251_),
    .ZN(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2600_ (.A1(_0211_),
    .A2(_0297_),
    .B(_0298_),
    .ZN(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2601_ (.A1(_0296_),
    .A2(_0299_),
    .Z(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2602_ (.A1(_0260_),
    .A2(_0300_),
    .Z(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2603_ (.A1(_0203_),
    .A2(_0256_),
    .ZN(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _2604_ (.A1(_0081_),
    .A2(_0153_),
    .A3(_0303_),
    .Z(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2605_ (.A1(_0086_),
    .A2(_0089_),
    .B(_0304_),
    .ZN(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _2606_ (.A1(_1169_),
    .A2(_1172_),
    .B(_0083_),
    .C(_0304_),
    .ZN(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2607_ (.A1(_0210_),
    .A2(_0208_),
    .ZN(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _2608_ (.A1(_0205_),
    .A2(_0303_),
    .B1(_0307_),
    .B2(_0255_),
    .ZN(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2609_ (.A1(_0305_),
    .A2(_0306_),
    .A3(_0308_),
    .ZN(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2610_ (.A1(_0302_),
    .A2(_0309_),
    .Z(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2611_ (.I(_0310_),
    .Z(net50));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2612_ (.I(_0260_),
    .ZN(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2613_ (.A1(_0312_),
    .A2(_0300_),
    .ZN(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2614_ (.I(_0302_),
    .ZN(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _2615_ (.A1(_0305_),
    .A2(_0306_),
    .A3(_0308_),
    .B(_0314_),
    .ZN(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2616_ (.I(_0188_),
    .ZN(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2617_ (.A1(_0316_),
    .A2(_0287_),
    .B(_0719_),
    .C(_1087_),
    .ZN(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2618_ (.I(_0317_),
    .ZN(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2619_ (.A1(_0271_),
    .A2(_0284_),
    .ZN(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2620_ (.A1(_0285_),
    .A2(_0289_),
    .B(_0319_),
    .ZN(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2621_ (.A1(_0848_),
    .A2(_0906_),
    .ZN(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2622_ (.A1(_0280_),
    .A2(_0282_),
    .Z(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2623_ (.A1(_0235_),
    .A2(_0321_),
    .B1(_0322_),
    .B2(_0281_),
    .ZN(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2624_ (.A1(_0274_),
    .A2(_0277_),
    .ZN(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2625_ (.A1(_0278_),
    .A2(_0283_),
    .B(_0324_),
    .ZN(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2626_ (.A1(_0692_),
    .A2(_1237_),
    .ZN(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2627_ (.A1(_0272_),
    .A2(_0276_),
    .Z(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2628_ (.A1(_0230_),
    .A2(_0326_),
    .B1(_0327_),
    .B2(_0275_),
    .ZN(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2629_ (.A1(_0813_),
    .A2(_0893_),
    .ZN(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2630_ (.A1(_0747_),
    .A2(_1383_),
    .ZN(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2631_ (.A1(_0326_),
    .A2(_0330_),
    .ZN(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2632_ (.A1(_0329_),
    .A2(_0331_),
    .Z(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2633_ (.A1(_0328_),
    .A2(_0333_),
    .ZN(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2634_ (.A1(_0724_),
    .A2(_1009_),
    .ZN(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2635_ (.A1(_0782_),
    .A2(_0944_),
    .ZN(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2636_ (.A1(_0321_),
    .A2(_0336_),
    .ZN(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2637_ (.A1(_0335_),
    .A2(_0337_),
    .ZN(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2638_ (.A1(_0334_),
    .A2(_0338_),
    .Z(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2639_ (.A1(_0325_),
    .A2(_0339_),
    .Z(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2640_ (.A1(_0323_),
    .A2(_0340_),
    .Z(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2641_ (.A1(_0320_),
    .A2(_0341_),
    .Z(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2642_ (.A1(_0318_),
    .A2(_0342_),
    .Z(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2643_ (.A1(_0269_),
    .A2(_0291_),
    .Z(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2644_ (.A1(_0266_),
    .A2(_0292_),
    .B(_0345_),
    .ZN(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2645_ (.A1(_0344_),
    .A2(_0346_),
    .ZN(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2646_ (.A1(_0296_),
    .A2(_0299_),
    .B(_0294_),
    .ZN(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2647_ (.A1(_0347_),
    .A2(_0348_),
    .ZN(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2648_ (.I(_0349_),
    .ZN(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2649_ (.A1(_0313_),
    .A2(_0315_),
    .B(_0350_),
    .ZN(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2650_ (.A1(_0313_),
    .A2(_0315_),
    .A3(_0350_),
    .Z(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2651_ (.A1(_0351_),
    .A2(_0352_),
    .ZN(net51));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2652_ (.A1(_0296_),
    .A2(_0299_),
    .A3(_0347_),
    .Z(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2653_ (.A1(_0354_),
    .A2(_0351_),
    .ZN(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2654_ (.A1(_0320_),
    .A2(_0341_),
    .ZN(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2655_ (.A1(_0318_),
    .A2(_0342_),
    .ZN(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2656_ (.A1(_0321_),
    .A2(_0336_),
    .ZN(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2657_ (.A1(_0335_),
    .A2(_0337_),
    .ZN(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2658_ (.A1(_0358_),
    .A2(_0359_),
    .ZN(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2659_ (.A1(_0328_),
    .A2(_0333_),
    .ZN(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2660_ (.A1(_0334_),
    .A2(_0338_),
    .B(_0361_),
    .ZN(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2661_ (.A1(_0848_),
    .A2(_1199_),
    .B1(_1009_),
    .B2(_0782_),
    .ZN(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2662_ (.A1(_0848_),
    .A2(_1009_),
    .ZN(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2663_ (.A1(_0336_),
    .A2(_0365_),
    .Z(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2664_ (.I(_0366_),
    .ZN(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2665_ (.A1(_0363_),
    .A2(_0367_),
    .ZN(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2666_ (.A1(_0747_),
    .A2(_1384_),
    .ZN(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2667_ (.A1(_0276_),
    .A2(_0369_),
    .B1(_0331_),
    .B2(_0329_),
    .ZN(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2668_ (.A1(_0893_),
    .A2(_0906_),
    .ZN(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2669_ (.A1(_0814_),
    .A2(_1384_),
    .ZN(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2670_ (.A1(_0330_),
    .A2(_0372_),
    .ZN(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2671_ (.A1(_0814_),
    .A2(_1383_),
    .B1(_1384_),
    .B2(_0747_),
    .ZN(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2672_ (.A1(_0373_),
    .A2(_0374_),
    .Z(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2673_ (.A1(_0371_),
    .A2(_0376_),
    .Z(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2674_ (.A1(_0370_),
    .A2(_0377_),
    .Z(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2675_ (.A1(_0368_),
    .A2(_0378_),
    .Z(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2676_ (.A1(_0362_),
    .A2(_0379_),
    .Z(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2677_ (.I(_0380_),
    .ZN(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2678_ (.A1(_0360_),
    .A2(_0381_),
    .Z(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2679_ (.A1(_0325_),
    .A2(_0339_),
    .ZN(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2680_ (.A1(_0323_),
    .A2(_0340_),
    .ZN(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2681_ (.A1(_0383_),
    .A2(_0384_),
    .ZN(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2682_ (.A1(_0382_),
    .A2(_0385_),
    .ZN(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2683_ (.A1(_0356_),
    .A2(_0357_),
    .B(_0387_),
    .ZN(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2684_ (.A1(_0356_),
    .A2(_0357_),
    .A3(_0387_),
    .Z(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2685_ (.A1(_0388_),
    .A2(_0389_),
    .ZN(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2686_ (.I(_0344_),
    .ZN(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2687_ (.A1(_0391_),
    .A2(_0346_),
    .ZN(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2688_ (.A1(_0294_),
    .A2(_0347_),
    .Z(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2689_ (.A1(_0392_),
    .A2(_0393_),
    .ZN(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2690_ (.A1(_0390_),
    .A2(_0394_),
    .Z(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2691_ (.A1(_0355_),
    .A2(_0395_),
    .Z(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2692_ (.I(_0396_),
    .Z(net52));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2693_ (.A1(_0370_),
    .A2(_0377_),
    .ZN(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2694_ (.A1(_0368_),
    .A2(_0378_),
    .ZN(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2695_ (.A1(_0398_),
    .A2(_0399_),
    .ZN(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2696_ (.A1(_0371_),
    .A2(_0376_),
    .ZN(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2697_ (.A1(_0373_),
    .A2(_0401_),
    .ZN(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2698_ (.A1(_0893_),
    .A2(_1199_),
    .ZN(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2699_ (.A1(_0906_),
    .A2(_1383_),
    .ZN(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2700_ (.A1(_0372_),
    .A2(_0404_),
    .ZN(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2701_ (.A1(_0403_),
    .A2(_0405_),
    .ZN(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2702_ (.A1(_0402_),
    .A2(_0406_),
    .Z(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2703_ (.A1(_0365_),
    .A2(_0408_),
    .Z(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2704_ (.A1(_0400_),
    .A2(_0409_),
    .Z(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2705_ (.A1(_0366_),
    .A2(_0410_),
    .Z(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2706_ (.A1(_0362_),
    .A2(_0379_),
    .ZN(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2707_ (.A1(_0360_),
    .A2(_0381_),
    .B(_0412_),
    .ZN(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2708_ (.A1(_0411_),
    .A2(_0413_),
    .Z(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2709_ (.A1(_0382_),
    .A2(_0385_),
    .Z(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2710_ (.A1(_0415_),
    .A2(_0388_),
    .ZN(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2711_ (.A1(_0414_),
    .A2(_0416_),
    .ZN(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2712_ (.A1(_0392_),
    .A2(_0390_),
    .B(_0417_),
    .ZN(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2713_ (.A1(_0392_),
    .A2(_0390_),
    .A3(_0417_),
    .Z(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2714_ (.A1(_0419_),
    .A2(_0420_),
    .ZN(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2715_ (.I(_0395_),
    .ZN(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2716_ (.A1(_0354_),
    .A2(_0351_),
    .B(_0422_),
    .ZN(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2717_ (.A1(_0393_),
    .A2(_0390_),
    .ZN(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2718_ (.A1(_0423_),
    .A2(_0424_),
    .ZN(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2719_ (.A1(_0421_),
    .A2(_0425_),
    .Z(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2720_ (.I(_0426_),
    .Z(net53));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2721_ (.A1(_0388_),
    .A2(_0414_),
    .ZN(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2722_ (.I(_0409_),
    .ZN(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2723_ (.A1(_0400_),
    .A2(_0429_),
    .ZN(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2724_ (.A1(_0366_),
    .A2(_0410_),
    .Z(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2725_ (.A1(_0906_),
    .A2(_1384_),
    .ZN(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2726_ (.A1(_1383_),
    .A2(_1199_),
    .ZN(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2727_ (.A1(_0893_),
    .A2(_1087_),
    .ZN(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2728_ (.A1(_0432_),
    .A2(_0433_),
    .A3(_0434_),
    .Z(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2729_ (.A1(_0372_),
    .A2(_0404_),
    .ZN(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2730_ (.A1(_0403_),
    .A2(_0405_),
    .ZN(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2731_ (.A1(_0436_),
    .A2(_0437_),
    .ZN(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2732_ (.A1(_0435_),
    .A2(_0438_),
    .Z(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2733_ (.A1(_0435_),
    .A2(_0438_),
    .ZN(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2734_ (.A1(_0440_),
    .A2(_0441_),
    .ZN(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2735_ (.A1(_0848_),
    .A2(_1087_),
    .A3(_0408_),
    .ZN(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2736_ (.A1(_0402_),
    .A2(_0406_),
    .B(_0443_),
    .ZN(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2737_ (.A1(_0442_),
    .A2(_0444_),
    .Z(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2738_ (.A1(_0430_),
    .A2(_0431_),
    .B(_0445_),
    .ZN(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2739_ (.I(_0446_),
    .ZN(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2740_ (.A1(_0430_),
    .A2(_0431_),
    .A3(_0445_),
    .ZN(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2741_ (.A1(_0447_),
    .A2(_0448_),
    .ZN(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2742_ (.A1(_0411_),
    .A2(_0413_),
    .ZN(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2743_ (.A1(_0415_),
    .A2(_0414_),
    .ZN(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2744_ (.A1(_0451_),
    .A2(_0452_),
    .ZN(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2745_ (.A1(_0449_),
    .A2(_0453_),
    .Z(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2746_ (.A1(_0427_),
    .A2(_0454_),
    .Z(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2747_ (.A1(_0422_),
    .A2(_0417_),
    .Z(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2748_ (.A1(_0349_),
    .A2(_0456_),
    .ZN(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2749_ (.A1(_0419_),
    .A2(_0424_),
    .ZN(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2750_ (.A1(_0420_),
    .A2(_0458_),
    .ZN(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2751_ (.A1(_0312_),
    .A2(_0300_),
    .A3(_0349_),
    .Z(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2752_ (.A1(_0354_),
    .A2(_0460_),
    .B(_0456_),
    .ZN(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _2753_ (.A1(_0315_),
    .A2(_0457_),
    .B(_0459_),
    .C(_0462_),
    .ZN(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2754_ (.A1(_0455_),
    .A2(_0463_),
    .Z(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2755_ (.I(_0464_),
    .Z(net54));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2756_ (.A1(_0452_),
    .A2(_0449_),
    .ZN(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2757_ (.I(_0442_),
    .ZN(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2758_ (.A1(_0466_),
    .A2(_0444_),
    .ZN(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2759_ (.A1(_0440_),
    .A2(_0467_),
    .ZN(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2760_ (.A1(_1199_),
    .A2(_1384_),
    .ZN(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2761_ (.A1(_0432_),
    .A2(_0433_),
    .Z(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2762_ (.A1(_0404_),
    .A2(_0469_),
    .B1(_0434_),
    .B2(_0470_),
    .ZN(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2763_ (.A1(_1383_),
    .A2(_1087_),
    .ZN(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2764_ (.A1(_0469_),
    .A2(_0473_),
    .Z(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2765_ (.A1(_0472_),
    .A2(_0474_),
    .ZN(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2766_ (.A1(_0468_),
    .A2(_0475_),
    .ZN(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2767_ (.I(_0476_),
    .ZN(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2768_ (.A1(_0451_),
    .A2(_0449_),
    .Z(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2769_ (.A1(_0447_),
    .A2(_0478_),
    .ZN(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2770_ (.A1(_0477_),
    .A2(_0479_),
    .Z(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2771_ (.I(_0480_),
    .ZN(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2772_ (.A1(_0427_),
    .A2(_0454_),
    .Z(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2773_ (.A1(_0455_),
    .A2(_0463_),
    .ZN(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2774_ (.A1(_0483_),
    .A2(_0484_),
    .ZN(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2775_ (.A1(_0465_),
    .A2(_0481_),
    .A3(_0485_),
    .Z(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2776_ (.I(_0486_),
    .Z(net55));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2777_ (.A1(_0477_),
    .A2(_0478_),
    .ZN(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2778_ (.A1(_0467_),
    .A2(_0475_),
    .ZN(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2779_ (.A1(_1384_),
    .A2(_1087_),
    .A3(_0433_),
    .ZN(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2780_ (.A1(_0472_),
    .A2(_0474_),
    .ZN(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2781_ (.A1(_0440_),
    .A2(_0475_),
    .B(_0490_),
    .ZN(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2782_ (.A1(_0489_),
    .A2(_0491_),
    .Z(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2783_ (.A1(_0488_),
    .A2(_0493_),
    .ZN(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2784_ (.A1(_0446_),
    .A2(_0476_),
    .A3(_0494_),
    .Z(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2785_ (.A1(_0446_),
    .A2(_0476_),
    .B(_0494_),
    .ZN(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2786_ (.A1(_0495_),
    .A2(_0496_),
    .Z(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2787_ (.A1(_0487_),
    .A2(_0497_),
    .Z(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2788_ (.I(_0483_),
    .ZN(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2789_ (.A1(_0465_),
    .A2(_0481_),
    .B(_0499_),
    .ZN(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2790_ (.A1(_0465_),
    .A2(_0481_),
    .ZN(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2791_ (.A1(_0484_),
    .A2(_0500_),
    .B(_0501_),
    .ZN(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2792_ (.A1(_0498_),
    .A2(_0502_),
    .ZN(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2793_ (.I(_0504_),
    .Z(net57));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2794_ (.A1(_0477_),
    .A2(_0478_),
    .A3(_0497_),
    .ZN(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2795_ (.A1(_0484_),
    .A2(_0500_),
    .B(_0498_),
    .C(_0501_),
    .ZN(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2796_ (.A1(_1383_),
    .A2(_1199_),
    .B(_0491_),
    .ZN(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2797_ (.A1(_1384_),
    .A2(_1087_),
    .ZN(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2798_ (.A1(_0467_),
    .A2(_0475_),
    .A3(_0493_),
    .B1(_0507_),
    .B2(_0508_),
    .ZN(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _2799_ (.A1(_0495_),
    .A2(_0505_),
    .A3(_0506_),
    .A4(_0509_),
    .Z(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2800_ (.I(_0510_),
    .Z(net58));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2801_ (.A1(_0624_),
    .A2(_0627_),
    .Z(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2802_ (.I(_0511_),
    .Z(net63));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2803_ (.I(_1246_),
    .ZN(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2804_ (.A1(_1062_),
    .A2(_1138_),
    .B1(_1192_),
    .B2(_1116_),
    .ZN(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2805_ (.A1(_0513_),
    .A2(_0514_),
    .ZN(net45));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2806_ (.D(net33),
    .CLK(clk),
    .Q(net66));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2807_ (.I(net34),
    .Z(net67));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2808_ (.I(net45),
    .Z(net74));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2809_ (.I(net56),
    .Z(net75));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2810_ (.I(net59),
    .Z(net76));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2811_ (.I(net60),
    .Z(net77));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2812_ (.I(net61),
    .Z(net78));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2813_ (.I(net62),
    .Z(net79));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2814_ (.I(net63),
    .Z(net80));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2815_ (.I(net64),
    .Z(net81));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2816_ (.I(net65),
    .Z(net82));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2817_ (.I(net35),
    .Z(net68));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2818_ (.I(net36),
    .Z(net69));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2819_ (.I(net37),
    .Z(net70));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2820_ (.I(net38),
    .Z(net71));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2821_ (.I(net39),
    .Z(net72));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2822_ (.I(net40),
    .Z(net73));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2823_ (.I(net41),
    .Z(net83));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2824_ (.I(net42),
    .Z(net90));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2825_ (.I(net43),
    .Z(net91));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2826_ (.I(net44),
    .Z(net92));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2827_ (.I(net46),
    .Z(net93));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2828_ (.I(net47),
    .Z(net94));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2829_ (.I(net48),
    .Z(net95));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2830_ (.I(net49),
    .Z(net96));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2831_ (.I(net50),
    .Z(net97));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2832_ (.I(net51),
    .Z(net98));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2833_ (.I(net52),
    .Z(net84));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2834_ (.I(net53),
    .Z(net85));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2835_ (.I(net54),
    .Z(net86));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2836_ (.I(net55),
    .Z(net87));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2837_ (.I(net57),
    .Z(net88));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2838_ (.I(net58),
    .Z(net89));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_85 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_86 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_87 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_88 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_89 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_90 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_91 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_92 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_93 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_94 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_95 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_96 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_97 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_98 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_99 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_512 ();
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input1 (.I(dba[0]),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input2 (.I(dba[10]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input3 (.I(dba[11]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input4 (.I(dba[12]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input5 (.I(dba[13]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input6 (.I(dba[14]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_1 input7 (.I(dba[15]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input8 (.I(dba[1]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input9 (.I(dba[2]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input10 (.I(dba[3]),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input11 (.I(dba[4]),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input12 (.I(dba[5]),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input13 (.I(dba[6]),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input14 (.I(dba[7]),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input15 (.I(dba[8]),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input16 (.I(dba[9]),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input17 (.I(dbb[0]),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input18 (.I(dbb[10]),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input19 (.I(dbb[11]),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input20 (.I(dbb[12]),
    .Z(net20));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input21 (.I(dbb[13]),
    .Z(net21));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input22 (.I(dbb[14]),
    .Z(net22));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input23 (.I(dbb[15]),
    .Z(net23));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input24 (.I(dbb[1]),
    .Z(net24));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input25 (.I(dbb[2]),
    .Z(net25));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input26 (.I(dbb[3]),
    .Z(net26));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input27 (.I(dbb[4]),
    .Z(net27));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input28 (.I(dbb[5]),
    .Z(net28));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input29 (.I(dbb[6]),
    .Z(net29));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input30 (.I(dbb[7]),
    .Z(net30));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input31 (.I(dbb[8]),
    .Z(net31));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input32 (.I(dbb[9]),
    .Z(net32));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input33 (.I(enable),
    .Z(net33));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output34 (.I(net34),
    .Z(Y[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output35 (.I(net35),
    .Z(Y[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output36 (.I(net36),
    .Z(Y[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output37 (.I(net37),
    .Z(Y[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output38 (.I(net38),
    .Z(Y[13]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output39 (.I(net39),
    .Z(Y[14]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output40 (.I(net40),
    .Z(Y[15]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output41 (.I(net41),
    .Z(Y[16]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output42 (.I(net42),
    .Z(Y[17]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output43 (.I(net43),
    .Z(Y[18]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output44 (.I(net44),
    .Z(Y[19]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output45 (.I(net45),
    .Z(Y[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output46 (.I(net46),
    .Z(Y[20]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output47 (.I(net47),
    .Z(Y[21]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output48 (.I(net48),
    .Z(Y[22]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output49 (.I(net49),
    .Z(Y[23]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output50 (.I(net50),
    .Z(Y[24]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output51 (.I(net51),
    .Z(Y[25]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output52 (.I(net52),
    .Z(Y[26]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output53 (.I(net53),
    .Z(Y[27]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output54 (.I(net54),
    .Z(Y[28]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output55 (.I(net55),
    .Z(Y[29]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output56 (.I(net56),
    .Z(Y[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output57 (.I(net57),
    .Z(Y[30]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output58 (.I(net58),
    .Z(Y[31]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output59 (.I(net59),
    .Z(Y[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output60 (.I(net60),
    .Z(Y[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output61 (.I(net61),
    .Z(Y[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output62 (.I(net62),
    .Z(Y[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output63 (.I(net63),
    .Z(Y[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output64 (.I(net64),
    .Z(Y[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output65 (.I(net65),
    .Z(Y[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output66 (.I(net66),
    .Z(done));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output67 (.I(net67),
    .Z(yA[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output68 (.I(net68),
    .Z(yA[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output69 (.I(net69),
    .Z(yA[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output70 (.I(net70),
    .Z(yA[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output71 (.I(net71),
    .Z(yA[13]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output72 (.I(net72),
    .Z(yA[14]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output73 (.I(net73),
    .Z(yA[15]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output74 (.I(net74),
    .Z(yA[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output75 (.I(net75),
    .Z(yA[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output76 (.I(net76),
    .Z(yA[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output77 (.I(net77),
    .Z(yA[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output78 (.I(net78),
    .Z(yA[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output79 (.I(net79),
    .Z(yA[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output80 (.I(net80),
    .Z(yA[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output81 (.I(net81),
    .Z(yA[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output82 (.I(net82),
    .Z(yA[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output83 (.I(net83),
    .Z(yB[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output84 (.I(net84),
    .Z(yB[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output85 (.I(net85),
    .Z(yB[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output86 (.I(net86),
    .Z(yB[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output87 (.I(net87),
    .Z(yB[13]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output88 (.I(net88),
    .Z(yB[14]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output89 (.I(net89),
    .Z(yB[15]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output90 (.I(net90),
    .Z(yB[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output91 (.I(net91),
    .Z(yB[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output92 (.I(net92),
    .Z(yB[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output93 (.I(net93),
    .Z(yB[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output94 (.I(net94),
    .Z(yB[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output95 (.I(net95),
    .Z(yB[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output96 (.I(net96),
    .Z(yB[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output97 (.I(net97),
    .Z(yB[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output98 (.I(net98),
    .Z(yB[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2416__A1 (.I(_0028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2357__A1 (.I(_0028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2519__A1 (.I(_0030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2474__A1 (.I(_0030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2352__A2 (.I(_0030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2418__A1 (.I(_0041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2390__A1 (.I(_0041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2371__A1 (.I(_0043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2363__A2 (.I(_0043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2386__A1 (.I(_0047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2368__A2 (.I(_0047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2421__A1 (.I(_0049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2373__A1 (.I(_0049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2495__A1 (.I(_0067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2386__A2 (.I(_0067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2513__A2 (.I(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2411__A2 (.I(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2408__A2 (.I(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2378__B2 (.I(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2318__A1 (.I(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1838__A1 (.I(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1837__A1 (.I(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1663__A1 (.I(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1601__A1 (.I(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1550__A2 (.I(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1431__I (.I(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2321__A1 (.I(_0106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1791__A1 (.I(_0106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1723__A1 (.I(_0106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1531__B1 (.I(_0106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1530__A4 (.I(_0106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1479__A2 (.I(_0106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1434__A2 (.I(_0106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1432__A2 (.I(_0106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2467__A4 (.I(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2424__A1 (.I(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2475__A1 (.I(_0115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2444__A1 (.I(_0115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2477__A1 (.I(_0119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2437__A1 (.I(_0119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2534__A1 (.I(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2436__A3 (.I(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2477__A2 (.I(_0122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2437__A2 (.I(_0122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2472__A1 (.I(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2454__A1 (.I(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2469__A2 (.I(_0144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2457__A2 (.I(_0144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2533__A1 (.I(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2484__A1 (.I(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2481__A2 (.I(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2530__A1 (.I(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2485__A1 (.I(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2577__A1 (.I(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2533__A2 (.I(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2484__A3 (.I(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2589__A1 (.I(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2547__A2 (.I(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2489__A3 (.I(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2616__I (.I(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2590__A3 (.I(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2498__A2 (.I(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1453__A1 (.I(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1452__A1 (.I(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1445__A1 (.I(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2155__A1 (.I(_0214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2070__A1 (.I(_0214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1914__A1 (.I(_0214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1612__A1 (.I(_0214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1550__A1 (.I(_0214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1490__A2 (.I(_0214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1461__A2 (.I(_0214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1442__I (.I(_0214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2566__A1 (.I(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2555__A1 (.I(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2565__A1 (.I(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2554__A1 (.I(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2571__A1 (.I(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2544__A1 (.I(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2291__A1 (.I(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2216__A1 (.I(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1600__A2 (.I(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1531__A2 (.I(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1530__A3 (.I(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1488__A2 (.I(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1462__B1 (.I(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1443__A2 (.I(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2576__A1 (.I(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2537__A1 (.I(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2534__A2 (.I(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2573__A1 (.I(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2538__A1 (.I(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2577__B2 (.I(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2537__A2 (.I(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2628__A1 (.I(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2576__A2 (.I(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2537__A3 (.I(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2588__A1 (.I(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2548__A2 (.I(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2542__A1 (.I(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2567__I (.I(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2551__A1 (.I(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1453__A2 (.I(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1452__A2 (.I(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1445__A2 (.I(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2608__B2 (.I(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2560__A2 (.I(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2612__I (.I(_0260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2602__A1 (.I(_0260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2644__A1 (.I(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2594__A1 (.I(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2627__A1 (.I(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2580__A1 (.I(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2577__A2 (.I(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2624__A1 (.I(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2581__A1 (.I(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2688__A1 (.I(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2646__B (.I(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2597__A1 (.I(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2652__A2 (.I(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2646__A2 (.I(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2601__A2 (.I(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2751__A2 (.I(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2613__A2 (.I(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2602__A2 (.I(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2606__C (.I(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2605__B (.I(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2615__A1 (.I(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2609__A1 (.I(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2615__A2 (.I(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2609__A2 (.I(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2615__A3 (.I(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2609__A3 (.I(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2680__A1 (.I(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2640__A1 (.I(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2660__A1 (.I(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2638__A1 (.I(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2687__A2 (.I(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2645__A2 (.I(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2751__A3 (.I(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2748__A1 (.I(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2648__I (.I(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2432__B2 (.I(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2378__A1 (.I(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2324__A1 (.I(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2168__A1 (.I(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1940__A1 (.I(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1847__A1 (.I(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1801__A1 (.I(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1456__I (.I(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1734__A1 (.I(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1674__A2 (.I(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1612__A2 (.I(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1551__A2 (.I(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1529__A2 (.I(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1508__A2 (.I(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1497__A2 (.I(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1457__A2 (.I(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2721__A1 (.I(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2710__A2 (.I(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2685__A1 (.I(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2785__A1 (.I(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2784__A1 (.I(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2739__I (.I(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1485__A1 (.I(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1469__A1 (.I(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2290__A1 (.I(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1917__A1 (.I(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1789__A1 (.I(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1601__A2 (.I(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1552__A2 (.I(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1523__A2 (.I(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1487__A2 (.I(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1466__I (.I(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2351__A1 (.I(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2350__B2 (.I(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2218__B2 (.I(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2217__A1 (.I(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1674__A1 (.I(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1521__A2 (.I(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1488__B1 (.I(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1467__A2 (.I(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2795__A1 (.I(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2791__A1 (.I(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2774__A2 (.I(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1485__A2 (.I(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1469__A2 (.I(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1583__A1 (.I(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1579__A1 (.I(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1478__A1 (.I(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1475__A1 (.I(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1581__A1 (.I(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1505__A1 (.I(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1475__A2 (.I(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2432__A1 (.I(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2323__A1 (.I(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2015__A1 (.I(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1933__A1 (.I(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1727__A2 (.I(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1666__A2 (.I(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1543__A2 (.I(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1482__I (.I(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2227__A1 (.I(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2180__A1 (.I(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1841__A1 (.I(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1795__A2 (.I(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1606__A2 (.I(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1567__A2 (.I(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1512__A2 (.I(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1483__A2 (.I(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2289__A1 (.I(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2217__A2 (.I(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1795__A1 (.I(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1663__A2 (.I(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1558__A2 (.I(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1555__I (.I(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1521__B1 (.I(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1492__A2 (.I(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1569__A2 (.I(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1568__A2 (.I(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1500__A3 (.I(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1517__A1 (.I(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1516__A1 (.I(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2480__A1 (.I(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2435__A1 (.I(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2380__A1 (.I(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2009__A2 (.I(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1926__A2 (.I(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1719__A2 (.I(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1660__A2 (.I(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1511__I (.I(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2304__A1 (.I(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2239__A1 (.I(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2179__A1 (.I(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1834__A2 (.I(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1789__A2 (.I(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1604__A2 (.I(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1513__A2 (.I(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1512__B1 (.I(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1536__A1 (.I(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1535__A1 (.I(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1548__A1 (.I(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1528__A1 (.I(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2499__A1 (.I(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2369__A1 (.I(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2307__A1 (.I(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2230__A1 (.I(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2171__A1 (.I(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1841__A2 (.I(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1618__A2 (.I(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1525__I (.I(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2450__A1 (.I(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1801__A2 (.I(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1723__A2 (.I(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1675__A2 (.I(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1616__B1 (.I(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1556__B1 (.I(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1554__A2 (.I(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1526__A2 (.I(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1548__A2 (.I(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1528__A2 (.I(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1538__A3 (.I(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1532__A2 (.I(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2532__A1 (.I(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2483__A1 (.I(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2366__A1 (.I(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2165__A1 (.I(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2085__A2 (.I(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2014__A2 (.I(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1840__A2 (.I(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1541__I (.I(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2316__A1 (.I(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2238__A1 (.I(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1932__A2 (.I(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1794__A2 (.I(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1726__A2 (.I(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1668__A2 (.I(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1605__A2 (.I(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1542__A2 (.I(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1662__A1 (.I(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1597__A2 (.I(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1544__A2 (.I(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2467__A1 (.I(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2423__A1 (.I(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2351__A2 (.I(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2350__A1 (.I(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2218__A1 (.I(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2214__A1 (.I(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1734__A2 (.I(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1556__A2 (.I(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2231__A1 (.I(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2172__A1 (.I(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2085__A1 (.I(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2009__A1 (.I(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1933__A2 (.I(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1681__A2 (.I(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1615__A2 (.I(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1560__I (.I(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2549__A1 (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1847__A2 (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1838__A2 (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1791__A2 (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1735__A2 (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1679__A2 (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1616__A2 (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1561__A2 (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1595__A2 (.I(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1594__A2 (.I(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1565__A3 (.I(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1632__A1 (.I(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1631__A1 (.I(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1578__A1 (.I(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1582__A1 (.I(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1576__A1 (.I(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1574__A1 (.I(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1632__A2 (.I(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1631__A2 (.I(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1578__A2 (.I(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1640__A2 (.I(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1633__A2 (.I(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1578__A3 (.I(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2801__A2 (.I(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1585__A2 (.I(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1643__A3 (.I(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1593__A1 (.I(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2575__A1 (.I(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2536__A1 (.I(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2315__A1 (.I(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2001__A2 (.I(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1917__A2 (.I(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1878__A2 (.I(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1780__A2 (.I(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1591__I (.I(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1644__A1 (.I(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1625__A1 (.I(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1673__A1 (.I(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1623__A1 (.I(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2225__A1 (.I(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2165__A2 (.I(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2015__A2 (.I(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1940__A2 (.I(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1837__A2 (.I(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1678__I (.I(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1677__A2 (.I(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1620__A2 (.I(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1658__A2 (.I(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1657__A2 (.I(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1624__A3 (.I(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1645__A2 (.I(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1626__A2 (.I(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1693__A2 (.I(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1630__A2 (.I(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1699__A1 (.I(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1656__A1 (.I(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2231__A2 (.I(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2171__A2 (.I(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2067__A2 (.I(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1997__A2 (.I(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1913__A2 (.I(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1874__A2 (.I(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1709__A2 (.I(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1651__I (.I(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2626__A1 (.I(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2579__A1 (.I(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2384__A2 (.I(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1914__B1 (.I(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1875__B1 (.I(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1711__B1 (.I(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1653__A4 (.I(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1652__A2 (.I(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1700__A1 (.I(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1689__A1 (.I(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1667__A1 (.I(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1662__A2 (.I(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1718__A1 (.I(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1688__A1 (.I(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1733__A1 (.I(_0717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1687__A1 (.I(_0717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2617__B (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2590__A1 (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2545__A1 (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1838__B1 (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1802__A2 (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1740__A2 (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1738__A2 (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1679__B1 (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2438__A1 (.I(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2315__A2 (.I(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2238__A2 (.I(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2179__A2 (.I(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1929__A2 (.I(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1848__A2 (.I(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1807__A2 (.I(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1683__I (.I(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2634__A1 (.I(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2583__A1 (.I(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2540__A1 (.I(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2384__A1 (.I(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1805__A2 (.I(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1738__B1 (.I(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1737__A2 (.I(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1684__A2 (.I(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1700__A2 (.I(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1689__A2 (.I(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1754__A1 (.I(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1695__A1 (.I(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1767__A1 (.I(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1750__A1 (.I(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1768__A1 (.I(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1715__A1 (.I(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2488__A2 (.I(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2438__A2 (.I(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2153__A2 (.I(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2071__A2 (.I(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2000__A2 (.I(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1916__A2 (.I(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1779__A2 (.I(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1707__I (.I(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2671__B2 (.I(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2666__A1 (.I(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2630__A1 (.I(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2578__A1 (.I(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2539__A1 (.I(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2230__A2 (.I(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1877__A2 (.I(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1708__A2 (.I(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1769__A1 (.I(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1748__A1 (.I(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1728__A1 (.I(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1720__A2 (.I(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1788__A1 (.I(_0771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1747__A1 (.I(_0771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1800__A1 (.I(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1746__A1 (.I(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2488__A1 (.I(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2385__A2 (.I(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2316__A2 (.I(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2239__A2 (.I(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2092__A2 (.I(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1941__A2 (.I(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1804__A2 (.I(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1742__I (.I(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2661__B2 (.I(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2635__A1 (.I(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2584__A1 (.I(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2541__A1 (.I(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2180__A2 (.I(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1851__A2 (.I(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1805__B1 (.I(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1743__A2 (.I(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1769__A2 (.I(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1748__A2 (.I(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2122__A1 (.I(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1763__A1 (.I(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2122__A2 (.I(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1763__A2 (.I(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1889__A1 (.I(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1816__A1 (.I(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1824__A1 (.I(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1784__A1 (.I(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2629__A1 (.I(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2541__A2 (.I(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2307__A2 (.I(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2218__A2 (.I(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2217__A3 (.I(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2070__A2 (.I(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1994__A2 (.I(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1775__I (.I(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2671__A1 (.I(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2669__A1 (.I(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2582__A2 (.I(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2214__A2 (.I(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1870__A3 (.I(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1869__A2 (.I(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1862__A2 (.I(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1776__A2 (.I(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1828__A1 (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1827__A1 (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1815__A2 (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1832__A1 (.I(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1814__A1 (.I(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1846__A1 (.I(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1813__A1 (.I(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2366__A2 (.I(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2304__A2 (.I(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2227__A2 (.I(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2168__A2 (.I(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2022__A2 (.I(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1944__A2 (.I(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1850__A2 (.I(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1809__I (.I(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2735__A1 (.I(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2662__A1 (.I(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2661__A1 (.I(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2621__A1 (.I(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2582__A1 (.I(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2539__A2 (.I(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1851__B1 (.I(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1810__A2 (.I(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1828__A2 (.I(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1827__A2 (.I(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1815__A3 (.I(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1896__A1 (.I(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1885__A1 (.I(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1900__A1 (.I(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1861__A1 (.I(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1925__A1 (.I(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1860__A1 (.I(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2535__A2 (.I(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2434__A2 (.I(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2380__A2 (.I(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2244__A2 (.I(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2186__A2 (.I(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2026__A2 (.I(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1943__A2 (.I(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1855__I (.I(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2727__A1 (.I(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2698__A1 (.I(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2668__A1 (.I(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2629__A2 (.I(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2578__A2 (.I(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2323__A2 (.I(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1944__B1 (.I(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1856__A2 (.I(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2027__A1 (.I(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1857__A3 (.I(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1924__A2 (.I(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1923__A2 (.I(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1860__A3 (.I(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1900__A2 (.I(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1861__A2 (.I(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1898__A1 (.I(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1882__A1 (.I(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2540__A2 (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2369__A2 (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2289__A2 (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2217__A4 (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2155__A2 (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1994__B1 (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1909__A2 (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1868__I (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2725__A1 (.I(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2699__A1 (.I(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2668__A2 (.I(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2621__A2 (.I(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2584__A2 (.I(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2218__B1 (.I(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1870__A4 (.I(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1869__B1 (.I(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1975__A1 (.I(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1921__A1 (.I(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2635__A2 (.I(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2545__A2 (.I(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2351__A3 (.I(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2350__A2 (.I(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2290__A2 (.I(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2148__I (.I(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1991__A2 (.I(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1908__A2 (.I(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1983__A1 (.I(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1954__A1 (.I(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2008__A1 (.I(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1953__A1 (.I(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2480__A2 (.I(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2435__A2 (.I(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2381__A2 (.I(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2245__A2 (.I(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2187__A2 (.I(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2095__A2 (.I(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2025__I (.I(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1948__A2 (.I(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2096__A1 (.I(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1949__A3 (.I(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1983__A2 (.I(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1954__A2 (.I(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1984__A2 (.I(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1955__A2 (.I(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1971__A2 (.I(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1970__A2 (.I(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1956__A3 (.I(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2116__A1 (.I(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1966__A1 (.I(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1963__A1 (.I(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2118__A1 (.I(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2117__A1 (.I(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2110__I (.I(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2041__A1 (.I(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2662__A2 (.I(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2661__B1 (.I(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2634__A2 (.I(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2590__A2 (.I(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2423__A2 (.I(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2350__B1 (.I(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2045__I (.I(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1974__A2 (.I(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1994__B2 (.I(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1877__A1 (.I(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1875__B2 (.I(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1711__A1 (.I(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1668__A1 (.I(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1604__A1 (.I(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1479__A1 (.I(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1388__I (.I(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1984__B (.I(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2050__A1 (.I(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2005__A1 (.I(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2149__B2 (.I(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1873__A1 (.I(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1529__A1 (.I(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1458__A1 (.I(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1440__A1 (.I(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1438__A1 (.I(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1418__A1 (.I(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1392__A1 (.I(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1851__B2 (.I(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1743__A1 (.I(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1684__A1 (.I(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1620__A1 (.I(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1616__A1 (.I(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1526__A1 (.I(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1492__A1 (.I(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1390__I (.I(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2167__A1 (.I(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2079__A1 (.I(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2016__A1 (.I(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2010__A2 (.I(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2170__A1 (.I(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2082__A1 (.I(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2023__A1 (.I(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2013__A2 (.I(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1805__B2 (.I(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1679__B2 (.I(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1561__A1 (.I(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1521__B2 (.I(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1488__B2 (.I(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1467__A1 (.I(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1443__A1 (.I(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1391__I (.I(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2061__A1 (.I(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2017__A1 (.I(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2077__A1 (.I(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2035__A1 (.I(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2083__B2 (.I(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2023__A2 (.I(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2804__A1 (.I(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1738__B2 (.I(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1556__B2 (.I(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1462__B2 (.I(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1438__B2 (.I(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1422__A1 (.I(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1406__A1 (.I(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1392__A2 (.I(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2185__A1 (.I(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2031__A1 (.I(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2027__A2 (.I(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2536__A2 (.I(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2432__A2 (.I(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2378__A2 (.I(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2324__A2 (.I(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2319__I (.I(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2242__A2 (.I(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2184__A2 (.I(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2026__B1 (.I(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2096__B2 (.I(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2031__A2 (.I(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2532__A2 (.I(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2480__B1 (.I(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2377__A2 (.I(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2241__A2 (.I(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2183__I (.I(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2182__A2 (.I(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2095__B1 (.I(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2030__A2 (.I(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2056__A2 (.I(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2037__A2 (.I(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2111__A2 (.I(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2040__A2 (.I(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2184__B2 (.I(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2095__A1 (.I(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2026__A1 (.I(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1944__A1 (.I(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1943__A1 (.I(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1850__A1 (.I(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1615__A1 (.I(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1394__I (.I(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2797__A2 (.I(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2779__A2 (.I(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2763__A2 (.I(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2735__A2 (.I(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2727__A2 (.I(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2617__C (.I(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2467__A2 (.I(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2046__A2 (.I(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2258__A1 (.I(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2128__A1 (.I(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2054__A1 (.I(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1851__A1 (.I(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1804__A1 (.I(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1737__A1 (.I(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1677__A1 (.I(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1554__A1 (.I(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1520__A1 (.I(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1487__A1 (.I(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1395__I (.I(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2056__B (.I(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1805__A1 (.I(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1738__A1 (.I(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1679__A1 (.I(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1616__B2 (.I(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1521__A1 (.I(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1488__A1 (.I(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1461__A1 (.I(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1396__I (.I(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2132__A1 (.I(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2131__A1 (.I(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2075__A2 (.I(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2144__A1 (.I(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2074__A1 (.I(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2804__B2 (.I(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1556__A1 (.I(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1462__A1 (.I(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1438__A2 (.I(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1437__A1 (.I(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1418__A2 (.I(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1408__A1 (.I(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1399__A1 (.I(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2140__A1 (.I(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2104__A1 (.I(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2166__A1 (.I(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2086__A1 (.I(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2080__A2 (.I(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2169__A1 (.I(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2093__A1 (.I(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2083__A2 (.I(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2063__A1 (.I(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1991__A1 (.I(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1870__A1 (.I(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1869__A1 (.I(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1649__A1 (.I(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1497__A1 (.I(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1434__A1 (.I(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1398__I (.I(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2146__A2 (.I(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2087__A2 (.I(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2164__A1 (.I(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2103__A1 (.I(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2163__A1 (.I(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2102__A1 (.I(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2170__B2 (.I(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2093__A2 (.I(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2804__A2 (.I(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1653__A1 (.I(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1512__A1 (.I(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1508__A1 (.I(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1429__A1 (.I(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1419__A1 (.I(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1408__A2 (.I(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1399__A2 (.I(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2177__A2 (.I(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2100__A2 (.I(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2129__A2 (.I(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2106__A2 (.I(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2242__B2 (.I(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2184__A1 (.I(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1946__A1 (.I(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1853__A1 (.I(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1807__A1 (.I(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1618__A1 (.I(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1523__A1 (.I(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1401__I (.I(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1740__A1 (.I(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1681__A1 (.I(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1558__A1 (.I(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1490__A1 (.I(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1464__A1 (.I(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1440__A2 (.I(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1419__A2 (.I(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1404__A1 (.I(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1862__A1 (.I(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1776__A1 (.I(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1653__A2 (.I(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1652__A1 (.I(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1512__B2 (.I(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1432__A1 (.I(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1414__A1 (.I(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1403__I (.I(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2138__A1 (.I(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2137__A1 (.I(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2202__A1 (.I(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2195__A1 (.I(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2804__B1 (.I(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2046__A1 (.I(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1974__A1 (.I(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1643__A1 (.I(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1592__A1 (.I(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1567__A1 (.I(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1406__A2 (.I(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1404__A2 (.I(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2204__A1 (.I(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2161__A1 (.I(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2796__A2 (.I(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2760__A1 (.I(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2726__A2 (.I(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2698__A2 (.I(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2661__A2 (.I(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2583__A2 (.I(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2216__A2 (.I(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2149__A2 (.I(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2210__A1 (.I(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2159__A1 (.I(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2208__A1 (.I(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2193__A1 (.I(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2301__A1 (.I(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2173__A2 (.I(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2224__A1 (.I(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2192__A1 (.I(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2626__A2 (.I(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2575__A2 (.I(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2432__B1 (.I(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2378__B1 (.I(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2320__I (.I(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2318__A2 (.I(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2242__B1 (.I(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2184__B1 (.I(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2203__A2 (.I(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2196__A2 (.I(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2203__B (.I(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2274__A2 (.I(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2207__A2 (.I(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2278__A1 (.I(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2277__A1 (.I(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2222__A2 (.I(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2284__A1 (.I(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2283__A1 (.I(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2221__A2 (.I(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2280__A1 (.I(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2251__A1 (.I(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2286__I (.I(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2235__A1 (.I(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2363__A1 (.I(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2232__A2 (.I(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1848__A1 (.I(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1838__B2 (.I(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1802__A1 (.I(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1735__A1 (.I(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1675__A1 (.I(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1613__A1 (.I(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1552__A1 (.I(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1413__I (.I(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2368__A1 (.I(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2305__A2 (.I(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2240__A3 (.I(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2321__B2 (.I(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1600__A1 (.I(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1531__A1 (.I(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1530__A2 (.I(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1495__A2 (.I(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1458__A2 (.I(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1429__A2 (.I(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1414__A2 (.I(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2344__A1 (.I(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2297__A1 (.I(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2343__A1 (.I(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2296__A1 (.I(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2467__A3 (.I(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2423__A3 (.I(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2354__A2 (.I(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2353__A2 (.I(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2292__A2 (.I(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2309__A1 (.I(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2301__A2 (.I(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2349__A1 (.I(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2312__A1 (.I(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2367__A1 (.I(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2317__A1 (.I(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2306__A2 (.I(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2348__A1 (.I(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2311__A1 (.I(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2446__A1 (.I(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2309__A2 (.I(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1914__B2 (.I(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1780__A1 (.I(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1606__A1 (.I(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1551__A1 (.I(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1530__A1 (.I(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1495__A1 (.I(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1464__A2 (.I(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1421__I (.I(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2449__A1 (.I(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2367__A2 (.I(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2317__A3 (.I(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2796__A1 (.I(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2763__A1 (.I(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2726__A1 (.I(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2699__A2 (.I(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2671__A2 (.I(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2630__A2 (.I(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2579__A2 (.I(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2321__A2 (.I(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2797__A1 (.I(_1384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2779__A1 (.I(_1384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2760__A2 (.I(_1384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2725__A2 (.I(_1384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2671__B1 (.I(_1384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2669__A2 (.I(_1384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2666__A2 (.I(_1384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2321__B1 (.I(_1384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2322__B1 (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2150__A1 (.I(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2149__A1 (.I(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1875__A1 (.I(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1531__B2 (.I(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1462__A2 (.I(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1438__B1 (.I(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1437__A2 (.I(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1422__A2 (.I(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2806__CLK (.I(clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(dba[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(dba[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(dba[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(dba[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(dba[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(dba[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(dba[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(dba[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(dba[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(dba[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input11_I (.I(dba[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input12_I (.I(dba[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input13_I (.I(dba[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input14_I (.I(dba[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input15_I (.I(dba[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input16_I (.I(dba[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input17_I (.I(dbb[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input18_I (.I(dbb[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input19_I (.I(dbb[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input20_I (.I(dbb[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input21_I (.I(dbb[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input22_I (.I(dbb[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input23_I (.I(dbb[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input24_I (.I(dbb[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input25_I (.I(dbb[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input26_I (.I(dbb[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input27_I (.I(dbb[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input28_I (.I(dbb[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input29_I (.I(dbb[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input30_I (.I(dbb[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input31_I (.I(dbb[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input32_I (.I(dbb[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input33_I (.I(enable));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1908__A1 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1870__A2 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1869__B2 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1708__A1 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1542__A1 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1483__A1 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1457__A1 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1402__I (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2487__A1 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2091__A2 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2021__A2 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1682__I (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2440__A2 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2011__A2 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1853__A2 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1741__I (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2486__A2 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2439__A2 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2081__A2 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1946__A2 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1808__I (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2482__A2 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2097__A2 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2028__A2 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1854__I (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2483__A2 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2098__A2 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2024__A2 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1947__I (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2479__A2 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2431__A2 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2094__A2 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2029__I (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1909__A1 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1779__A1 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1711__B2 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1605__A1 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1513__A1 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1397__I (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2064__A1 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1910__A1 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1709__A1 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1543__A1 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1387__I (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1994__A1 (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1992__A1 (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1916__A1 (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1874__A1 (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1726__A1 (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1660__A1 (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1420__I (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2000__A1 (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1913__A1 (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1878__A1 (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1794__A1 (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1719__A1 (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1666__A1 (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1441__I (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2156__A1 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2071__A1 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1997__A1 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1840__A1 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1727__A1 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1465__I (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2153__A1 (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2067__A1 (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2001__A1 (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1932__A1 (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1834__A1 (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1613__A2 (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1520__A2 (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1491__I (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2084__A1 (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2014__A1 (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1926__A1 (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1524__I (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2497__A1 (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2451__A1 (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2370__A1 (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2308__A1 (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1559__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2496__A1 (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2445__A1 (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2362__A1 (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2300__A1 (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2078__A2 (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1619__I (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2095__B2 (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2030__A1 (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2026__B2 (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1948__A1 (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1944__B2 (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1856__A1 (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1810__A1 (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1389__I (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2535__A1 (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2486__A1 (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2440__A1 (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2300__A2 (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1650__I (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2487__A2 (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2445__A2 (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2370__A2 (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2156__A2 (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1910__A2 (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1774__I (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2496__A2 (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2451__A2 (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1992__A2 (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1867__I (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2497__A2 (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2450__A2 (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2064__A2 (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1907__I (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2549__A2 (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2499__A2 (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2351__A4 (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2291__A2 (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2150__A2 (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2149__B1 (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2063__A2 (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1973__I (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2182__A1 (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2098__A1 (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2028__A1 (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1400__I (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2242__A1 (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2241__A1 (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2187__A1 (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2097__A1 (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2022__A1 (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1941__A1 (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1412__I (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2245__A1 (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2186__A1 (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2081__A1 (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2011__A1 (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1929__A1 (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1430__I (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2377__A1 (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2244__A1 (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2092__A1 (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2021__A1 (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1455__I (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2482__A1 (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2439__A1 (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2385__A1 (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2225__A2 (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2172__A2 (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2084__A2 (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1590__I (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output34_I (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2807__I (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1408__A3 (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output35_I (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2817__I (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output36_I (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2818__I (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output37_I (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2819__I (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output38_I (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2820__I (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output39_I (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2821__I (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output40_I (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2822__I (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output41_I (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2823__I (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output42_I (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2824__I (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output43_I (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2825__I (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output44_I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2826__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output45_I (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2808__I (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output46_I (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2827__I (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output47_I (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2828__I (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output48_I (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2829__I (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output49_I (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2830__I (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output50_I (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2831__I (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output51_I (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2832__I (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output52_I (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2833__I (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output53_I (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2834__I (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output54_I (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2835__I (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output55_I (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2836__I (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output56_I (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2809__I (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output57_I (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2837__I (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output58_I (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2838__I (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output59_I (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2810__I (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output60_I (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2811__I (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output61_I (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2812__I (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output62_I (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2813__I (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output63_I (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2814__I (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output64_I (.I(net64));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2815__I (.I(net64));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output65_I (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2816__I (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output68_I (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output76_I (.I(net76));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output77_I (.I(net77));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output78_I (.I(net78));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output79_I (.I(net79));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output80_I (.I(net80));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output81_I (.I(net81));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output82_I (.I(net82));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output97_I (.I(net97));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_686 ();
endmodule

