* NGSPICE file created from DiffDigota.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyb_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyb_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VSS
.ends

.subckt DiffDigota INmb INpb OUTm OUTp cmnmos cmpmos oe omnmos ompmos opnmos oppmos
+ vdd vss
XFILLER_9_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput7 net7 cmpmos vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_6_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput10 net10 opnmos vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput8 net8 omnmos vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA_input3_I OUTm vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput9 net9 ompmos vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_11_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput11 net11 oppmos vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_3_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input1_I INmb vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09__A1 net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_5_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09_ net5 _00_ _01_ net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_4_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08_ net2 _01_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_5_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07_ net1 _00_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_5_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_2_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput1 INmb net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XPHY_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xinput2 INpb net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XPHY_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_4_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput3 OUTm net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_4_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput4 OUTp net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_1_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput5 oe net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__17__A1 net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__19__B net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input4_I OUTp vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input2_I INpb vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10__I net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_19_ _00_ _06_ net5 net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_5_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_18_ net4 net3 net2 _06_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_11_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_17_ net5 _00_ _05_ net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_5_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_16_ net4 net3 net2 _05_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_2_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15_ _02_ _01_ _04_ net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_5_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_14_ net4 net3 net1 _04_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_3_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13_ _01_ _03_ _02_ net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_6_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12_ net4 net3 net1 _03_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_3_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_7_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11_ _02_ _00_ _01_ net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_3_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_3_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10_ net5 _02_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_3_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input5_I oe vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput6 net6 cmnmos vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
.ends

