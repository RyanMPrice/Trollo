// This is the unpowered netlist.
module WavePWM (clk,
    enable,
    qcomplex,
    qcos,
    qsin,
    rst,
    divSel);
 input clk;
 input enable;
 output qcomplex;
 output qcos;
 output qsin;
 input rst;
 input [3:0] divSel;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire \csTable.address[0] ;
 wire \csTable.address[1] ;
 wire \csTable.address[2] ;
 wire \csTable.address[3] ;
 wire \csTable.address[4] ;
 wire \csTable.address[5] ;
 wire \csTable.address[6] ;
 wire \csTable.address[7] ;
 wire \freeRunCntr[0] ;
 wire \freeRunCntr[10] ;
 wire \freeRunCntr[11] ;
 wire \freeRunCntr[12] ;
 wire \freeRunCntr[13] ;
 wire \freeRunCntr[14] ;
 wire \freeRunCntr[15] ;
 wire \freeRunCntr[16] ;
 wire \freeRunCntr[17] ;
 wire \freeRunCntr[1] ;
 wire \freeRunCntr[26] ;
 wire \freeRunCntr[27] ;
 wire \freeRunCntr[28] ;
 wire \freeRunCntr[2] ;
 wire \freeRunCntr[3] ;
 wire \freeRunCntr[4] ;
 wire \freeRunCntr[5] ;
 wire \freeRunCntr[6] ;
 wire \freeRunCntr[7] ;
 wire \freeRunCntr[8] ;
 wire \freeRunCntr[9] ;
 wire \sigRom.address[0] ;
 wire \sigRom.address[1] ;
 wire \sigRom.address[2] ;
 wire \sigRom.address[3] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;

 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1599_ (.I(\csTable.address[7] ),
    .Z(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1600_ (.I(\csTable.address[6] ),
    .Z(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _1601_ (.I(_1334_),
    .Z(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1602_ (.A1(_1323_),
    .A2(_1345_),
    .Z(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _1603_ (.I(_1356_),
    .Z(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _1604_ (.I(_1367_),
    .Z(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _1605_ (.A1(_1345_),
    .A2(\csTable.address[5] ),
    .ZN(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _1606_ (.I(_1389_),
    .Z(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _1607_ (.I(\csTable.address[2] ),
    .Z(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_4 _1608_ (.A1(_1334_),
    .A2(_1411_),
    .Z(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1609_ (.I(\csTable.address[0] ),
    .Z(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1610_ (.A1(_1334_),
    .A2(_1433_),
    .Z(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1611_ (.A1(_1422_),
    .A2(_1444_),
    .ZN(_1455_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1612_ (.I(\csTable.address[1] ),
    .Z(_1466_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_4 _1613_ (.A1(_1334_),
    .A2(_1466_),
    .Z(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1614_ (.A1(_1334_),
    .A2(\csTable.address[3] ),
    .Z(_1488_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1615_ (.A1(_1477_),
    .A2(_1422_),
    .B(_1488_),
    .ZN(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1616_ (.A1(_1455_),
    .A2(_1499_),
    .ZN(_1510_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1617_ (.I(_1488_),
    .Z(_1521_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1618_ (.I(_1521_),
    .Z(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_4 _1619_ (.A1(_1334_),
    .A2(_1466_),
    .ZN(_1543_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _1620_ (.I(_1543_),
    .Z(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _1621_ (.I(_1554_),
    .Z(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_4 _1622_ (.A1(_1345_),
    .A2(_1433_),
    .ZN(_1576_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _1623_ (.I(_1576_),
    .Z(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1624_ (.I(_1587_),
    .Z(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _1625_ (.A1(_1334_),
    .A2(_1411_),
    .ZN(_0043_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1626_ (.I(_0043_),
    .Z(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _1627_ (.I(_0054_),
    .Z(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1628_ (.A1(_1565_),
    .A2(_1598_),
    .B(_0065_),
    .ZN(_0076_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1629_ (.A1(_1345_),
    .A2(\csTable.address[4] ),
    .Z(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1630_ (.I(_0087_),
    .Z(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1631_ (.A1(_1532_),
    .A2(_0076_),
    .B(_0098_),
    .ZN(_0109_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_4 _1632_ (.A1(_1345_),
    .A2(\csTable.address[3] ),
    .ZN(_0120_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1633_ (.I(_0120_),
    .Z(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _1634_ (.I(_1444_),
    .Z(_0142_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _1635_ (.I(_1422_),
    .Z(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1636_ (.A1(_1477_),
    .A2(_0142_),
    .B(_0153_),
    .ZN(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1637_ (.I(_1477_),
    .Z(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _1638_ (.I(_0142_),
    .Z(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1639_ (.A1(_0175_),
    .A2(_0153_),
    .A3(_0186_),
    .ZN(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1640_ (.A1(_1554_),
    .A2(_0054_),
    .B(_0120_),
    .ZN(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1641_ (.A1(_0131_),
    .A2(_0164_),
    .B1(_0197_),
    .B2(_0208_),
    .ZN(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1642_ (.I(_0098_),
    .Z(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1643_ (.A1(_1510_),
    .A2(_0109_),
    .B1(_0219_),
    .B2(_0230_),
    .ZN(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1644_ (.I(_1521_),
    .Z(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1645_ (.A1(_1554_),
    .A2(_0065_),
    .ZN(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1646_ (.A1(_0252_),
    .A2(_0263_),
    .ZN(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1647_ (.I(_0098_),
    .Z(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _1648_ (.A1(_1400_),
    .A2(_0274_),
    .A3(_0285_),
    .A4(_1510_),
    .ZN(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1649_ (.A1(_1400_),
    .A2(_0241_),
    .B(_0296_),
    .ZN(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_4 _1650_ (.A1(_1356_),
    .A2(_0307_),
    .Z(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_4 _1651_ (.A1(_1345_),
    .A2(\csTable.address[4] ),
    .ZN(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1652_ (.A1(_0131_),
    .A2(_0164_),
    .B(_0329_),
    .ZN(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1653_ (.A1(_0285_),
    .A2(_0208_),
    .ZN(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1654_ (.A1(_1400_),
    .A2(_0274_),
    .B1(_0340_),
    .B2(_0351_),
    .ZN(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_4 _1655_ (.A1(_1356_),
    .A2(_0362_),
    .Z(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1656_ (.A1(\freeRunCntr[13] ),
    .A2(_0318_),
    .B1(_0373_),
    .B2(\freeRunCntr[14] ),
    .ZN(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _1657_ (.I(_1323_),
    .ZN(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1658_ (.A1(_0395_),
    .A2(_1345_),
    .Z(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _1659_ (.I(_0406_),
    .Z(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1660_ (.A1(_1345_),
    .A2(\csTable.address[5] ),
    .Z(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1661_ (.I(_0428_),
    .Z(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1662_ (.I(_0439_),
    .Z(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1663_ (.A1(_0450_),
    .A2(_0340_),
    .ZN(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1664_ (.A1(_0417_),
    .A2(_0461_),
    .Z(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1665_ (.A1(\freeRunCntr[14] ),
    .A2(_0373_),
    .B1(_0472_),
    .B2(\freeRunCntr[15] ),
    .ZN(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1666_ (.A1(\freeRunCntr[16] ),
    .A2(_1378_),
    .B1(_0472_),
    .B2(\freeRunCntr[15] ),
    .ZN(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1667_ (.A1(_0384_),
    .A2(_0483_),
    .B(_0494_),
    .ZN(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1668_ (.A1(\freeRunCntr[16] ),
    .A2(_1378_),
    .B(_0505_),
    .ZN(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1669_ (.A1(\freeRunCntr[16] ),
    .A2(_1378_),
    .ZN(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1670_ (.A1(\freeRunCntr[13] ),
    .A2(_0318_),
    .B(_0384_),
    .C(_0494_),
    .ZN(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1671_ (.A1(_0483_),
    .A2(_0527_),
    .A3(_0538_),
    .ZN(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1672_ (.I(\freeRunCntr[9] ),
    .Z(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1673_ (.I(_0131_),
    .Z(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _1674_ (.I(_1422_),
    .Z(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1675_ (.I0(_0175_),
    .I1(_0582_),
    .S(_0186_),
    .Z(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1676_ (.I(_0329_),
    .Z(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1677_ (.A1(_0571_),
    .A2(_0592_),
    .B(_0602_),
    .ZN(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1678_ (.A1(_1422_),
    .A2(_1576_),
    .ZN(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_4 _1679_ (.A1(_1466_),
    .A2(_1433_),
    .Z(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1680_ (.A1(_0043_),
    .A2(_0631_),
    .B(_0120_),
    .ZN(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1681_ (.I(_0285_),
    .Z(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1682_ (.A1(_0622_),
    .A2(_0641_),
    .B(_0651_),
    .C(_1499_),
    .ZN(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _1683_ (.I(_1400_),
    .Z(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1684_ (.A1(_0612_),
    .A2(_0660_),
    .B(_0670_),
    .ZN(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1685_ (.A1(_1433_),
    .A2(_1411_),
    .Z(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _1686_ (.I(_0120_),
    .Z(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1687_ (.A1(_0175_),
    .A2(_0186_),
    .B(_0698_),
    .ZN(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1688_ (.A1(_0252_),
    .A2(_1587_),
    .B(_0098_),
    .ZN(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1689_ (.A1(_0689_),
    .A2(_0707_),
    .B(_0715_),
    .ZN(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _1690_ (.A1(_1565_),
    .A2(_0582_),
    .A3(_0186_),
    .ZN(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1691_ (.A1(_1477_),
    .A2(_1576_),
    .B(_0043_),
    .ZN(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1692_ (.A1(_0582_),
    .A2(_1598_),
    .ZN(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1693_ (.A1(_1565_),
    .A2(_0698_),
    .ZN(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _1694_ (.A1(_0571_),
    .A2(_0730_),
    .A3(_0738_),
    .B1(_0742_),
    .B2(_0743_),
    .ZN(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _1695_ (.A1(_1389_),
    .A2(_0087_),
    .ZN(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1696_ (.A1(_0450_),
    .A2(_0722_),
    .B1(_0744_),
    .B2(_0745_),
    .ZN(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1697_ (.A1(_1378_),
    .A2(_0679_),
    .A3(_0746_),
    .Z(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1698_ (.A1(_0679_),
    .A2(_0746_),
    .B(_1378_),
    .ZN(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__or2_4 _1699_ (.A1(_0747_),
    .A2(_0748_),
    .Z(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1700_ (.I(_1400_),
    .Z(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1701_ (.A1(_1565_),
    .A2(_1598_),
    .B(_0689_),
    .C(_0131_),
    .ZN(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1702_ (.A1(_0571_),
    .A2(_1598_),
    .B(_0751_),
    .C(_0230_),
    .ZN(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1703_ (.A1(_0175_),
    .A2(_0065_),
    .A3(_0186_),
    .ZN(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _1704_ (.A1(_1543_),
    .A2(_1576_),
    .B(_1488_),
    .ZN(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1705_ (.A1(_0753_),
    .A2(_0754_),
    .B(_0602_),
    .ZN(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1706_ (.A1(_0750_),
    .A2(_0752_),
    .A3(_0755_),
    .Z(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _1707_ (.A1(_1543_),
    .A2(_1444_),
    .ZN(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1708_ (.A1(_0730_),
    .A2(_0738_),
    .B(_0757_),
    .C(_0571_),
    .ZN(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1709_ (.A1(_0175_),
    .A2(_0153_),
    .B(_0698_),
    .ZN(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1710_ (.A1(_0631_),
    .A2(_0759_),
    .B(_0651_),
    .ZN(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1711_ (.A1(_1466_),
    .A2(_1411_),
    .Z(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1712_ (.A1(_1598_),
    .A2(_0761_),
    .ZN(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1713_ (.I(_1477_),
    .Z(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1714_ (.I(_0252_),
    .Z(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1715_ (.A1(_0763_),
    .A2(_0764_),
    .B(_0230_),
    .ZN(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1716_ (.A1(_0762_),
    .A2(_0707_),
    .B(_0765_),
    .ZN(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _1717_ (.A1(_0758_),
    .A2(_0760_),
    .B(_0766_),
    .C(_0670_),
    .ZN(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1718_ (.A1(_0756_),
    .A2(_0767_),
    .B(_0417_),
    .ZN(_0768_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _1719_ (.A1(_0406_),
    .A2(_0756_),
    .A3(_0767_),
    .Z(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _1720_ (.A1(_0768_),
    .A2(_0769_),
    .ZN(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1721_ (.A1(_0560_),
    .A2(_0749_),
    .B1(_0770_),
    .B2(\freeRunCntr[10] ),
    .ZN(_0771_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1722_ (.A1(\freeRunCntr[10] ),
    .A2(_0770_),
    .ZN(_0772_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1723_ (.A1(_1554_),
    .A2(_1587_),
    .ZN(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _1724_ (.A1(_1466_),
    .A2(_1411_),
    .ZN(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1725_ (.A1(_0142_),
    .A2(_0774_),
    .ZN(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1726_ (.A1(_0763_),
    .A2(_1532_),
    .B(_0329_),
    .ZN(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1727_ (.A1(_0764_),
    .A2(_0773_),
    .A3(_0775_),
    .B(_0776_),
    .ZN(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1728_ (.I(_1532_),
    .Z(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1729_ (.I(_0329_),
    .Z(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1730_ (.I0(_1422_),
    .I1(_0761_),
    .S(_1444_),
    .Z(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1731_ (.A1(_0778_),
    .A2(_0779_),
    .A3(_0780_),
    .ZN(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1732_ (.A1(_0777_),
    .A2(_0781_),
    .B(_0439_),
    .ZN(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1733_ (.I(_0698_),
    .Z(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _1734_ (.A1(_0783_),
    .A2(_0730_),
    .A3(_0738_),
    .B(_0208_),
    .ZN(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1735_ (.A1(_1532_),
    .A2(_0631_),
    .ZN(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1736_ (.A1(_0230_),
    .A2(_0785_),
    .ZN(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _1737_ (.A1(_1433_),
    .A2(_1411_),
    .ZN(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1738_ (.A1(_0779_),
    .A2(_0787_),
    .ZN(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1739_ (.A1(_0175_),
    .A2(_0065_),
    .ZN(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1740_ (.A1(_0764_),
    .A2(_0789_),
    .ZN(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1741_ (.A1(_0784_),
    .A2(_0786_),
    .B1(_0788_),
    .B2(_0790_),
    .C(_1400_),
    .ZN(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1742_ (.A1(_0782_),
    .A2(_0791_),
    .B(_1367_),
    .ZN(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _1743_ (.A1(_1367_),
    .A2(_0782_),
    .A3(_0791_),
    .Z(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _1744_ (.A1(_0792_),
    .A2(_0793_),
    .Z(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _1745_ (.A1(_1455_),
    .A2(_1499_),
    .B1(_0761_),
    .B2(_1532_),
    .C(_0329_),
    .ZN(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1746_ (.A1(_1554_),
    .A2(_0120_),
    .ZN(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1747_ (.A1(_0065_),
    .A2(_1598_),
    .ZN(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1748_ (.A1(_0796_),
    .A2(_0797_),
    .B(_0285_),
    .ZN(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1749_ (.A1(_0795_),
    .A2(_0798_),
    .B(_1400_),
    .ZN(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1750_ (.A1(_1543_),
    .A2(_1576_),
    .B(_1422_),
    .ZN(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1751_ (.A1(_1488_),
    .A2(_0761_),
    .ZN(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1752_ (.A1(_0153_),
    .A2(_0186_),
    .ZN(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _1753_ (.A1(_1532_),
    .A2(_0800_),
    .A3(_0753_),
    .B1(_0801_),
    .B2(_0802_),
    .ZN(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1754_ (.A1(_1466_),
    .A2(_1433_),
    .ZN(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1755_ (.A1(_0582_),
    .A2(_0804_),
    .B(_0252_),
    .ZN(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _1756_ (.A1(_1477_),
    .A2(_0043_),
    .B(_0120_),
    .ZN(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1757_ (.A1(_0153_),
    .A2(_0631_),
    .ZN(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _1758_ (.A1(_0263_),
    .A2(_0805_),
    .B1(_0806_),
    .B2(_0807_),
    .C(_0098_),
    .ZN(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _1759_ (.A1(_0230_),
    .A2(_0803_),
    .B(_0808_),
    .C(_0439_),
    .ZN(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1760_ (.A1(_1356_),
    .A2(_0799_),
    .A3(_0809_),
    .Z(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1761_ (.A1(_0799_),
    .A2(_0809_),
    .B(_1367_),
    .ZN(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _1762_ (.A1(_0810_),
    .A2(_0811_),
    .ZN(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1763_ (.A1(\freeRunCntr[11] ),
    .A2(_0794_),
    .B1(_0812_),
    .B2(\freeRunCntr[12] ),
    .ZN(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1764_ (.I(\freeRunCntr[11] ),
    .ZN(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1765_ (.A1(_0792_),
    .A2(_0793_),
    .ZN(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1766_ (.A1(\freeRunCntr[12] ),
    .A2(_0812_),
    .ZN(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1767_ (.A1(_0814_),
    .A2(_0815_),
    .B(_0816_),
    .ZN(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1768_ (.A1(_0813_),
    .A2(_0817_),
    .ZN(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _1769_ (.A1(_0771_),
    .A2(_0772_),
    .A3(_0818_),
    .B1(_0816_),
    .B2(_0813_),
    .ZN(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1770_ (.A1(_0730_),
    .A2(_0738_),
    .B(_0757_),
    .ZN(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1771_ (.A1(_0065_),
    .A2(_1587_),
    .ZN(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1772_ (.A1(_1532_),
    .A2(_0821_),
    .B(_0779_),
    .ZN(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1773_ (.A1(_0778_),
    .A2(_0820_),
    .B(_0822_),
    .ZN(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _1774_ (.A1(_1565_),
    .A2(_0065_),
    .A3(_1587_),
    .ZN(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _1775_ (.A1(_1499_),
    .A2(_0824_),
    .B1(_0631_),
    .B2(_0778_),
    .C(_0779_),
    .ZN(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1776_ (.A1(_0054_),
    .A2(_0142_),
    .B(_0774_),
    .ZN(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1777_ (.I(_0186_),
    .Z(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1778_ (.A1(_0763_),
    .A2(_0827_),
    .ZN(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1779_ (.A1(_0783_),
    .A2(_0828_),
    .ZN(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1780_ (.A1(_0821_),
    .A2(_0743_),
    .ZN(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _1781_ (.A1(_0826_),
    .A2(_0829_),
    .B(_0830_),
    .C(_0602_),
    .ZN(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1782_ (.A1(_0175_),
    .A2(_0186_),
    .B(_0698_),
    .ZN(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _1783_ (.A1(_0783_),
    .A2(_0821_),
    .B1(_0164_),
    .B2(_0832_),
    .C(_0779_),
    .ZN(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1784_ (.A1(_0750_),
    .A2(_0833_),
    .ZN(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _1785_ (.A1(_0750_),
    .A2(_0823_),
    .A3(_0825_),
    .B1(_0831_),
    .B2(_0834_),
    .ZN(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_4 _1786_ (.A1(_1367_),
    .A2(_0835_),
    .Z(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _1787_ (.A1(_0698_),
    .A2(_0780_),
    .B1(_0800_),
    .B2(_0806_),
    .C(_0087_),
    .ZN(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1788_ (.A1(_0120_),
    .A2(_0054_),
    .A3(_0804_),
    .ZN(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1789_ (.A1(_0153_),
    .A2(_0142_),
    .B1(_0631_),
    .B2(_1521_),
    .C(_0087_),
    .ZN(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1790_ (.A1(_0838_),
    .A2(_0839_),
    .B(_1389_),
    .ZN(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1791_ (.A1(_1521_),
    .A2(_1587_),
    .ZN(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _1792_ (.A1(_0120_),
    .A2(_0142_),
    .A3(_0761_),
    .ZN(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1793_ (.A1(_0826_),
    .A2(_0841_),
    .B(_0842_),
    .C(_0098_),
    .ZN(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1794_ (.A1(_0153_),
    .A2(_0142_),
    .B(_0087_),
    .ZN(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1795_ (.I0(_0120_),
    .I1(_0054_),
    .S(_1543_),
    .Z(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1796_ (.A1(_0844_),
    .A2(_0845_),
    .B(_0428_),
    .ZN(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1797_ (.A1(_0837_),
    .A2(_0840_),
    .B1(_0843_),
    .B2(_0846_),
    .ZN(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_4 _1798_ (.A1(_0406_),
    .A2(_0847_),
    .Z(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1799_ (.I(_0054_),
    .Z(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1800_ (.A1(_0763_),
    .A2(_0849_),
    .B(_1598_),
    .ZN(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1801_ (.A1(_0775_),
    .A2(_0850_),
    .B(_0764_),
    .ZN(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1802_ (.A1(_0153_),
    .A2(_1587_),
    .B(_1521_),
    .ZN(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1803_ (.A1(_0450_),
    .A2(_0852_),
    .ZN(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1804_ (.A1(_0065_),
    .A2(_0186_),
    .B(_0698_),
    .ZN(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1805_ (.A1(_0763_),
    .A2(_1598_),
    .ZN(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _1806_ (.A1(_1499_),
    .A2(_0757_),
    .B1(_0854_),
    .B2(_0855_),
    .C(_0750_),
    .ZN(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1807_ (.I(_0779_),
    .Z(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _1808_ (.A1(_0851_),
    .A2(_0853_),
    .B(_0856_),
    .C(_0857_),
    .ZN(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _1809_ (.A1(_0750_),
    .A2(_0263_),
    .A3(_0807_),
    .Z(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1810_ (.A1(_0670_),
    .A2(_0850_),
    .B(_0571_),
    .ZN(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1811_ (.A1(_0208_),
    .A2(_0828_),
    .B(_0857_),
    .ZN(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1812_ (.A1(_0859_),
    .A2(_0860_),
    .B(_0861_),
    .ZN(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _1813_ (.A1(_0417_),
    .A2(_0858_),
    .A3(_0862_),
    .Z(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1814_ (.A1(_0858_),
    .A2(_0862_),
    .B(_0417_),
    .ZN(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1815_ (.A1(_0863_),
    .A2(_0864_),
    .Z(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1816_ (.A1(_0778_),
    .A2(_0802_),
    .B(_0651_),
    .ZN(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1817_ (.A1(_1422_),
    .A2(_1444_),
    .B(_1488_),
    .ZN(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1818_ (.A1(_0763_),
    .A2(_0849_),
    .ZN(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1819_ (.A1(_0763_),
    .A2(_1598_),
    .B(_0783_),
    .ZN(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _1820_ (.A1(_0867_),
    .A2(_0868_),
    .B1(_0787_),
    .B2(_0869_),
    .C(_0602_),
    .ZN(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _1821_ (.A1(_0866_),
    .A2(_0842_),
    .B(_0439_),
    .C(_0870_),
    .ZN(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1822_ (.A1(_1565_),
    .A2(_0582_),
    .ZN(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1823_ (.A1(_1477_),
    .A2(_1576_),
    .ZN(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1824_ (.A1(_1422_),
    .A2(_1587_),
    .B(_1521_),
    .ZN(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _1825_ (.A1(_0778_),
    .A2(_0797_),
    .A3(_0872_),
    .B1(_0873_),
    .B2(_0874_),
    .ZN(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1826_ (.A1(_1477_),
    .A2(_0142_),
    .B(_0054_),
    .ZN(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1827_ (.A1(_0876_),
    .A2(_0707_),
    .B(_0715_),
    .C(_1499_),
    .ZN(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _1828_ (.A1(_0857_),
    .A2(_0875_),
    .B(_0877_),
    .C(_0750_),
    .ZN(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _1829_ (.A1(_1367_),
    .A2(_0871_),
    .A3(_0878_),
    .Z(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1830_ (.A1(_0871_),
    .A2(_0878_),
    .B(_1367_),
    .ZN(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1831_ (.A1(_0879_),
    .A2(_0880_),
    .Z(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1832_ (.I(\freeRunCntr[5] ),
    .Z(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1833_ (.I(\freeRunCntr[4] ),
    .ZN(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _1834_ (.A1(_0863_),
    .A2(_0864_),
    .ZN(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1835_ (.I(\freeRunCntr[3] ),
    .ZN(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1836_ (.A1(_0592_),
    .A2(_0765_),
    .Z(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1837_ (.A1(_0775_),
    .A2(_0754_),
    .B(_0857_),
    .C(_0208_),
    .ZN(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1838_ (.A1(_0886_),
    .A2(_0887_),
    .B(_0450_),
    .ZN(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1839_ (.A1(_0428_),
    .A2(_0285_),
    .ZN(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1840_ (.A1(_1565_),
    .A2(_0582_),
    .A3(_0827_),
    .B(_0131_),
    .ZN(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1841_ (.A1(_0738_),
    .A2(_0873_),
    .A3(_0890_),
    .ZN(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1842_ (.A1(_0571_),
    .A2(_0849_),
    .A3(_0631_),
    .ZN(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1843_ (.A1(_0849_),
    .A2(_0827_),
    .ZN(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1844_ (.A1(_0175_),
    .A2(_0252_),
    .ZN(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1845_ (.A1(_0893_),
    .A2(_0894_),
    .B1(_0757_),
    .B2(_0759_),
    .ZN(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1846_ (.A1(_0428_),
    .A2(_0329_),
    .ZN(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _1847_ (.A1(_0889_),
    .A2(_0891_),
    .A3(_0892_),
    .B1(_0895_),
    .B2(_0896_),
    .ZN(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _1848_ (.A1(_0417_),
    .A2(_0888_),
    .A3(_0897_),
    .Z(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1849_ (.A1(_0888_),
    .A2(_0897_),
    .B(_0417_),
    .ZN(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _1850_ (.A1(_0898_),
    .A2(_0899_),
    .Z(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1851_ (.A1(_0885_),
    .A2(_0900_),
    .ZN(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1852_ (.A1(_0175_),
    .A2(_0582_),
    .ZN(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _1853_ (.A1(_0763_),
    .A2(_0827_),
    .B1(_0902_),
    .B2(_0754_),
    .C(_0651_),
    .ZN(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1854_ (.A1(_0873_),
    .A2(_0874_),
    .B(_0890_),
    .C(_0857_),
    .ZN(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1855_ (.A1(_0903_),
    .A2(_0904_),
    .B(_0670_),
    .ZN(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1856_ (.A1(_0698_),
    .A2(_0065_),
    .A3(_0631_),
    .ZN(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1857_ (.A1(_0805_),
    .A2(_0906_),
    .B(_0775_),
    .ZN(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1858_ (.A1(_0263_),
    .A2(_0742_),
    .B(_0571_),
    .ZN(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1859_ (.A1(_0651_),
    .A2(_0707_),
    .ZN(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _1860_ (.A1(_0651_),
    .A2(_0907_),
    .B1(_0908_),
    .B2(_0909_),
    .C(_0450_),
    .ZN(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _1861_ (.A1(_1378_),
    .A2(_0905_),
    .A3(_0910_),
    .Z(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1862_ (.A1(_0905_),
    .A2(_0910_),
    .B(_1378_),
    .ZN(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _1863_ (.A1(_0911_),
    .A2(_0912_),
    .Z(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1864_ (.A1(\freeRunCntr[2] ),
    .A2(_0913_),
    .ZN(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1865_ (.A1(_0043_),
    .A2(_1444_),
    .ZN(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _1866_ (.A1(_0802_),
    .A2(_0789_),
    .B1(_0915_),
    .B2(_0743_),
    .C(_0602_),
    .ZN(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1867_ (.A1(_1554_),
    .A2(_1521_),
    .B(_0329_),
    .ZN(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1868_ (.A1(_0571_),
    .A2(_0821_),
    .B(_0751_),
    .C(_0917_),
    .ZN(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1869_ (.A1(_0916_),
    .A2(_0918_),
    .Z(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1870_ (.A1(_0827_),
    .A2(_0774_),
    .ZN(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1871_ (.A1(_0873_),
    .A2(_0874_),
    .B(_0920_),
    .C(_0762_),
    .ZN(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1872_ (.A1(_0730_),
    .A2(_0738_),
    .B(_0757_),
    .C(_0854_),
    .ZN(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1873_ (.A1(_0651_),
    .A2(_0921_),
    .A3(_0922_),
    .Z(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1874_ (.A1(_0651_),
    .A2(_0867_),
    .A3(_0775_),
    .B(_0750_),
    .ZN(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _1875_ (.A1(_0670_),
    .A2(_0919_),
    .B1(_0923_),
    .B2(_0924_),
    .ZN(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1876_ (.A1(_0417_),
    .A2(_0925_),
    .Z(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1877_ (.A1(\freeRunCntr[2] ),
    .A2(_0913_),
    .B(_0926_),
    .C(\freeRunCntr[1] ),
    .ZN(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1878_ (.A1(_0885_),
    .A2(_0900_),
    .B1(_0914_),
    .B2(_0927_),
    .ZN(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1879_ (.A1(_0901_),
    .A2(_0928_),
    .ZN(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1880_ (.A1(_0883_),
    .A2(_0884_),
    .B(_0929_),
    .ZN(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _1881_ (.A1(\freeRunCntr[4] ),
    .A2(_0865_),
    .B1(_0881_),
    .B2(_0882_),
    .C(_0930_),
    .ZN(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1882_ (.A1(_1565_),
    .A2(_0827_),
    .B(_1532_),
    .ZN(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _1883_ (.A1(_0764_),
    .A2(_0775_),
    .B1(_0932_),
    .B2(_0802_),
    .C(_0230_),
    .ZN(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1884_ (.A1(_1554_),
    .A2(_0142_),
    .B(_0054_),
    .ZN(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _1885_ (.A1(_0902_),
    .A2(_0754_),
    .B1(_0934_),
    .B2(_0764_),
    .C(_0779_),
    .ZN(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1886_ (.A1(_0933_),
    .A2(_0935_),
    .B(_0439_),
    .ZN(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1887_ (.I0(_0175_),
    .I1(_0582_),
    .S(_1598_),
    .Z(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1888_ (.A1(_0783_),
    .A2(_0937_),
    .B(_0230_),
    .ZN(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _1889_ (.A1(_1499_),
    .A2(_0824_),
    .B1(_0757_),
    .B2(_0854_),
    .C(_0779_),
    .ZN(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _1890_ (.A1(_0851_),
    .A2(_0938_),
    .B(_0939_),
    .C(_0750_),
    .ZN(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _1891_ (.A1(_1367_),
    .A2(_0936_),
    .A3(_0940_),
    .Z(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1892_ (.A1(_0936_),
    .A2(_0940_),
    .B(_1367_),
    .ZN(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1893_ (.A1(_0941_),
    .A2(_0942_),
    .Z(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1894_ (.A1(_0882_),
    .A2(_0881_),
    .B1(_0943_),
    .B2(\freeRunCntr[6] ),
    .ZN(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1895_ (.A1(_0406_),
    .A2(_0835_),
    .Z(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1896_ (.I(\freeRunCntr[7] ),
    .ZN(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1897_ (.A1(\freeRunCntr[6] ),
    .A2(_0943_),
    .ZN(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1898_ (.A1(_0931_),
    .A2(_0944_),
    .B1(_0945_),
    .B2(_0946_),
    .C(_0947_),
    .ZN(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1899_ (.A1(\freeRunCntr[7] ),
    .A2(_0836_),
    .B1(_0848_),
    .B2(\freeRunCntr[8] ),
    .C(_0948_),
    .ZN(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _1900_ (.A1(_0560_),
    .A2(_0749_),
    .B1(_0770_),
    .B2(\freeRunCntr[10] ),
    .C(_0549_),
    .ZN(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1901_ (.A1(\freeRunCntr[8] ),
    .A2(_0848_),
    .B(_0771_),
    .ZN(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _1902_ (.A1(_0818_),
    .A2(_0949_),
    .A3(_0950_),
    .A4(_0951_),
    .ZN(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1903_ (.A1(_0549_),
    .A2(_0819_),
    .B(_0952_),
    .ZN(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1904_ (.A1(_0516_),
    .A2(_0953_),
    .Z(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1905_ (.I(_0954_),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _1906_ (.I(_1323_),
    .Z(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1907_ (.A1(_0783_),
    .A2(_0849_),
    .ZN(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1908_ (.A1(_0956_),
    .A2(_0351_),
    .ZN(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1909_ (.A1(_0857_),
    .A2(_0219_),
    .B(_0957_),
    .ZN(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1910_ (.A1(_0783_),
    .A2(_0164_),
    .ZN(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1911_ (.A1(_0745_),
    .A2(_0959_),
    .ZN(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1912_ (.A1(_0450_),
    .A2(_0958_),
    .B1(_0960_),
    .B2(_0956_),
    .ZN(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1913_ (.A1(_0955_),
    .A2(_0961_),
    .Z(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1914_ (.A1(_0340_),
    .A2(_0351_),
    .Z(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _1915_ (.A1(_0450_),
    .A2(_0963_),
    .A3(_0830_),
    .B1(_0959_),
    .B2(_0896_),
    .ZN(_0964_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1916_ (.A1(_0955_),
    .A2(_0964_),
    .Z(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1917_ (.A1(\freeRunCntr[13] ),
    .A2(_0962_),
    .B1(_0965_),
    .B2(\freeRunCntr[14] ),
    .ZN(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1918_ (.A1(_0857_),
    .A2(_0830_),
    .ZN(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1919_ (.A1(_0670_),
    .A2(_0351_),
    .A3(_0967_),
    .ZN(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1920_ (.A1(_0395_),
    .A2(_0968_),
    .Z(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1921_ (.A1(\freeRunCntr[15] ),
    .A2(_0969_),
    .B1(_0965_),
    .B2(\freeRunCntr[14] ),
    .ZN(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1922_ (.A1(_0450_),
    .A2(_0967_),
    .ZN(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1923_ (.A1(_0955_),
    .A2(_0971_),
    .Z(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1924_ (.A1(\freeRunCntr[16] ),
    .A2(_0972_),
    .B1(_0969_),
    .B2(\freeRunCntr[15] ),
    .ZN(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1925_ (.A1(_0966_),
    .A2(_0970_),
    .B(_0973_),
    .ZN(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1926_ (.A1(\freeRunCntr[16] ),
    .A2(_0972_),
    .Z(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1927_ (.A1(_0131_),
    .A2(_0902_),
    .ZN(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1928_ (.A1(_0849_),
    .A2(_0841_),
    .B(_0842_),
    .ZN(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1929_ (.A1(_0745_),
    .A2(_0977_),
    .ZN(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1930_ (.A1(_1554_),
    .A2(_0054_),
    .B(_1521_),
    .ZN(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _1931_ (.A1(_0787_),
    .A2(_0979_),
    .A3(_0873_),
    .B1(_0807_),
    .B2(_0806_),
    .ZN(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1932_ (.A1(_0800_),
    .A2(_0754_),
    .B(_0098_),
    .ZN(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1933_ (.A1(_0065_),
    .A2(_0773_),
    .B(_0806_),
    .ZN(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _1934_ (.A1(_0285_),
    .A2(_0980_),
    .B1(_0981_),
    .B2(_0982_),
    .C(_1389_),
    .ZN(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1935_ (.A1(_0889_),
    .A2(_0976_),
    .B(_0978_),
    .C(_0983_),
    .ZN(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1936_ (.A1(_1323_),
    .A2(_0984_),
    .Z(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1937_ (.A1(_1554_),
    .A2(_0142_),
    .B(_0153_),
    .ZN(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1938_ (.A1(_0986_),
    .A2(_0757_),
    .B(_0698_),
    .ZN(_0987_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1939_ (.A1(_1587_),
    .A2(_0774_),
    .Z(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _1940_ (.A1(_0787_),
    .A2(_0806_),
    .B1(_0988_),
    .B2(_0783_),
    .C(_0602_),
    .ZN(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1941_ (.A1(_0602_),
    .A2(_0891_),
    .A3(_0987_),
    .B(_0989_),
    .ZN(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1942_ (.A1(_0131_),
    .A2(_0804_),
    .ZN(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1943_ (.A1(_0800_),
    .A2(_0754_),
    .B(_0991_),
    .ZN(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1944_ (.A1(_0902_),
    .A2(_0889_),
    .ZN(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1945_ (.A1(_0745_),
    .A2(_0992_),
    .B1(_0993_),
    .B2(_1499_),
    .ZN(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1946_ (.A1(_0450_),
    .A2(_0990_),
    .B(_0994_),
    .ZN(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1947_ (.A1(_0955_),
    .A2(_0995_),
    .Z(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1948_ (.A1(\freeRunCntr[12] ),
    .A2(_0985_),
    .B1(_0996_),
    .B2(\freeRunCntr[11] ),
    .ZN(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1949_ (.A1(_1565_),
    .A2(_0827_),
    .ZN(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1950_ (.A1(_0915_),
    .A2(_0743_),
    .B(_0602_),
    .ZN(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1951_ (.A1(_0764_),
    .A2(_0988_),
    .ZN(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1952_ (.A1(_0991_),
    .A2(_0976_),
    .A3(_1000_),
    .Z(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _1953_ (.A1(_0796_),
    .A2(_0998_),
    .A3(_0999_),
    .B1(_1001_),
    .B2(_0857_),
    .ZN(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1954_ (.A1(_0778_),
    .A2(_0824_),
    .B(_0765_),
    .C(_0750_),
    .ZN(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1955_ (.A1(_0915_),
    .A2(_0759_),
    .B1(_0801_),
    .B2(_0827_),
    .ZN(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1956_ (.A1(_0896_),
    .A2(_1004_),
    .ZN(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1957_ (.A1(_0670_),
    .A2(_1002_),
    .B(_1003_),
    .C(_1005_),
    .ZN(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1958_ (.A1(_0395_),
    .A2(_1006_),
    .Z(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1959_ (.A1(_0582_),
    .A2(_1587_),
    .B(_0761_),
    .ZN(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1960_ (.A1(_0252_),
    .A2(_1008_),
    .B(_0329_),
    .ZN(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1961_ (.A1(_0764_),
    .A2(_0988_),
    .B(_1009_),
    .ZN(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _1962_ (.A1(_0787_),
    .A2(_0979_),
    .B1(_0806_),
    .B2(_0800_),
    .C(_0098_),
    .ZN(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1963_ (.A1(_0439_),
    .A2(_1011_),
    .ZN(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1964_ (.A1(_0773_),
    .A2(_0775_),
    .ZN(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _1965_ (.A1(_0783_),
    .A2(_1013_),
    .B1(_0641_),
    .B2(_1455_),
    .C(_0329_),
    .ZN(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1966_ (.A1(_1532_),
    .A2(_0285_),
    .A3(_0800_),
    .B(_1400_),
    .ZN(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _1967_ (.A1(_1010_),
    .A2(_1012_),
    .B1(_1014_),
    .B2(_1015_),
    .ZN(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1968_ (.A1(_0955_),
    .A2(_1016_),
    .Z(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1969_ (.A1(_0764_),
    .A2(_0937_),
    .Z(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1970_ (.A1(_0641_),
    .A2(_0715_),
    .B1(_1009_),
    .B2(_1018_),
    .ZN(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1971_ (.A1(_1477_),
    .A2(_1422_),
    .ZN(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1972_ (.A1(_0689_),
    .A2(_0894_),
    .B(_0779_),
    .C(_0998_),
    .ZN(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1973_ (.A1(_0764_),
    .A2(_0827_),
    .B1(_0867_),
    .B2(_0934_),
    .C(_0285_),
    .ZN(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1974_ (.A1(_1020_),
    .A2(_1021_),
    .B(_1022_),
    .C(_0439_),
    .ZN(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1975_ (.A1(_0450_),
    .A2(_1019_),
    .B(_1023_),
    .ZN(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1976_ (.A1(_0395_),
    .A2(_1024_),
    .Z(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1977_ (.A1(_0131_),
    .A2(_0780_),
    .Z(_1026_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1978_ (.A1(_0821_),
    .A2(_0894_),
    .ZN(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1979_ (.A1(_1026_),
    .A2(_1027_),
    .B(_0439_),
    .C(_0230_),
    .ZN(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1980_ (.A1(_0631_),
    .A2(_0689_),
    .B(_0698_),
    .ZN(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1981_ (.A1(_0131_),
    .A2(_0826_),
    .B(_1029_),
    .C(_0285_),
    .ZN(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1982_ (.A1(_1499_),
    .A2(_0824_),
    .B1(_0622_),
    .B2(_0759_),
    .C(_0715_),
    .ZN(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1983_ (.A1(_0774_),
    .A2(_0832_),
    .B(_0917_),
    .C(_1389_),
    .ZN(_1032_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1984_ (.A1(_1400_),
    .A2(_1030_),
    .A3(_1031_),
    .B(_1032_),
    .ZN(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1985_ (.A1(_1028_),
    .A2(_1033_),
    .ZN(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1986_ (.A1(_1323_),
    .A2(_1034_),
    .Z(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1987_ (.A1(_1521_),
    .A2(_0915_),
    .B1(_0641_),
    .B2(_1020_),
    .ZN(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1988_ (.A1(_0867_),
    .A2(_0934_),
    .B(_0087_),
    .ZN(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1989_ (.A1(_1477_),
    .A2(_1576_),
    .B(_0787_),
    .ZN(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1990_ (.A1(_0787_),
    .A2(_0754_),
    .B1(_1038_),
    .B2(_1521_),
    .ZN(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1991_ (.A1(_1036_),
    .A2(_1037_),
    .B1(_1039_),
    .B2(_0098_),
    .C(_0428_),
    .ZN(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1992_ (.A1(_0186_),
    .A2(_0806_),
    .B1(_0801_),
    .B2(_0689_),
    .ZN(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1993_ (.A1(_0745_),
    .A2(_1041_),
    .Z(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _1994_ (.A1(_0428_),
    .A2(_1510_),
    .A3(_0874_),
    .A4(_0917_),
    .Z(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _1995_ (.A1(_1040_),
    .A2(_1042_),
    .A3(_1043_),
    .Z(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1996_ (.A1(_1323_),
    .A2(_1044_),
    .Z(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1997_ (.A1(_0849_),
    .A2(_0785_),
    .ZN(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1998_ (.A1(_1565_),
    .A2(_0849_),
    .ZN(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1999_ (.I0(_0054_),
    .I1(_0761_),
    .S(_1576_),
    .Z(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2000_ (.A1(_1047_),
    .A2(_0841_),
    .B1(_1048_),
    .B2(_1532_),
    .ZN(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2001_ (.A1(_0822_),
    .A2(_1046_),
    .B1(_1049_),
    .B2(_0602_),
    .ZN(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2002_ (.A1(_0763_),
    .A2(_0689_),
    .B(_0285_),
    .ZN(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _2003_ (.A1(_0252_),
    .A2(_0802_),
    .A3(_0773_),
    .A4(_0789_),
    .Z(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2004_ (.A1(_1047_),
    .A2(_0707_),
    .B(_0779_),
    .ZN(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2005_ (.A1(_1036_),
    .A2(_1051_),
    .B1(_1052_),
    .B2(_1053_),
    .C(_1400_),
    .ZN(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2006_ (.A1(_0750_),
    .A2(_1050_),
    .B(_1054_),
    .ZN(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _2007_ (.A1(_0395_),
    .A2(_1055_),
    .Z(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2008_ (.A1(_0852_),
    .A2(_0876_),
    .B1(_1048_),
    .B2(_0252_),
    .ZN(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2009_ (.A1(_0896_),
    .A2(_1057_),
    .ZN(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2010_ (.A1(_0252_),
    .A2(_1038_),
    .B(_0098_),
    .ZN(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2011_ (.A1(_0796_),
    .A2(_0622_),
    .B(_0867_),
    .C(_0329_),
    .ZN(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _2012_ (.A1(_0906_),
    .A2(_1059_),
    .B(_1060_),
    .C(_0428_),
    .ZN(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2013_ (.A1(_0252_),
    .A2(_0738_),
    .A3(_0873_),
    .ZN(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _2014_ (.A1(_1554_),
    .A2(_0120_),
    .A3(_0153_),
    .B(_0087_),
    .ZN(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _2015_ (.A1(_1389_),
    .A2(_1062_),
    .A3(_0987_),
    .A4(_1063_),
    .ZN(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _2016_ (.A1(_0395_),
    .A2(_1058_),
    .A3(_1061_),
    .A4(_1064_),
    .Z(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _2017_ (.A1(_1058_),
    .A2(_1061_),
    .A3(_1064_),
    .B(_0395_),
    .ZN(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2018_ (.A1(_1065_),
    .A2(_1066_),
    .ZN(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2019_ (.A1(_0857_),
    .A2(_0890_),
    .ZN(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2020_ (.A1(_0797_),
    .A2(_0979_),
    .A3(_0807_),
    .ZN(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2021_ (.A1(_0796_),
    .A2(_0797_),
    .B1(_0805_),
    .B2(_0920_),
    .ZN(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2022_ (.A1(_1068_),
    .A2(_1069_),
    .B1(_1070_),
    .B2(_0857_),
    .ZN(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2023_ (.A1(_0274_),
    .A2(_0612_),
    .ZN(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2024_ (.A1(_0571_),
    .A2(_0876_),
    .A3(_0757_),
    .ZN(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2025_ (.A1(_0778_),
    .A2(_0800_),
    .B(_0651_),
    .ZN(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2026_ (.A1(_1073_),
    .A2(_1074_),
    .B(_0670_),
    .ZN(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2027_ (.A1(_0670_),
    .A2(_1071_),
    .B1(_1072_),
    .B2(_1075_),
    .ZN(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2028_ (.A1(_0955_),
    .A2(_1076_),
    .Z(_1077_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2029_ (.I(_1077_),
    .Z(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2030_ (.I(_1078_),
    .ZN(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2031_ (.A1(_0778_),
    .A2(_0762_),
    .B1(_0631_),
    .B2(_0821_),
    .ZN(_1080_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2032_ (.A1(_0778_),
    .A2(_1047_),
    .B(_0991_),
    .C(_0917_),
    .ZN(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2033_ (.A1(_0651_),
    .A2(_1080_),
    .B(_1081_),
    .ZN(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2034_ (.A1(_0571_),
    .A2(_0937_),
    .Z(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _2035_ (.A1(_0849_),
    .A2(_0991_),
    .B1(_1083_),
    .B2(_0738_),
    .ZN(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2036_ (.A1(_0778_),
    .A2(_0787_),
    .ZN(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2037_ (.A1(_1085_),
    .A2(_0757_),
    .B1(_0854_),
    .B2(_0855_),
    .C(_0889_),
    .ZN(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2038_ (.A1(_0670_),
    .A2(_1082_),
    .B1(_1084_),
    .B2(_0745_),
    .C(_1086_),
    .ZN(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2039_ (.A1(_0395_),
    .A2(_1087_),
    .Z(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2040_ (.A1(\freeRunCntr[2] ),
    .A2(_1079_),
    .B(_1088_),
    .C(\freeRunCntr[1] ),
    .ZN(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2041_ (.A1(_0783_),
    .A2(_0988_),
    .ZN(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2042_ (.A1(_0790_),
    .A2(_1090_),
    .B(_0602_),
    .ZN(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2043_ (.A1(_0763_),
    .A2(_0131_),
    .A3(_0827_),
    .B(_0842_),
    .ZN(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _2044_ (.A1(_0582_),
    .A2(_0998_),
    .B(_1092_),
    .C(_0230_),
    .ZN(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _2045_ (.A1(_0230_),
    .A2(_0592_),
    .B1(_0754_),
    .B2(_0849_),
    .C(_1063_),
    .ZN(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2046_ (.A1(_0439_),
    .A2(_1094_),
    .ZN(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _2047_ (.A1(_0439_),
    .A2(_1091_),
    .A3(_1093_),
    .B(_1095_),
    .ZN(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _2048_ (.A1(_1323_),
    .A2(_1096_),
    .Z(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2049_ (.A1(\freeRunCntr[2] ),
    .A2(_1079_),
    .B1(_1097_),
    .B2(\freeRunCntr[3] ),
    .ZN(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2050_ (.A1(\freeRunCntr[3] ),
    .A2(_1097_),
    .B1(_1056_),
    .B2(\freeRunCntr[4] ),
    .ZN(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2051_ (.A1(_1089_),
    .A2(_1098_),
    .B(_1099_),
    .ZN(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _2052_ (.A1(\freeRunCntr[4] ),
    .A2(_1056_),
    .B1(_1067_),
    .B2(_0882_),
    .C(_1100_),
    .ZN(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2053_ (.A1(_0882_),
    .A2(_1067_),
    .B1(_1045_),
    .B2(\freeRunCntr[6] ),
    .ZN(_1102_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2054_ (.A1(_1101_),
    .A2(_1102_),
    .B1(_1035_),
    .B2(_0946_),
    .ZN(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2055_ (.A1(\freeRunCntr[6] ),
    .A2(_1045_),
    .B(_1103_),
    .ZN(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2056_ (.A1(\freeRunCntr[8] ),
    .A2(_1017_),
    .ZN(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2057_ (.A1(_0946_),
    .A2(_1035_),
    .B(_1104_),
    .C(_1105_),
    .ZN(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _2058_ (.A1(\freeRunCntr[8] ),
    .A2(_1017_),
    .B1(_1025_),
    .B2(_0560_),
    .C(_1106_),
    .ZN(_1107_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2059_ (.A1(_0560_),
    .A2(_1025_),
    .B1(_1007_),
    .B2(\freeRunCntr[10] ),
    .ZN(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2060_ (.A1(_1107_),
    .A2(_1108_),
    .ZN(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _2061_ (.A1(\freeRunCntr[11] ),
    .A2(_0996_),
    .B1(_1007_),
    .B2(\freeRunCntr[10] ),
    .C(_1109_),
    .ZN(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2062_ (.A1(\freeRunCntr[13] ),
    .A2(_0962_),
    .B(_0975_),
    .C(_0973_),
    .ZN(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2063_ (.A1(_0970_),
    .A2(_1111_),
    .ZN(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2064_ (.A1(\freeRunCntr[12] ),
    .A2(_0985_),
    .B(_1112_),
    .ZN(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2065_ (.A1(_0997_),
    .A2(_1110_),
    .B(_1113_),
    .ZN(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2066_ (.A1(_0974_),
    .A2(_0975_),
    .B1(_1114_),
    .B2(_0966_),
    .ZN(net8));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2067_ (.I(\sigRom.address[2] ),
    .Z(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _2068_ (.I(_1115_),
    .ZN(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2069_ (.I(\sigRom.address[1] ),
    .Z(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _2070_ (.I(\sigRom.address[3] ),
    .Z(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _2071_ (.A1(_1116_),
    .A2(_1117_),
    .A3(_1118_),
    .ZN(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _2072_ (.A1(_0985_),
    .A2(_1119_),
    .ZN(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _2073_ (.A1(_1007_),
    .A2(_1119_),
    .ZN(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _2074_ (.A1(_1115_),
    .A2(\sigRom.address[0] ),
    .A3(_1117_),
    .B(_1118_),
    .ZN(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _2075_ (.I(_1118_),
    .ZN(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2076_ (.A1(_1115_),
    .A2(\sigRom.address[0] ),
    .A3(_1117_),
    .ZN(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2077_ (.A1(_1123_),
    .A2(_1124_),
    .ZN(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2078_ (.A1(_1122_),
    .A2(_1125_),
    .ZN(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2079_ (.A1(_1045_),
    .A2(_1119_),
    .B1(_1126_),
    .B2(_1067_),
    .ZN(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2080_ (.A1(_1121_),
    .A2(_1127_),
    .Z(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2081_ (.A1(_0996_),
    .A2(_1119_),
    .Z(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2082_ (.A1(_1117_),
    .A2(_1118_),
    .ZN(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2083_ (.A1(_1115_),
    .A2(_1130_),
    .ZN(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _2084_ (.A1(_1035_),
    .A2(_1131_),
    .Z(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2085_ (.A1(_1045_),
    .A2(_1126_),
    .ZN(_1133_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2086_ (.A1(_1132_),
    .A2(_1133_),
    .ZN(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2087_ (.A1(_1129_),
    .A2(_1134_),
    .Z(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2088_ (.A1(_1128_),
    .A2(_1135_),
    .Z(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2089_ (.A1(_1128_),
    .A2(_1135_),
    .Z(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2090_ (.A1(_1120_),
    .A2(_1136_),
    .B(_1137_),
    .ZN(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2091_ (.A1(_0417_),
    .A2(_0307_),
    .Z(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _2092_ (.I(\sigRom.address[0] ),
    .ZN(_1140_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _2093_ (.A1(_1115_),
    .A2(_1140_),
    .A3(_1123_),
    .ZN(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _2094_ (.I(_1141_),
    .Z(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2095_ (.A1(_1139_),
    .A2(_1142_),
    .ZN(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2096_ (.A1(_1115_),
    .A2(_1123_),
    .ZN(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2097_ (.A1(_1117_),
    .A2(_1144_),
    .ZN(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2098_ (.A1(_1077_),
    .A2(_1145_),
    .ZN(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2099_ (.A1(_1140_),
    .A2(_1118_),
    .ZN(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2100_ (.A1(\sigRom.address[1] ),
    .A2(_1147_),
    .Z(_1148_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2101_ (.A1(\sigRom.address[1] ),
    .A2(_1147_),
    .B(_1115_),
    .ZN(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2102_ (.A1(_1148_),
    .A2(_1149_),
    .ZN(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2103_ (.I(_1150_),
    .Z(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _2104_ (.A1(_1143_),
    .A2(_1146_),
    .B(_1097_),
    .C(_1151_),
    .ZN(_1152_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2105_ (.I(_1152_),
    .ZN(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2106_ (.A1(_0941_),
    .A2(_0942_),
    .ZN(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2107_ (.A1(_1154_),
    .A2(_1142_),
    .ZN(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _2108_ (.A1(_0768_),
    .A2(_0769_),
    .A3(_1141_),
    .ZN(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2109_ (.A1(_0768_),
    .A2(_0769_),
    .Z(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _2110_ (.A1(_1116_),
    .A2(\sigRom.address[0] ),
    .A3(_1118_),
    .ZN(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _2111_ (.A1(_0941_),
    .A2(_0942_),
    .B(_1158_),
    .ZN(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2112_ (.I0(_1156_),
    .I1(_1157_),
    .S(_1159_),
    .Z(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2113_ (.A1(_0815_),
    .A2(_1142_),
    .ZN(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2114_ (.A1(_0770_),
    .A2(_1155_),
    .B1(_1160_),
    .B2(_1161_),
    .ZN(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2115_ (.A1(_1056_),
    .A2(_1150_),
    .ZN(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2116_ (.A1(_1117_),
    .A2(_1144_),
    .Z(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2117_ (.A1(_0373_),
    .A2(_1158_),
    .Z(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2118_ (.A1(_1097_),
    .A2(_1164_),
    .B(_1165_),
    .ZN(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2119_ (.A1(_1163_),
    .A2(_1166_),
    .Z(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2120_ (.A1(_1162_),
    .A2(_1167_),
    .ZN(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2121_ (.A1(_1162_),
    .A2(_1167_),
    .ZN(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2122_ (.A1(_1153_),
    .A2(_1168_),
    .B(_1169_),
    .ZN(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _2123_ (.I(_1119_),
    .Z(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _2124_ (.A1(_0962_),
    .A2(_1171_),
    .ZN(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2125_ (.A1(_0996_),
    .A2(_1119_),
    .ZN(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2126_ (.A1(_1132_),
    .A2(_1133_),
    .B(_1173_),
    .ZN(_1174_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _2127_ (.A1(_0395_),
    .A2(_1016_),
    .Z(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2128_ (.A1(_1122_),
    .A2(_1125_),
    .Z(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2129_ (.A1(_1175_),
    .A2(_1131_),
    .B1(_1176_),
    .B2(_1035_),
    .ZN(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2130_ (.A1(_1120_),
    .A2(_1177_),
    .Z(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2131_ (.A1(_1174_),
    .A2(_1178_),
    .Z(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2132_ (.A1(_1172_),
    .A2(_1179_),
    .Z(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2133_ (.A1(_1170_),
    .A2(_1180_),
    .ZN(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2134_ (.A1(_1170_),
    .A2(_1180_),
    .ZN(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2135_ (.A1(_1138_),
    .A2(_1181_),
    .B(_1182_),
    .ZN(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _2136_ (.A1(_0792_),
    .A2(_0793_),
    .B(_1158_),
    .ZN(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2137_ (.A1(_1184_),
    .A2(_1160_),
    .Z(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2138_ (.A1(_1115_),
    .A2(\sigRom.address[0] ),
    .ZN(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_4 _2139_ (.A1(_1118_),
    .A2(_1186_),
    .Z(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _2140_ (.A1(_1115_),
    .A2(_1117_),
    .Z(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _2141_ (.A1(_1147_),
    .A2(_1188_),
    .Z(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2142_ (.A1(_0911_),
    .A2(_0912_),
    .ZN(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2143_ (.A1(_1115_),
    .A2(_1117_),
    .ZN(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2144_ (.A1(\sigRom.address[0] ),
    .A2(_1191_),
    .B(_1123_),
    .ZN(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _2145_ (.A1(_1122_),
    .A2(_1192_),
    .Z(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2146_ (.A1(_0879_),
    .A2(_0880_),
    .ZN(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _2147_ (.A1(_0900_),
    .A2(_1187_),
    .B1(_1189_),
    .B2(_1190_),
    .C1(_1193_),
    .C2(_1194_),
    .ZN(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2148_ (.A1(_1185_),
    .A2(_1195_),
    .ZN(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2149_ (.I(_1158_),
    .Z(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2150_ (.A1(_0812_),
    .A2(_1197_),
    .ZN(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2151_ (.A1(_0945_),
    .A2(_1184_),
    .ZN(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2152_ (.A1(_0794_),
    .A2(_0836_),
    .B(_1197_),
    .ZN(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2153_ (.A1(_1199_),
    .A2(_1200_),
    .ZN(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _2154_ (.A1(_0884_),
    .A2(_1187_),
    .B1(_1189_),
    .B2(_0900_),
    .C1(_1193_),
    .C2(_1154_),
    .ZN(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2155_ (.A1(_1198_),
    .A2(_1201_),
    .A3(_1202_),
    .Z(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2156_ (.A1(_1196_),
    .A2(_1203_),
    .ZN(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2157_ (.A1(_1152_),
    .A2(_1168_),
    .Z(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2158_ (.A1(_1196_),
    .A2(_1203_),
    .ZN(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2159_ (.A1(_1204_),
    .A2(_1205_),
    .B(_1206_),
    .ZN(_1207_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2160_ (.A1(_1198_),
    .A2(_1199_),
    .A3(_1200_),
    .Z(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2161_ (.A1(_1199_),
    .A2(_1200_),
    .B(_1198_),
    .ZN(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2162_ (.A1(_1208_),
    .A2(_1209_),
    .A3(_1202_),
    .ZN(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2163_ (.A1(_0318_),
    .A2(_1158_),
    .ZN(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2164_ (.A1(_0810_),
    .A2(_0811_),
    .Z(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2165_ (.A1(_0810_),
    .A2(_0811_),
    .B(_1141_),
    .ZN(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _2166_ (.A1(_0848_),
    .A2(_1158_),
    .Z(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2167_ (.I0(_1212_),
    .I1(_1213_),
    .S(_1214_),
    .Z(_1215_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2168_ (.A1(_1211_),
    .A2(_1215_),
    .Z(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _2169_ (.A1(_1194_),
    .A2(_1187_),
    .B1(_1193_),
    .B2(_0945_),
    .C1(_1189_),
    .C2(_0884_),
    .ZN(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2170_ (.A1(_1216_),
    .A2(_1217_),
    .Z(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2171_ (.A1(_1210_),
    .A2(_1218_),
    .ZN(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2172_ (.A1(_1163_),
    .A2(_1166_),
    .ZN(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2173_ (.A1(_0945_),
    .A2(_1142_),
    .B(_1184_),
    .ZN(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2174_ (.A1(_1213_),
    .A2(_1221_),
    .B(_1199_),
    .ZN(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2175_ (.A1(_1067_),
    .A2(_1150_),
    .ZN(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2176_ (.A1(_0472_),
    .A2(_1197_),
    .Z(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2177_ (.A1(_1056_),
    .A2(_1164_),
    .B(_1224_),
    .ZN(_1225_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2178_ (.A1(_1223_),
    .A2(_1225_),
    .Z(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2179_ (.A1(_1220_),
    .A2(_1222_),
    .A3(_1226_),
    .Z(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2180_ (.A1(_1219_),
    .A2(_1227_),
    .Z(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2181_ (.A1(_1207_),
    .A2(_1228_),
    .Z(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2182_ (.A1(_1138_),
    .A2(_1181_),
    .Z(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2183_ (.A1(_1207_),
    .A2(_1228_),
    .Z(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2184_ (.A1(_1229_),
    .A2(_1230_),
    .B(_1231_),
    .ZN(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2185_ (.A1(_1210_),
    .A2(_1218_),
    .ZN(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2186_ (.A1(_1219_),
    .A2(_1227_),
    .B(_1233_),
    .ZN(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2187_ (.A1(_1216_),
    .A2(_1217_),
    .ZN(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2188_ (.A1(_1223_),
    .A2(_1225_),
    .Z(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2189_ (.A1(_0848_),
    .A2(_1197_),
    .ZN(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2190_ (.A1(_1213_),
    .A2(_1214_),
    .ZN(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2191_ (.A1(_1212_),
    .A2(_1237_),
    .B1(_1238_),
    .B2(_1211_),
    .ZN(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2192_ (.A1(_1045_),
    .A2(_1150_),
    .ZN(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2193_ (.A1(_0406_),
    .A2(_1141_),
    .ZN(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2194_ (.A1(_1067_),
    .A2(_1164_),
    .B(_1241_),
    .ZN(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2195_ (.A1(_1240_),
    .A2(_1242_),
    .ZN(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2196_ (.A1(_1239_),
    .A2(_1243_),
    .ZN(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2197_ (.A1(_1236_),
    .A2(_1244_),
    .Z(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2198_ (.A1(_0747_),
    .A2(_0748_),
    .A3(_1197_),
    .ZN(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2199_ (.A1(_1139_),
    .A2(_1246_),
    .ZN(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2200_ (.I(_1197_),
    .Z(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2201_ (.A1(_0318_),
    .A2(_0749_),
    .B(_1248_),
    .ZN(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2202_ (.A1(_1247_),
    .A2(_1249_),
    .Z(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2203_ (.A1(_1122_),
    .A2(_1192_),
    .ZN(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _2204_ (.I(_1251_),
    .Z(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2205_ (.A1(_0848_),
    .A2(_1252_),
    .ZN(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2206_ (.A1(_1154_),
    .A2(_1187_),
    .B1(_1189_),
    .B2(_1194_),
    .C(_1253_),
    .ZN(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2207_ (.A1(_1165_),
    .A2(_1250_),
    .A3(_1254_),
    .Z(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _2208_ (.A1(_1235_),
    .A2(_1245_),
    .A3(_1255_),
    .ZN(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2209_ (.A1(_1234_),
    .A2(_1256_),
    .Z(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2210_ (.A1(_1174_),
    .A2(_1178_),
    .ZN(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2211_ (.A1(_1172_),
    .A2(_1179_),
    .B(_1258_),
    .ZN(_1259_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2212_ (.A1(_1222_),
    .A2(_1226_),
    .ZN(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2213_ (.A1(_1222_),
    .A2(_1226_),
    .ZN(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2214_ (.A1(_1220_),
    .A2(_1260_),
    .B(_1261_),
    .ZN(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2215_ (.A1(_0965_),
    .A2(_1171_),
    .ZN(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _2216_ (.A1(_0962_),
    .A2(_1119_),
    .Z(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2217_ (.A1(_0985_),
    .A2(_1119_),
    .Z(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2218_ (.A1(_1265_),
    .A2(_1177_),
    .Z(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _2219_ (.A1(_1025_),
    .A2(_1119_),
    .Z(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2220_ (.A1(_1017_),
    .A2(_1126_),
    .B(_1267_),
    .ZN(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2221_ (.A1(_1264_),
    .A2(_1266_),
    .A3(_1268_),
    .Z(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2222_ (.A1(_1263_),
    .A2(_1269_),
    .Z(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2223_ (.A1(_1262_),
    .A2(_1270_),
    .ZN(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2224_ (.A1(_1259_),
    .A2(_1271_),
    .Z(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2225_ (.A1(_1257_),
    .A2(_1272_),
    .ZN(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2226_ (.A1(_1232_),
    .A2(_1273_),
    .Z(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2227_ (.A1(_1232_),
    .A2(_1273_),
    .ZN(_1275_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2228_ (.A1(_1183_),
    .A2(_1274_),
    .B(_1275_),
    .ZN(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2229_ (.A1(_1262_),
    .A2(_1270_),
    .ZN(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2230_ (.A1(_1259_),
    .A2(_1271_),
    .B(_1277_),
    .ZN(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2231_ (.A1(_1234_),
    .A2(_1256_),
    .Z(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2232_ (.A1(_1257_),
    .A2(_1272_),
    .B(_1279_),
    .ZN(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2233_ (.A1(_1264_),
    .A2(_1268_),
    .Z(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2234_ (.A1(_1266_),
    .A2(_1281_),
    .ZN(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2235_ (.A1(_1263_),
    .A2(_1269_),
    .B(_1282_),
    .ZN(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2236_ (.I(_1236_),
    .ZN(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2237_ (.A1(_1239_),
    .A2(_1243_),
    .Z(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2238_ (.A1(_1284_),
    .A2(_1244_),
    .B(_1285_),
    .ZN(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2239_ (.A1(_1172_),
    .A2(_1268_),
    .ZN(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2240_ (.A1(_0955_),
    .A2(_0968_),
    .Z(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2241_ (.I(_1131_),
    .Z(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2242_ (.A1(_1288_),
    .A2(_1289_),
    .ZN(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _2243_ (.A1(_0965_),
    .A2(_1007_),
    .A3(_1171_),
    .Z(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2244_ (.A1(_1121_),
    .A2(_1263_),
    .B(_1291_),
    .ZN(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _2245_ (.A1(_1287_),
    .A2(_1290_),
    .A3(_1292_),
    .ZN(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2246_ (.A1(_1286_),
    .A2(_1293_),
    .ZN(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2247_ (.A1(_1283_),
    .A2(_1294_),
    .Z(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2248_ (.A1(_1235_),
    .A2(_1255_),
    .ZN(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2249_ (.A1(_1235_),
    .A2(_1255_),
    .ZN(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2250_ (.A1(_1245_),
    .A2(_1296_),
    .B(_1297_),
    .ZN(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2251_ (.A1(_1240_),
    .A2(_1242_),
    .ZN(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2252_ (.A1(_0747_),
    .A2(_0748_),
    .ZN(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2253_ (.A1(_1139_),
    .A2(_1300_),
    .B(_1142_),
    .ZN(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2254_ (.A1(_1165_),
    .A2(_1301_),
    .B(_1247_),
    .ZN(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2255_ (.A1(_1148_),
    .A2(_1149_),
    .Z(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2256_ (.I(_1164_),
    .Z(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2257_ (.I(_1126_),
    .Z(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2258_ (.A1(_1045_),
    .A2(_1304_),
    .B1(_1305_),
    .B2(_1025_),
    .ZN(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2259_ (.A1(_1035_),
    .A2(_1303_),
    .B(_1306_),
    .ZN(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2260_ (.A1(_1302_),
    .A2(_1307_),
    .Z(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2261_ (.A1(_1299_),
    .A2(_1308_),
    .Z(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2262_ (.A1(_0373_),
    .A2(_1197_),
    .ZN(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2263_ (.A1(_1310_),
    .A2(_1247_),
    .A3(_1249_),
    .Z(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2264_ (.A1(_1247_),
    .A2(_1249_),
    .B(_1310_),
    .ZN(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2265_ (.A1(_1311_),
    .A2(_1312_),
    .A3(_1254_),
    .ZN(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2266_ (.A1(_0472_),
    .A2(_1197_),
    .ZN(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2267_ (.I0(_0373_),
    .I1(_1310_),
    .S(_1156_),
    .Z(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2268_ (.A1(_1314_),
    .A2(_1315_),
    .Z(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_4 _2269_ (.A1(_1123_),
    .A2(_1186_),
    .Z(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _2270_ (.A1(_1147_),
    .A2(_1188_),
    .ZN(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_4 _2271_ (.A1(_0836_),
    .A2(_1317_),
    .B1(_1318_),
    .B2(_0943_),
    .C1(_0749_),
    .C2(_1252_),
    .ZN(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2272_ (.A1(_1316_),
    .A2(_1319_),
    .Z(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2273_ (.A1(_1313_),
    .A2(_1320_),
    .Z(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2274_ (.A1(_1309_),
    .A2(_1321_),
    .Z(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2275_ (.A1(_1298_),
    .A2(_1322_),
    .Z(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2276_ (.A1(_1295_),
    .A2(_1324_),
    .ZN(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _2277_ (.A1(_1278_),
    .A2(_1280_),
    .A3(_1325_),
    .ZN(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2278_ (.A1(_1276_),
    .A2(_1326_),
    .ZN(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2279_ (.A1(_1286_),
    .A2(_1293_),
    .ZN(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2280_ (.A1(_1283_),
    .A2(_1294_),
    .B(_1328_),
    .ZN(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2281_ (.A1(_1298_),
    .A2(_1322_),
    .ZN(_1330_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2282_ (.A1(_1295_),
    .A2(_1324_),
    .ZN(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2283_ (.A1(_1330_),
    .A2(_1331_),
    .ZN(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2284_ (.A1(_1290_),
    .A2(_1292_),
    .Z(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2285_ (.A1(_1172_),
    .A2(_1268_),
    .A3(_1333_),
    .ZN(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2286_ (.I(_1307_),
    .ZN(_1336_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2287_ (.A1(_1302_),
    .A2(_1336_),
    .ZN(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2288_ (.A1(_1299_),
    .A2(_1308_),
    .B(_1337_),
    .ZN(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2289_ (.A1(_1290_),
    .A2(_1292_),
    .B(_1291_),
    .ZN(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _2290_ (.A1(_0972_),
    .A2(_1171_),
    .Z(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2291_ (.A1(_1129_),
    .A2(_1290_),
    .Z(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2292_ (.A1(_1288_),
    .A2(_1173_),
    .B(_1341_),
    .ZN(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2293_ (.A1(_1340_),
    .A2(_1342_),
    .ZN(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2294_ (.A1(_1339_),
    .A2(_1343_),
    .Z(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2295_ (.A1(_1338_),
    .A2(_1344_),
    .ZN(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2296_ (.A1(_1335_),
    .A2(_1346_),
    .Z(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2297_ (.A1(_1313_),
    .A2(_1320_),
    .ZN(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2298_ (.A1(_1309_),
    .A2(_1321_),
    .ZN(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2299_ (.A1(_1348_),
    .A2(_1349_),
    .ZN(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2300_ (.A1(_1157_),
    .A2(_1310_),
    .B1(_1314_),
    .B2(_1315_),
    .ZN(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2301_ (.A1(_1007_),
    .A2(_1305_),
    .ZN(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _2302_ (.A1(_1175_),
    .A2(_1303_),
    .B1(_1145_),
    .B2(_1035_),
    .C(_1352_),
    .ZN(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2303_ (.A1(_1351_),
    .A2(_1353_),
    .ZN(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2304_ (.A1(_1316_),
    .A2(_1319_),
    .ZN(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2305_ (.A1(_1378_),
    .A2(_1248_),
    .ZN(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2306_ (.I0(_1314_),
    .I1(_0472_),
    .S(_1184_),
    .Z(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2307_ (.A1(_1357_),
    .A2(_1358_),
    .Z(_1359_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_4 _2308_ (.A1(_0848_),
    .A2(_1317_),
    .B1(_1318_),
    .B2(_0836_),
    .C1(_0770_),
    .C2(_1252_),
    .ZN(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2309_ (.A1(_1359_),
    .A2(_1360_),
    .ZN(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2310_ (.A1(_1355_),
    .A2(_1361_),
    .Z(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2311_ (.A1(_1355_),
    .A2(_1361_),
    .ZN(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2312_ (.A1(_1362_),
    .A2(_1363_),
    .ZN(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2313_ (.A1(_1354_),
    .A2(_1364_),
    .Z(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2314_ (.A1(_1350_),
    .A2(_1365_),
    .Z(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2315_ (.A1(_1347_),
    .A2(_1366_),
    .Z(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2316_ (.A1(_1332_),
    .A2(_1368_),
    .Z(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2317_ (.A1(_1329_),
    .A2(_1369_),
    .ZN(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2318_ (.A1(_1280_),
    .A2(_1325_),
    .ZN(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2319_ (.A1(_1280_),
    .A2(_1325_),
    .ZN(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2320_ (.A1(_1278_),
    .A2(_1371_),
    .B(_1372_),
    .ZN(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2321_ (.A1(_1370_),
    .A2(_1373_),
    .Z(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2322_ (.A1(_1327_),
    .A2(_1374_),
    .Z(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2323_ (.A1(_1276_),
    .A2(_1326_),
    .Z(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2324_ (.A1(_1025_),
    .A2(_1171_),
    .ZN(_1377_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _2325_ (.A1(_1065_),
    .A2(_1066_),
    .A3(_1289_),
    .ZN(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2326_ (.A1(_1056_),
    .A2(_1305_),
    .B(_1379_),
    .ZN(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2327_ (.A1(_1377_),
    .A2(_1380_),
    .ZN(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2328_ (.A1(_1121_),
    .A2(_1127_),
    .ZN(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2329_ (.A1(_1121_),
    .A2(_1127_),
    .A3(_1381_),
    .Z(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2330_ (.A1(_1128_),
    .A2(_1381_),
    .A3(_1382_),
    .B1(_1383_),
    .B2(_1129_),
    .ZN(_1384_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _2331_ (.A1(_0879_),
    .A2(_0880_),
    .B(_1197_),
    .ZN(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2332_ (.I0(_1246_),
    .I1(_0749_),
    .S(_1385_),
    .Z(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2333_ (.A1(_0770_),
    .A2(_1248_),
    .ZN(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2334_ (.A1(_1300_),
    .A2(_1385_),
    .B1(_1386_),
    .B2(_1387_),
    .ZN(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2335_ (.A1(_1097_),
    .A2(_1150_),
    .ZN(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2336_ (.A1(_1143_),
    .A2(_1146_),
    .ZN(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2337_ (.A1(_1390_),
    .A2(_1391_),
    .ZN(_1392_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2338_ (.A1(_1390_),
    .A2(_1391_),
    .A3(_1388_),
    .Z(_1393_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2339_ (.A1(_1088_),
    .A2(_1164_),
    .B(_1213_),
    .ZN(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2340_ (.A1(_1078_),
    .A2(_1303_),
    .A3(_1394_),
    .ZN(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2341_ (.A1(_1152_),
    .A2(_1388_),
    .A3(_1392_),
    .B1(_1393_),
    .B2(_1395_),
    .ZN(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2342_ (.A1(_1120_),
    .A2(_1136_),
    .Z(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2343_ (.A1(_1396_),
    .A2(_1397_),
    .Z(_1398_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2344_ (.A1(_1396_),
    .A2(_1397_),
    .Z(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2345_ (.A1(_1384_),
    .A2(_1398_),
    .B(_1399_),
    .ZN(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2346_ (.A1(_0884_),
    .A2(_1142_),
    .ZN(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _2347_ (.A1(_1367_),
    .A2(_0925_),
    .Z(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2348_ (.A1(_1403_),
    .A2(_1187_),
    .B1(_1193_),
    .B2(_0900_),
    .ZN(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _2349_ (.A1(_1190_),
    .A2(_1187_),
    .B1(_1189_),
    .B2(_1403_),
    .C1(_1193_),
    .C2(_0884_),
    .ZN(_1405_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2350_ (.A1(_1402_),
    .A2(_1404_),
    .B(_1405_),
    .ZN(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2351_ (.A1(_1387_),
    .A2(_1386_),
    .Z(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2352_ (.A1(_1402_),
    .A2(_1404_),
    .A3(_1405_),
    .ZN(_1408_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2353_ (.A1(_1406_),
    .A2(_1407_),
    .B(_1408_),
    .ZN(_1409_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2354_ (.A1(_1185_),
    .A2(_1195_),
    .ZN(_1410_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2355_ (.A1(_1409_),
    .A2(_1410_),
    .ZN(_1412_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2356_ (.A1(_1395_),
    .A2(_1393_),
    .Z(_1413_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2357_ (.A1(_1409_),
    .A2(_1410_),
    .ZN(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2358_ (.A1(_1412_),
    .A2(_1413_),
    .B(_1414_),
    .ZN(_1415_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2359_ (.A1(_1204_),
    .A2(_1205_),
    .ZN(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2360_ (.A1(_1415_),
    .A2(_1416_),
    .ZN(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _2361_ (.A1(_1384_),
    .A2(_1396_),
    .A3(_1397_),
    .ZN(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2362_ (.A1(_1415_),
    .A2(_1416_),
    .Z(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2363_ (.A1(_1417_),
    .A2(_1418_),
    .B(_1419_),
    .ZN(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2364_ (.A1(_1229_),
    .A2(_1230_),
    .Z(_1421_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2365_ (.A1(_1420_),
    .A2(_1421_),
    .ZN(_1423_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2366_ (.A1(_1420_),
    .A2(_1421_),
    .ZN(_1424_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2367_ (.A1(_1401_),
    .A2(_1423_),
    .B(_1424_),
    .ZN(_1425_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2368_ (.A1(_1183_),
    .A2(_1274_),
    .Z(_1426_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2369_ (.A1(_1425_),
    .A2(_1426_),
    .ZN(_1427_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2370_ (.A1(_1425_),
    .A2(_1426_),
    .ZN(_1428_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2371_ (.A1(_1340_),
    .A2(_1427_),
    .B(_1428_),
    .ZN(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2372_ (.A1(_1376_),
    .A2(_1429_),
    .Z(_1430_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2373_ (.A1(_1375_),
    .A2(_1430_),
    .ZN(_1431_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _2374_ (.A1(_1056_),
    .A2(_1171_),
    .Z(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2375_ (.A1(_0955_),
    .A2(_1087_),
    .Z(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _2376_ (.A1(_0395_),
    .A2(_1096_),
    .Z(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2377_ (.A1(_1434_),
    .A2(_1303_),
    .B1(_1176_),
    .B2(_1435_),
    .ZN(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2378_ (.I0(_0749_),
    .I1(_1246_),
    .S(_1214_),
    .Z(_1437_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2379_ (.A1(_1300_),
    .A2(_1237_),
    .B1(_1437_),
    .B2(_1184_),
    .ZN(_1438_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2380_ (.A1(_1077_),
    .A2(_1303_),
    .ZN(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2381_ (.A1(_1439_),
    .A2(_1394_),
    .Z(_1440_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2382_ (.A1(_1438_),
    .A2(_1440_),
    .ZN(_1441_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2383_ (.A1(_1432_),
    .A2(_1436_),
    .A3(_1441_),
    .B1(_1440_),
    .B2(_1438_),
    .ZN(_1442_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2384_ (.A1(_1129_),
    .A2(_1383_),
    .Z(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2385_ (.A1(_1017_),
    .A2(_1171_),
    .ZN(_1445_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2386_ (.I0(_1017_),
    .I1(_1445_),
    .S(_1267_),
    .Z(_1446_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2387_ (.A1(_1175_),
    .A2(_1377_),
    .B1(_1446_),
    .B2(_1173_),
    .ZN(_1447_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2388_ (.A1(_1267_),
    .A2(_1380_),
    .Z(_1448_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2389_ (.A1(_1447_),
    .A2(_1448_),
    .ZN(_1449_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2390_ (.A1(_1447_),
    .A2(_1448_),
    .ZN(_1450_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2391_ (.A1(_1121_),
    .A2(_1449_),
    .B(_1450_),
    .ZN(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2392_ (.A1(_1442_),
    .A2(_1443_),
    .ZN(_1452_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2393_ (.A1(_1451_),
    .A2(_1452_),
    .ZN(_1453_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2394_ (.A1(_1442_),
    .A2(_1443_),
    .B(_1453_),
    .ZN(_1454_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2395_ (.A1(_1402_),
    .A2(_1404_),
    .ZN(_1456_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2396_ (.A1(_0911_),
    .A2(_0912_),
    .B(_1251_),
    .ZN(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _2397_ (.A1(_0900_),
    .A2(_1457_),
    .B(_1142_),
    .C(_0945_),
    .ZN(_1458_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2398_ (.A1(_1402_),
    .A2(_1404_),
    .Z(_1459_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2399_ (.A1(_1402_),
    .A2(_1404_),
    .A3(_1458_),
    .Z(_1460_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2400_ (.A1(_1161_),
    .A2(_1437_),
    .Z(_1461_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2401_ (.A1(_1456_),
    .A2(_1458_),
    .A3(_1459_),
    .B1(_1460_),
    .B2(_1461_),
    .ZN(_1462_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _2402_ (.A1(_1456_),
    .A2(_1405_),
    .A3(_1407_),
    .ZN(_1463_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2403_ (.A1(_1462_),
    .A2(_1463_),
    .Z(_1464_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2404_ (.A1(_1432_),
    .A2(_1436_),
    .ZN(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2405_ (.A1(_1465_),
    .A2(_1441_),
    .ZN(_1467_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2406_ (.A1(_1462_),
    .A2(_1463_),
    .Z(_1468_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2407_ (.A1(_1464_),
    .A2(_1467_),
    .B(_1468_),
    .ZN(_1469_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _2408_ (.A1(_1409_),
    .A2(_1410_),
    .A3(_1413_),
    .ZN(_1470_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2409_ (.A1(_1469_),
    .A2(_1470_),
    .Z(_1471_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2410_ (.A1(_1451_),
    .A2(_1452_),
    .Z(_1472_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2411_ (.A1(_1469_),
    .A2(_1470_),
    .ZN(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2412_ (.A1(_1471_),
    .A2(_1472_),
    .B(_1473_),
    .ZN(_1474_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2413_ (.A1(_1417_),
    .A2(_1418_),
    .ZN(_1475_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2414_ (.A1(_1474_),
    .A2(_1475_),
    .ZN(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2415_ (.A1(_1474_),
    .A2(_1475_),
    .Z(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2416_ (.A1(_1454_),
    .A2(_1476_),
    .B(_1478_),
    .ZN(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2417_ (.A1(_1401_),
    .A2(_1423_),
    .Z(_1480_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2418_ (.A1(_1479_),
    .A2(_1480_),
    .ZN(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2419_ (.A1(_1479_),
    .A2(_1480_),
    .ZN(_1482_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2420_ (.A1(_1290_),
    .A2(_1481_),
    .B(_1482_),
    .ZN(_1483_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2421_ (.A1(_1340_),
    .A2(_1427_),
    .Z(_1484_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2422_ (.A1(_1483_),
    .A2(_1484_),
    .ZN(_1485_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2423_ (.A1(_1290_),
    .A2(_1481_),
    .Z(_1486_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2424_ (.A1(_1435_),
    .A2(_1035_),
    .A3(_1289_),
    .ZN(_1487_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2425_ (.A1(_1097_),
    .A2(_1171_),
    .ZN(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2426_ (.A1(_1132_),
    .A2(_1489_),
    .B(_1487_),
    .C(_1445_),
    .ZN(_1490_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2427_ (.A1(_1487_),
    .A2(_1490_),
    .Z(_1491_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2428_ (.A1(_0770_),
    .A2(_1214_),
    .ZN(_1492_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2429_ (.A1(_1432_),
    .A2(_1436_),
    .Z(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2430_ (.A1(_1492_),
    .A2(_1493_),
    .Z(_1494_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2431_ (.I(_1494_),
    .ZN(_1495_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2432_ (.A1(_1492_),
    .A2(_1493_),
    .ZN(_1496_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2433_ (.A1(_1491_),
    .A2(_1495_),
    .B(_1496_),
    .ZN(_1497_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2434_ (.A1(_1121_),
    .A2(_1447_),
    .A3(_1448_),
    .Z(_1498_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2435_ (.A1(_1497_),
    .A2(_1498_),
    .ZN(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2436_ (.A1(_1497_),
    .A2(_1498_),
    .Z(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2437_ (.A1(_1157_),
    .A2(_1237_),
    .ZN(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2438_ (.A1(_1156_),
    .A2(_1214_),
    .ZN(_1503_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2439_ (.A1(_1078_),
    .A2(_1176_),
    .B1(_1502_),
    .B2(_1503_),
    .ZN(_1504_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _2440_ (.A1(_0913_),
    .A2(_1248_),
    .B1(_1252_),
    .B2(_0926_),
    .ZN(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _2441_ (.A1(_0898_),
    .A2(_0899_),
    .A3(_1142_),
    .ZN(_1506_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _2442_ (.A1(_0836_),
    .A2(_1248_),
    .B1(_1252_),
    .B2(_0913_),
    .C(_1506_),
    .ZN(_1507_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2443_ (.A1(_1159_),
    .A2(_1505_),
    .B1(_1507_),
    .B2(_1458_),
    .ZN(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2444_ (.A1(_1159_),
    .A2(_1458_),
    .A3(_1505_),
    .A4(_1507_),
    .ZN(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2445_ (.A1(_1504_),
    .A2(_1508_),
    .B(_1509_),
    .ZN(_1511_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2446_ (.A1(_1460_),
    .A2(_1461_),
    .Z(_1512_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2447_ (.A1(_1511_),
    .A2(_1512_),
    .ZN(_1513_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2448_ (.A1(_1491_),
    .A2(_1494_),
    .Z(_1514_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2449_ (.A1(_1511_),
    .A2(_1512_),
    .ZN(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2450_ (.A1(_1513_),
    .A2(_1514_),
    .B(_1515_),
    .ZN(_1516_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2451_ (.A1(_1464_),
    .A2(_1467_),
    .Z(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2452_ (.A1(_1516_),
    .A2(_1517_),
    .Z(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2453_ (.A1(_1516_),
    .A2(_1517_),
    .Z(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2454_ (.A1(_1501_),
    .A2(_1518_),
    .B(_1519_),
    .ZN(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2455_ (.A1(_1471_),
    .A2(_1472_),
    .ZN(_1522_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2456_ (.A1(_1520_),
    .A2(_1522_),
    .ZN(_1523_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2457_ (.A1(_1520_),
    .A2(_1522_),
    .Z(_1524_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2458_ (.A1(_1500_),
    .A2(_1523_),
    .B(_1524_),
    .ZN(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2459_ (.A1(_1454_),
    .A2(_1476_),
    .Z(_1526_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2460_ (.A1(_1525_),
    .A2(_1526_),
    .ZN(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2461_ (.A1(_1525_),
    .A2(_1526_),
    .ZN(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _2462_ (.A1(_0965_),
    .A2(_1171_),
    .A3(_1527_),
    .B(_1528_),
    .ZN(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2463_ (.A1(_1483_),
    .A2(_1484_),
    .B1(_1486_),
    .B2(_1529_),
    .ZN(_1530_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2464_ (.A1(_1485_),
    .A2(_1530_),
    .Z(_1531_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2465_ (.A1(_1431_),
    .A2(_1531_),
    .Z(_1533_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2466_ (.A1(_1045_),
    .A2(_1171_),
    .ZN(_1534_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2467_ (.I(_1534_),
    .ZN(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2468_ (.A1(_1077_),
    .A2(_1289_),
    .ZN(_1536_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2469_ (.A1(_1535_),
    .A2(_1536_),
    .ZN(_1537_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2470_ (.A1(_1078_),
    .A2(_1534_),
    .B1(_1132_),
    .B2(_1537_),
    .ZN(_1538_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2471_ (.A1(_0945_),
    .A2(_1142_),
    .ZN(_1539_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2472_ (.A1(_0749_),
    .A2(_1539_),
    .ZN(_1540_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2473_ (.A1(_1175_),
    .A2(_1289_),
    .ZN(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2474_ (.A1(_1132_),
    .A2(_1489_),
    .B(_1487_),
    .ZN(_1542_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2475_ (.A1(_1541_),
    .A2(_1542_),
    .Z(_1544_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2476_ (.A1(_1540_),
    .A2(_1544_),
    .ZN(_1545_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2477_ (.A1(_1540_),
    .A2(_1544_),
    .ZN(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2478_ (.A1(_1538_),
    .A2(_1545_),
    .B(_1546_),
    .ZN(_1547_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2479_ (.A1(_1173_),
    .A2(_1446_),
    .Z(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2480_ (.A1(_1547_),
    .A2(_1548_),
    .ZN(_1549_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2481_ (.A1(_1547_),
    .A2(_1548_),
    .Z(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2482_ (.I(_1550_),
    .ZN(_1551_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2483_ (.A1(_0836_),
    .A2(_1248_),
    .ZN(_1552_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2484_ (.A1(_1552_),
    .A2(_1246_),
    .ZN(_1553_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2485_ (.A1(_1088_),
    .A2(_1305_),
    .B1(_1540_),
    .B2(_1553_),
    .ZN(_1555_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2486_ (.A1(_0926_),
    .A2(_1248_),
    .ZN(_1556_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2487_ (.A1(_0926_),
    .A2(_0881_),
    .B(_1248_),
    .ZN(_1557_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2488_ (.A1(_1194_),
    .A2(_1556_),
    .B1(_1557_),
    .B2(_1159_),
    .ZN(_1558_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2489_ (.A1(_1155_),
    .A2(_1505_),
    .Z(_1559_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2490_ (.A1(_1558_),
    .A2(_1559_),
    .Z(_1560_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2491_ (.A1(_1558_),
    .A2(_1559_),
    .ZN(_1561_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2492_ (.A1(_1555_),
    .A2(_1560_),
    .B(_1561_),
    .ZN(_1562_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2493_ (.A1(_1159_),
    .A2(_1505_),
    .ZN(_1563_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2494_ (.A1(_1458_),
    .A2(_1507_),
    .ZN(_1564_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2495_ (.A1(_1563_),
    .A2(_1564_),
    .A3(_1504_),
    .Z(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2496_ (.A1(_1562_),
    .A2(_1566_),
    .ZN(_1567_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2497_ (.A1(_1538_),
    .A2(_1545_),
    .ZN(_1568_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2498_ (.A1(_1562_),
    .A2(_1566_),
    .Z(_1569_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2499_ (.A1(_1567_),
    .A2(_1568_),
    .B(_1569_),
    .ZN(_1570_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _2500_ (.A1(_1511_),
    .A2(_1512_),
    .A3(_1514_),
    .ZN(_1571_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2501_ (.A1(_1570_),
    .A2(_1571_),
    .ZN(_1572_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2502_ (.A1(_1570_),
    .A2(_1571_),
    .ZN(_1573_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2503_ (.A1(_1551_),
    .A2(_1572_),
    .B(_1573_),
    .ZN(_1574_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2504_ (.A1(_1501_),
    .A2(_1518_),
    .Z(_1575_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2505_ (.A1(_1574_),
    .A2(_1575_),
    .ZN(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2506_ (.A1(_1574_),
    .A2(_1575_),
    .ZN(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2507_ (.A1(_1549_),
    .A2(_1577_),
    .B(_1578_),
    .ZN(_1579_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _2508_ (.A1(_1500_),
    .A2(_1523_),
    .Z(_1580_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2509_ (.A1(_1579_),
    .A2(_1580_),
    .Z(_1581_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2510_ (.A1(_1579_),
    .A2(_1580_),
    .Z(_1582_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2511_ (.A1(_1263_),
    .A2(_1525_),
    .A3(_1526_),
    .Z(_1583_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _2512_ (.A1(_1172_),
    .A2(_1581_),
    .B(_1582_),
    .C(_1583_),
    .ZN(_1584_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2513_ (.A1(_1579_),
    .A2(_1580_),
    .ZN(_1585_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2514_ (.A1(_1579_),
    .A2(_1580_),
    .ZN(_1586_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2515_ (.A1(_1264_),
    .A2(_1585_),
    .B(_1586_),
    .ZN(_1588_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2516_ (.A1(_1434_),
    .A2(_1237_),
    .A3(_1289_),
    .ZN(_1589_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2517_ (.A1(_1434_),
    .A2(_1289_),
    .ZN(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2518_ (.A1(_1237_),
    .A2(_1590_),
    .Z(_1591_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2519_ (.A1(_1379_),
    .A2(_1591_),
    .Z(_1592_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2520_ (.I0(_1536_),
    .I1(_1078_),
    .S(_1534_),
    .Z(_1593_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2521_ (.A1(_1132_),
    .A2(_1593_),
    .Z(_1594_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2522_ (.A1(_1589_),
    .A2(_1592_),
    .B(_1594_),
    .ZN(_1595_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2523_ (.A1(_1045_),
    .A2(_1541_),
    .ZN(_1596_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2524_ (.I(_1596_),
    .ZN(_1597_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2525_ (.A1(_1379_),
    .A2(_1591_),
    .B(_1589_),
    .ZN(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2526_ (.A1(_0033_),
    .A2(_1594_),
    .Z(_0034_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2527_ (.A1(_1597_),
    .A2(_0034_),
    .ZN(_0035_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2528_ (.A1(_1595_),
    .A2(_0035_),
    .B(_1121_),
    .ZN(_0036_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2529_ (.A1(_1595_),
    .A2(_0035_),
    .ZN(_0037_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2530_ (.A1(_1121_),
    .A2(_0037_),
    .ZN(_0038_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2531_ (.A1(_1403_),
    .A2(_1385_),
    .ZN(_0039_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2532_ (.A1(_1159_),
    .A2(_0039_),
    .A3(_1557_),
    .Z(_0040_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2533_ (.A1(_0039_),
    .A2(_1557_),
    .B(_1159_),
    .ZN(_0041_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2534_ (.A1(_0863_),
    .A2(_0864_),
    .B(_1197_),
    .ZN(_0042_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2535_ (.I0(_1385_),
    .I1(_0881_),
    .S(_0042_),
    .Z(_0044_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2536_ (.A1(_1194_),
    .A2(_0042_),
    .B1(_0044_),
    .B2(_1552_),
    .ZN(_0045_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2537_ (.A1(_0040_),
    .A2(_0041_),
    .B(_0045_),
    .ZN(_0046_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2538_ (.A1(_1379_),
    .A2(_1591_),
    .Z(_0047_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2539_ (.A1(_0040_),
    .A2(_0045_),
    .A3(_0041_),
    .ZN(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2540_ (.A1(_0046_),
    .A2(_0047_),
    .B(_0048_),
    .ZN(_0049_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2541_ (.A1(_1555_),
    .A2(_1560_),
    .ZN(_0050_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2542_ (.A1(_0049_),
    .A2(_0050_),
    .ZN(_0051_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2543_ (.A1(_1597_),
    .A2(_0034_),
    .Z(_0052_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2544_ (.A1(_0049_),
    .A2(_0050_),
    .ZN(_0053_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2545_ (.A1(_0051_),
    .A2(_0052_),
    .B(_0053_),
    .ZN(_0055_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2546_ (.A1(_1567_),
    .A2(_1568_),
    .ZN(_0056_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2547_ (.A1(_0055_),
    .A2(_0056_),
    .Z(_0057_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2548_ (.A1(_0055_),
    .A2(_0056_),
    .ZN(_0058_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2549_ (.A1(_0038_),
    .A2(_0057_),
    .B(_0058_),
    .ZN(_0059_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2550_ (.A1(_1550_),
    .A2(_1572_),
    .Z(_0060_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2551_ (.A1(_0059_),
    .A2(_0060_),
    .Z(_0061_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2552_ (.A1(_0059_),
    .A2(_0060_),
    .Z(_0062_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2553_ (.A1(_0036_),
    .A2(_0061_),
    .B(_0062_),
    .ZN(_0063_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2554_ (.A1(_1549_),
    .A2(_1577_),
    .Z(_0064_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2555_ (.A1(_0063_),
    .A2(_0064_),
    .ZN(_0066_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2556_ (.A1(_0063_),
    .A2(_0064_),
    .ZN(_0067_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2557_ (.A1(_1265_),
    .A2(_0066_),
    .B(_0067_),
    .ZN(_0068_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2558_ (.A1(_1172_),
    .A2(_1579_),
    .A3(_1580_),
    .Z(_0069_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2559_ (.A1(_1583_),
    .A2(_1588_),
    .B1(_0068_),
    .B2(_0069_),
    .ZN(_0070_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2560_ (.A1(_0063_),
    .A2(_0064_),
    .Z(_0071_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2561_ (.A1(_1265_),
    .A2(_0071_),
    .Z(_0072_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2562_ (.A1(_1056_),
    .A2(_1379_),
    .ZN(_0073_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2563_ (.A1(_1379_),
    .A2(_1432_),
    .B(_0073_),
    .ZN(_0074_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2564_ (.A1(_1132_),
    .A2(_0074_),
    .Z(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2565_ (.A1(_1535_),
    .A2(_1541_),
    .B(_1596_),
    .ZN(_0077_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2566_ (.A1(_0073_),
    .A2(_0075_),
    .B(_0077_),
    .ZN(_0078_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2567_ (.A1(_1267_),
    .A2(_0078_),
    .ZN(_0079_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2568_ (.A1(_1267_),
    .A2(_0078_),
    .Z(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2569_ (.A1(_0073_),
    .A2(_0075_),
    .ZN(_0081_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2570_ (.A1(_0081_),
    .A2(_0077_),
    .ZN(_0082_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2571_ (.I0(_0865_),
    .I1(_0042_),
    .S(_1506_),
    .Z(_0083_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2572_ (.A1(_0900_),
    .A2(_0042_),
    .B1(_0083_),
    .B2(_1159_),
    .ZN(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2573_ (.A1(_1539_),
    .A2(_0044_),
    .Z(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2574_ (.A1(_0084_),
    .A2(_0085_),
    .Z(_0086_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2575_ (.A1(_1132_),
    .A2(_0074_),
    .Z(_0088_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2576_ (.A1(_0084_),
    .A2(_0085_),
    .ZN(_0089_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2577_ (.A1(_0086_),
    .A2(_0088_),
    .B(_0089_),
    .ZN(_0090_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2578_ (.A1(_0040_),
    .A2(_0041_),
    .ZN(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2579_ (.A1(_0045_),
    .A2(_0091_),
    .A3(_0047_),
    .Z(_0092_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2580_ (.A1(_0090_),
    .A2(_0092_),
    .Z(_0093_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2581_ (.A1(_0090_),
    .A2(_0092_),
    .ZN(_0094_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2582_ (.A1(_0082_),
    .A2(_0093_),
    .B(_0094_),
    .ZN(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _2583_ (.A1(_0049_),
    .A2(_0050_),
    .A3(_0052_),
    .ZN(_0096_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2584_ (.A1(_0095_),
    .A2(_0096_),
    .Z(_0097_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2585_ (.A1(_0095_),
    .A2(_0096_),
    .ZN(_0099_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2586_ (.A1(_0080_),
    .A2(_0097_),
    .B(_0099_),
    .ZN(_0100_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2587_ (.A1(_0038_),
    .A2(_0057_),
    .ZN(_0101_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2588_ (.A1(_0100_),
    .A2(_0101_),
    .Z(_0102_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _2589_ (.A1(_0036_),
    .A2(_0059_),
    .A3(_0060_),
    .ZN(_0103_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2590_ (.A1(_0100_),
    .A2(_0101_),
    .ZN(_0104_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _2591_ (.A1(_0079_),
    .A2(_0102_),
    .B(_0103_),
    .C(_0104_),
    .ZN(_0105_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2592_ (.A1(_0080_),
    .A2(_0097_),
    .ZN(_0106_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2593_ (.A1(_1159_),
    .A2(_0083_),
    .Z(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2594_ (.A1(_0913_),
    .A2(_1248_),
    .ZN(_0108_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2595_ (.I0(_0913_),
    .I1(_0108_),
    .S(_1506_),
    .Z(_0110_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2596_ (.A1(_0900_),
    .A2(_0108_),
    .B1(_0110_),
    .B2(_1385_),
    .ZN(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2597_ (.A1(_1159_),
    .A2(_0083_),
    .ZN(_0112_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2598_ (.A1(_1435_),
    .A2(_1289_),
    .ZN(_0113_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2599_ (.A1(_1432_),
    .A2(_0113_),
    .ZN(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2600_ (.A1(_1056_),
    .A2(_0113_),
    .B(_0114_),
    .ZN(_0115_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2601_ (.A1(_1534_),
    .A2(_0115_),
    .Z(_0116_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2602_ (.A1(_0107_),
    .A2(_0112_),
    .ZN(_0117_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2603_ (.A1(_0111_),
    .A2(_0117_),
    .Z(_0118_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2604_ (.A1(_0107_),
    .A2(_0111_),
    .A3(_0112_),
    .B1(_0116_),
    .B2(_0118_),
    .ZN(_0119_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2605_ (.A1(_0086_),
    .A2(_0088_),
    .Z(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2606_ (.A1(_0119_),
    .A2(_0121_),
    .ZN(_0122_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2607_ (.A1(_1056_),
    .A2(_0113_),
    .B1(_0115_),
    .B2(_1535_),
    .ZN(_0123_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2608_ (.A1(_0119_),
    .A2(_0121_),
    .Z(_0124_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2609_ (.A1(_0123_),
    .A2(_0124_),
    .ZN(_0125_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2610_ (.A1(_0082_),
    .A2(_0093_),
    .ZN(_0126_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2611_ (.A1(_0122_),
    .A2(_0125_),
    .B(_0126_),
    .ZN(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2612_ (.A1(_0080_),
    .A2(_0097_),
    .Z(_0128_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2613_ (.I(_0079_),
    .ZN(_0129_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2614_ (.A1(_0038_),
    .A2(_0057_),
    .Z(_0130_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2615_ (.A1(_0129_),
    .A2(_0100_),
    .A3(_0130_),
    .Z(_0132_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _2616_ (.A1(_0106_),
    .A2(_0127_),
    .A3(_0128_),
    .A4(_0132_),
    .ZN(_0133_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2617_ (.A1(_0100_),
    .A2(_0130_),
    .Z(_0134_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2618_ (.A1(_0100_),
    .A2(_0101_),
    .Z(_0135_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2619_ (.A1(_0129_),
    .A2(_0134_),
    .B(_0135_),
    .ZN(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2620_ (.A1(_0136_),
    .A2(_0103_),
    .ZN(_0137_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2621_ (.A1(_0105_),
    .A2(_0133_),
    .B(_0137_),
    .ZN(_0138_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2622_ (.A1(_0136_),
    .A2(_0103_),
    .ZN(_0139_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2623_ (.A1(_1403_),
    .A2(_1142_),
    .ZN(_0140_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2624_ (.A1(_0108_),
    .A2(_1556_),
    .ZN(_0141_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2625_ (.A1(_0913_),
    .A2(_0140_),
    .B1(_0141_),
    .B2(_1402_),
    .ZN(_0143_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2626_ (.I(_0143_),
    .ZN(_0144_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2627_ (.A1(_1385_),
    .A2(_0110_),
    .ZN(_0145_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2628_ (.A1(_0144_),
    .A2(_0145_),
    .ZN(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2629_ (.A1(_1078_),
    .A2(_1435_),
    .B(_1289_),
    .ZN(_0147_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2630_ (.A1(_1078_),
    .A2(_1489_),
    .B(_0147_),
    .ZN(_0148_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2631_ (.A1(_1379_),
    .A2(_0148_),
    .Z(_0149_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2632_ (.A1(_0143_),
    .A2(_0145_),
    .Z(_0150_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2633_ (.A1(_0149_),
    .A2(_0150_),
    .ZN(_0151_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2634_ (.A1(_0116_),
    .A2(_0118_),
    .Z(_0152_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2635_ (.A1(_0146_),
    .A2(_0151_),
    .B(_0152_),
    .ZN(_0154_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2636_ (.A1(_1079_),
    .A2(_0113_),
    .B1(_0147_),
    .B2(_1379_),
    .ZN(_0155_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _2637_ (.A1(_0146_),
    .A2(_0151_),
    .A3(_0152_),
    .Z(_0156_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2638_ (.A1(_0154_),
    .A2(_0156_),
    .Z(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2639_ (.A1(_0155_),
    .A2(_0157_),
    .ZN(_0158_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2640_ (.A1(_0154_),
    .A2(_0158_),
    .ZN(_0159_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2641_ (.A1(_0123_),
    .A2(_0124_),
    .Z(_0160_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2642_ (.A1(_0155_),
    .A2(_0157_),
    .ZN(_0161_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2643_ (.I(_1590_),
    .ZN(_0162_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2644_ (.A1(_0926_),
    .A2(_1506_),
    .ZN(_0163_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2645_ (.A1(_1506_),
    .A2(_0140_),
    .B(_0163_),
    .ZN(_0165_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2646_ (.A1(_0162_),
    .A2(_0165_),
    .B(_0163_),
    .ZN(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2647_ (.I0(_1556_),
    .I1(_0926_),
    .S(_0108_),
    .Z(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2648_ (.A1(_1402_),
    .A2(_0167_),
    .Z(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2649_ (.A1(_0166_),
    .A2(_0168_),
    .ZN(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2650_ (.A1(_1536_),
    .A2(_1590_),
    .ZN(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2651_ (.A1(_1079_),
    .A2(_1590_),
    .B(_0170_),
    .ZN(_0171_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2652_ (.A1(_1432_),
    .A2(_0171_),
    .Z(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2653_ (.A1(_0166_),
    .A2(_0168_),
    .Z(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2654_ (.A1(_0172_),
    .A2(_0173_),
    .Z(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2655_ (.A1(_0149_),
    .A2(_0150_),
    .Z(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2656_ (.A1(_0169_),
    .A2(_0174_),
    .B(_0176_),
    .ZN(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _2657_ (.A1(_0176_),
    .A2(_0169_),
    .A3(_0174_),
    .Z(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2658_ (.A1(_0178_),
    .A2(_0177_),
    .ZN(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2659_ (.A1(_1432_),
    .A2(_0171_),
    .ZN(_0180_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2660_ (.A1(_1078_),
    .A2(_0162_),
    .B(_0180_),
    .ZN(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2661_ (.A1(_1078_),
    .A2(_0108_),
    .B(_1556_),
    .C(_0162_),
    .ZN(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2662_ (.A1(_1078_),
    .A2(_1289_),
    .A3(_0108_),
    .ZN(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2663_ (.A1(_0182_),
    .A2(_0183_),
    .Z(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2664_ (.A1(_0162_),
    .A2(_0165_),
    .Z(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2665_ (.A1(_0113_),
    .A2(_0184_),
    .ZN(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2666_ (.A1(_0185_),
    .A2(_0187_),
    .ZN(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2667_ (.A1(_0113_),
    .A2(_0184_),
    .B(_0188_),
    .C(_0174_),
    .ZN(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2668_ (.A1(_0172_),
    .A2(_0173_),
    .B(_0189_),
    .ZN(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2669_ (.A1(_0161_),
    .A2(_0177_),
    .B1(_0179_),
    .B2(_0181_),
    .C(_0190_),
    .ZN(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2670_ (.A1(_0181_),
    .A2(_0179_),
    .Z(_0192_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2671_ (.A1(_0177_),
    .A2(_0192_),
    .B(_0161_),
    .ZN(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2672_ (.A1(_0159_),
    .A2(_0160_),
    .B(_0191_),
    .C(_0193_),
    .ZN(_0194_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2673_ (.A1(_0122_),
    .A2(_0125_),
    .ZN(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2674_ (.A1(_0126_),
    .A2(_0195_),
    .Z(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2675_ (.A1(_0159_),
    .A2(_0160_),
    .ZN(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _2676_ (.A1(_0194_),
    .A2(_0196_),
    .A3(_0198_),
    .Z(_0199_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2677_ (.A1(_0129_),
    .A2(_0134_),
    .ZN(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2678_ (.A1(_0106_),
    .A2(_0128_),
    .ZN(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2679_ (.A1(_0079_),
    .A2(_0102_),
    .B(_0201_),
    .ZN(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2680_ (.A1(_0200_),
    .A2(_0202_),
    .ZN(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2681_ (.A1(_0133_),
    .A2(_0139_),
    .B(_0199_),
    .C(_0203_),
    .ZN(_0204_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _2682_ (.A1(_1263_),
    .A2(_1525_),
    .A3(_1526_),
    .ZN(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _2683_ (.A1(_1264_),
    .A2(_1585_),
    .B(_1586_),
    .C(_0205_),
    .ZN(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _2684_ (.A1(_0068_),
    .A2(_0069_),
    .B1(_0138_),
    .B2(_0204_),
    .C(_0206_),
    .ZN(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2685_ (.A1(_1584_),
    .A2(_0070_),
    .B1(_0072_),
    .B2(_0207_),
    .ZN(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2686_ (.A1(_1483_),
    .A2(_1484_),
    .ZN(_0210_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2687_ (.A1(_1486_),
    .A2(_1529_),
    .ZN(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2688_ (.A1(_1431_),
    .A2(_0210_),
    .A3(_0211_),
    .ZN(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2689_ (.A1(_1327_),
    .A2(_1374_),
    .ZN(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2690_ (.A1(_1376_),
    .A2(_1429_),
    .Z(_0214_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2691_ (.A1(_1374_),
    .A2(_0214_),
    .ZN(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2692_ (.A1(_0213_),
    .A2(_0215_),
    .ZN(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2693_ (.A1(_0209_),
    .A2(_0212_),
    .B(_0216_),
    .ZN(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2694_ (.A1(_1351_),
    .A2(_1353_),
    .ZN(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2695_ (.A1(_1288_),
    .A2(_1173_),
    .ZN(_0220_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2696_ (.A1(_1340_),
    .A2(_1341_),
    .ZN(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2697_ (.A1(_1340_),
    .A2(_0220_),
    .B(_0221_),
    .ZN(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2698_ (.A1(_1339_),
    .A2(_1343_),
    .ZN(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2699_ (.A1(_0218_),
    .A2(_0222_),
    .Z(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2700_ (.I(_0224_),
    .ZN(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2701_ (.A1(_0223_),
    .A2(_0225_),
    .ZN(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2702_ (.A1(_0218_),
    .A2(_0222_),
    .B(_0226_),
    .ZN(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2703_ (.A1(_1354_),
    .A2(_1364_),
    .B(_1362_),
    .ZN(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2704_ (.A1(_0815_),
    .A2(_1314_),
    .B1(_1357_),
    .B2(_1358_),
    .ZN(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _2705_ (.A1(_1025_),
    .A2(_1151_),
    .B1(_1305_),
    .B2(_0996_),
    .ZN(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2706_ (.A1(_1265_),
    .A2(_0231_),
    .Z(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2707_ (.A1(_0229_),
    .A2(_0232_),
    .Z(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2708_ (.A1(_1359_),
    .A2(_1360_),
    .ZN(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2709_ (.A1(_0799_),
    .A2(_0809_),
    .ZN(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2710_ (.A1(_0235_),
    .A2(_1248_),
    .B1(_1304_),
    .B2(_1017_),
    .ZN(_0236_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_4 _2711_ (.A1(_0749_),
    .A2(_1317_),
    .B1(_1318_),
    .B2(_0848_),
    .C1(_1252_),
    .C2(_0794_),
    .ZN(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2712_ (.A1(_0236_),
    .A2(_0237_),
    .ZN(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2713_ (.A1(_0234_),
    .A2(_0238_),
    .Z(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2714_ (.A1(_0233_),
    .A2(_0239_),
    .Z(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2715_ (.A1(_0228_),
    .A2(_0240_),
    .ZN(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2716_ (.A1(_0223_),
    .A2(_0225_),
    .Z(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2717_ (.A1(_0228_),
    .A2(_0240_),
    .Z(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2718_ (.A1(_0243_),
    .A2(_0244_),
    .ZN(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2719_ (.A1(_0242_),
    .A2(_0245_),
    .ZN(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2720_ (.A1(_0229_),
    .A2(_0232_),
    .ZN(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2721_ (.A1(_0221_),
    .A2(_0247_),
    .ZN(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2722_ (.A1(_0234_),
    .A2(_0238_),
    .ZN(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2723_ (.A1(_0233_),
    .A2(_0239_),
    .B(_0249_),
    .ZN(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2724_ (.A1(_1120_),
    .A2(_0231_),
    .ZN(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2725_ (.A1(_0985_),
    .A2(_1305_),
    .ZN(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2726_ (.A1(_1172_),
    .A2(_0253_),
    .ZN(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2727_ (.A1(_0235_),
    .A2(_1357_),
    .ZN(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2728_ (.A1(_0254_),
    .A2(_0255_),
    .Z(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2729_ (.A1(_0251_),
    .A2(_0256_),
    .ZN(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2730_ (.A1(_0236_),
    .A2(_0237_),
    .ZN(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2731_ (.A1(_1007_),
    .A2(_1151_),
    .ZN(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2732_ (.A1(_1025_),
    .A2(_1164_),
    .B(_1143_),
    .ZN(_0260_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2733_ (.A1(_0259_),
    .A2(_0260_),
    .ZN(_0261_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _2734_ (.A1(_1157_),
    .A2(_1187_),
    .B1(_1189_),
    .B2(_1300_),
    .C1(_1212_),
    .C2(_1193_),
    .ZN(_0262_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2735_ (.A1(_0261_),
    .A2(_0262_),
    .ZN(_0264_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2736_ (.A1(_0258_),
    .A2(_0264_),
    .Z(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2737_ (.A1(_0257_),
    .A2(_0265_),
    .ZN(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2738_ (.A1(_0250_),
    .A2(_0266_),
    .ZN(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2739_ (.A1(_0248_),
    .A2(_0267_),
    .ZN(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2740_ (.A1(_0227_),
    .A2(_0246_),
    .A3(_0268_),
    .Z(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2741_ (.A1(_1338_),
    .A2(_1344_),
    .ZN(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2742_ (.A1(_1335_),
    .A2(_1346_),
    .B(_0270_),
    .ZN(_0271_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2743_ (.I(_0271_),
    .ZN(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2744_ (.A1(_1347_),
    .A2(_1366_),
    .Z(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2745_ (.A1(_1350_),
    .A2(_1365_),
    .B(_0273_),
    .ZN(_0275_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2746_ (.A1(_0243_),
    .A2(_0244_),
    .ZN(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2747_ (.A1(_0275_),
    .A2(_0276_),
    .Z(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2748_ (.A1(_0275_),
    .A2(_0276_),
    .Z(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2749_ (.A1(_0272_),
    .A2(_0277_),
    .B(_0278_),
    .ZN(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2750_ (.A1(_0269_),
    .A2(_0279_),
    .ZN(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2751_ (.I(_0268_),
    .ZN(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2752_ (.A1(_0246_),
    .A2(_0281_),
    .ZN(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2753_ (.A1(_0246_),
    .A2(_0281_),
    .ZN(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2754_ (.A1(_0227_),
    .A2(_0282_),
    .B(_0283_),
    .ZN(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2755_ (.A1(_0221_),
    .A2(_0247_),
    .Z(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2756_ (.A1(_0250_),
    .A2(_0266_),
    .ZN(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2757_ (.A1(_0248_),
    .A2(_0267_),
    .ZN(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2758_ (.A1(_0287_),
    .A2(_0288_),
    .ZN(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2759_ (.A1(_1120_),
    .A2(_0231_),
    .A3(_0256_),
    .ZN(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2760_ (.A1(_0254_),
    .A2(_0255_),
    .B(_0290_),
    .ZN(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2761_ (.A1(_0257_),
    .A2(_0265_),
    .ZN(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2762_ (.A1(_0258_),
    .A2(_0264_),
    .B(_0292_),
    .ZN(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2763_ (.A1(_0259_),
    .A2(_0260_),
    .ZN(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2764_ (.A1(_0962_),
    .A2(_1305_),
    .ZN(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2765_ (.A1(_1263_),
    .A2(_0295_),
    .ZN(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2766_ (.A1(_0294_),
    .A2(_0297_),
    .Z(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2767_ (.A1(_0261_),
    .A2(_0262_),
    .ZN(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2768_ (.A1(_0996_),
    .A2(_1151_),
    .ZN(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2769_ (.A1(_1007_),
    .A2(_1304_),
    .B(_1165_),
    .ZN(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2770_ (.A1(_0300_),
    .A2(_0301_),
    .Z(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_4 _2771_ (.A1(_0794_),
    .A2(_1317_),
    .B1(_1318_),
    .B2(_0770_),
    .C1(_1252_),
    .C2(_0318_),
    .ZN(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2772_ (.A1(_0302_),
    .A2(_0303_),
    .Z(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2773_ (.A1(_0299_),
    .A2(_0304_),
    .Z(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2774_ (.A1(_0298_),
    .A2(_0305_),
    .Z(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2775_ (.A1(_0293_),
    .A2(_0306_),
    .Z(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2776_ (.A1(_0291_),
    .A2(_0308_),
    .ZN(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2777_ (.A1(_0286_),
    .A2(_0289_),
    .A3(_0309_),
    .Z(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2778_ (.A1(_0284_),
    .A2(_0310_),
    .Z(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2779_ (.A1(_0280_),
    .A2(_0311_),
    .Z(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2780_ (.A1(_0284_),
    .A2(_0310_),
    .ZN(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2781_ (.A1(_0294_),
    .A2(_0297_),
    .ZN(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2782_ (.A1(_0299_),
    .A2(_0304_),
    .Z(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2783_ (.A1(_0298_),
    .A2(_0305_),
    .B(_0315_),
    .ZN(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2784_ (.A1(_0300_),
    .A2(_0301_),
    .Z(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2785_ (.A1(_0965_),
    .A2(_1305_),
    .B(_1290_),
    .ZN(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2786_ (.A1(_0302_),
    .A2(_0303_),
    .ZN(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2787_ (.A1(_0985_),
    .A2(_1151_),
    .ZN(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2788_ (.A1(_0996_),
    .A2(_1304_),
    .B(_1224_),
    .ZN(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2789_ (.A1(_0321_),
    .A2(_0322_),
    .Z(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_4 _2790_ (.A1(_0812_),
    .A2(_1317_),
    .B1(_1318_),
    .B2(_0794_),
    .C1(_0373_),
    .C2(_1252_),
    .ZN(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2791_ (.A1(_0323_),
    .A2(_0324_),
    .ZN(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2792_ (.A1(_0320_),
    .A2(_0325_),
    .ZN(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2793_ (.A1(_0317_),
    .A2(_0319_),
    .A3(_0326_),
    .Z(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _2794_ (.A1(_0314_),
    .A2(_0316_),
    .A3(_0327_),
    .ZN(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2795_ (.A1(_0293_),
    .A2(_0306_),
    .Z(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2796_ (.A1(_0291_),
    .A2(_0308_),
    .B(_0330_),
    .ZN(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2797_ (.A1(_0328_),
    .A2(_0331_),
    .ZN(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2798_ (.A1(_0289_),
    .A2(_0309_),
    .ZN(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2799_ (.A1(_0289_),
    .A2(_0309_),
    .ZN(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2800_ (.A1(_0286_),
    .A2(_0333_),
    .B(_0334_),
    .ZN(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2801_ (.A1(_0332_),
    .A2(_0335_),
    .ZN(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2802_ (.A1(_0313_),
    .A2(_0336_),
    .ZN(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2803_ (.A1(_0312_),
    .A2(_0337_),
    .ZN(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2804_ (.I(_0338_),
    .ZN(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2805_ (.A1(_1370_),
    .A2(_1373_),
    .ZN(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2806_ (.A1(_1332_),
    .A2(_1368_),
    .Z(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2807_ (.A1(_1329_),
    .A2(_1369_),
    .B(_0342_),
    .ZN(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2808_ (.A1(_0275_),
    .A2(_0276_),
    .A3(_0272_),
    .Z(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2809_ (.A1(_0343_),
    .A2(_0344_),
    .Z(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2810_ (.A1(_0341_),
    .A2(_0345_),
    .Z(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2811_ (.A1(_0343_),
    .A2(_0344_),
    .Z(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2812_ (.A1(_0269_),
    .A2(_0279_),
    .ZN(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2813_ (.A1(_0347_),
    .A2(_0348_),
    .Z(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2814_ (.A1(_0346_),
    .A2(_0349_),
    .ZN(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _2815_ (.A1(_1533_),
    .A2(_0217_),
    .B(_0339_),
    .C(_0350_),
    .ZN(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2816_ (.A1(_0341_),
    .A2(_0345_),
    .ZN(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2817_ (.A1(_0347_),
    .A2(_0353_),
    .B(_0348_),
    .ZN(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2818_ (.A1(_0338_),
    .A2(_0354_),
    .Z(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2819_ (.A1(_0269_),
    .A2(_0279_),
    .A3(_0311_),
    .ZN(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2820_ (.A1(_0313_),
    .A2(_0356_),
    .B(_0336_),
    .ZN(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2821_ (.A1(_0355_),
    .A2(_0357_),
    .Z(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2822_ (.A1(_0317_),
    .A2(_0319_),
    .ZN(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2823_ (.I(_0359_),
    .ZN(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2824_ (.A1(_0317_),
    .A2(_0319_),
    .ZN(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2825_ (.A1(_0360_),
    .A2(_0361_),
    .A3(_0326_),
    .B1(_0325_),
    .B2(_0320_),
    .ZN(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2826_ (.I(_0363_),
    .ZN(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2827_ (.A1(_0321_),
    .A2(_0322_),
    .ZN(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2828_ (.I(_0365_),
    .ZN(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2829_ (.A1(_0969_),
    .A2(_1305_),
    .B(_1340_),
    .ZN(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2830_ (.A1(_0366_),
    .A2(_0367_),
    .Z(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2831_ (.A1(_0323_),
    .A2(_0324_),
    .ZN(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_4 _2832_ (.A1(_0318_),
    .A2(_1317_),
    .B1(_1318_),
    .B2(_0812_),
    .C1(_1252_),
    .C2(_0472_),
    .ZN(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2833_ (.A1(_0962_),
    .A2(_1151_),
    .ZN(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2834_ (.A1(_0985_),
    .A2(_1304_),
    .B(_1241_),
    .ZN(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2835_ (.A1(_0371_),
    .A2(_0372_),
    .Z(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2836_ (.A1(_0370_),
    .A2(_0374_),
    .Z(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2837_ (.A1(_0369_),
    .A2(_0375_),
    .Z(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2838_ (.A1(_0368_),
    .A2(_0376_),
    .Z(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2839_ (.A1(_0364_),
    .A2(_0377_),
    .Z(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2840_ (.A1(_0359_),
    .A2(_0378_),
    .Z(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2841_ (.A1(_0316_),
    .A2(_0327_),
    .ZN(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2842_ (.A1(_0316_),
    .A2(_0327_),
    .ZN(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2843_ (.A1(_0314_),
    .A2(_0380_),
    .B(_0381_),
    .ZN(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2844_ (.A1(_0379_),
    .A2(_0382_),
    .Z(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2845_ (.A1(_0328_),
    .A2(_0331_),
    .ZN(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2846_ (.A1(_0332_),
    .A2(_0335_),
    .ZN(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2847_ (.A1(_0385_),
    .A2(_0386_),
    .ZN(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2848_ (.A1(_0383_),
    .A2(_0387_),
    .Z(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2849_ (.A1(_0366_),
    .A2(_0367_),
    .ZN(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2850_ (.I(_0368_),
    .ZN(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2851_ (.A1(_0323_),
    .A2(_0324_),
    .A3(_0375_),
    .ZN(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2852_ (.A1(_0390_),
    .A2(_0376_),
    .B(_0391_),
    .ZN(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2853_ (.A1(_0972_),
    .A2(_1305_),
    .ZN(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2854_ (.A1(_0965_),
    .A2(_1151_),
    .B1(_1304_),
    .B2(_0962_),
    .ZN(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2855_ (.A1(_0393_),
    .A2(_0394_),
    .ZN(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_4 _2856_ (.A1(_0373_),
    .A2(_1317_),
    .B1(_1318_),
    .B2(_0318_),
    .C1(_1378_),
    .C2(_1252_),
    .ZN(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2857_ (.A1(_0396_),
    .A2(_0397_),
    .Z(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2858_ (.A1(_0371_),
    .A2(_0372_),
    .Z(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2859_ (.A1(_0370_),
    .A2(_0374_),
    .B(_0399_),
    .ZN(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2860_ (.A1(_0398_),
    .A2(_0400_),
    .Z(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2861_ (.A1(_0392_),
    .A2(_0401_),
    .Z(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2862_ (.A1(_0389_),
    .A2(_0402_),
    .Z(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2863_ (.A1(_0364_),
    .A2(_0377_),
    .ZN(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2864_ (.A1(_0360_),
    .A2(_0378_),
    .B(_0404_),
    .ZN(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2865_ (.A1(_0403_),
    .A2(_0405_),
    .Z(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2866_ (.A1(_0379_),
    .A2(_0382_),
    .ZN(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2867_ (.A1(_0385_),
    .A2(_0383_),
    .Z(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2868_ (.A1(_0408_),
    .A2(_0409_),
    .ZN(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2869_ (.A1(_0407_),
    .A2(_0410_),
    .Z(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2870_ (.A1(_0388_),
    .A2(_0411_),
    .Z(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2871_ (.I(_0412_),
    .ZN(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2872_ (.A1(_0352_),
    .A2(_0358_),
    .B(_0413_),
    .ZN(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2873_ (.A1(_0386_),
    .A2(_0383_),
    .ZN(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2874_ (.A1(_0415_),
    .A2(_0411_),
    .Z(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2875_ (.A1(_0409_),
    .A2(_0407_),
    .ZN(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2876_ (.A1(_0416_),
    .A2(_0418_),
    .ZN(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2877_ (.I(_0419_),
    .ZN(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2878_ (.A1(_0403_),
    .A2(_0405_),
    .ZN(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2879_ (.A1(_0366_),
    .A2(_0367_),
    .A3(_0402_),
    .Z(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2880_ (.A1(_0392_),
    .A2(_0401_),
    .B(_0422_),
    .ZN(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2881_ (.A1(_0969_),
    .A2(_1151_),
    .ZN(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2882_ (.A1(_0965_),
    .A2(_1304_),
    .ZN(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _2883_ (.A1(_0472_),
    .A2(_1317_),
    .B1(_1318_),
    .B2(_0373_),
    .ZN(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2884_ (.A1(_0425_),
    .A2(_0426_),
    .Z(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2885_ (.A1(_0424_),
    .A2(_0427_),
    .Z(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2886_ (.I(_0397_),
    .ZN(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2887_ (.A1(_0396_),
    .A2(_0430_),
    .ZN(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2888_ (.A1(_0398_),
    .A2(_0400_),
    .ZN(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2889_ (.A1(_0431_),
    .A2(_0432_),
    .ZN(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2890_ (.A1(_0429_),
    .A2(_0433_),
    .Z(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2891_ (.A1(_0423_),
    .A2(_0434_),
    .Z(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2892_ (.A1(_0421_),
    .A2(_0435_),
    .ZN(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2893_ (.A1(_0408_),
    .A2(_0407_),
    .ZN(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2894_ (.A1(_0421_),
    .A2(_0435_),
    .ZN(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2895_ (.A1(_0437_),
    .A2(_0438_),
    .ZN(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2896_ (.A1(_0408_),
    .A2(_0407_),
    .A3(_0435_),
    .ZN(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2897_ (.A1(_0440_),
    .A2(_0441_),
    .Z(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2898_ (.A1(_0436_),
    .A2(_0442_),
    .ZN(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2899_ (.A1(_0414_),
    .A2(_0420_),
    .B(_0443_),
    .ZN(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2900_ (.I(_1533_),
    .ZN(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2901_ (.A1(_1172_),
    .A2(_1581_),
    .B(_1582_),
    .ZN(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2902_ (.A1(_0063_),
    .A2(_0064_),
    .Z(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2903_ (.A1(_1120_),
    .A2(_0071_),
    .B(_0447_),
    .ZN(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _2904_ (.A1(_1264_),
    .A2(_1579_),
    .A3(_1580_),
    .Z(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _2905_ (.A1(_0205_),
    .A2(_0446_),
    .B1(_0448_),
    .B2(_0449_),
    .ZN(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2906_ (.A1(_1120_),
    .A2(_0071_),
    .Z(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2907_ (.A1(_0105_),
    .A2(_0133_),
    .ZN(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2908_ (.A1(_0136_),
    .A2(_0103_),
    .B(_0453_),
    .ZN(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2909_ (.A1(_0136_),
    .A2(_0103_),
    .Z(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2910_ (.A1(_0194_),
    .A2(_0196_),
    .A3(_0198_),
    .ZN(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2911_ (.A1(_0200_),
    .A2(_0202_),
    .Z(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _2912_ (.A1(_0127_),
    .A2(_0455_),
    .B(_0456_),
    .C(_0457_),
    .ZN(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2913_ (.A1(_0448_),
    .A2(_0449_),
    .B1(_0454_),
    .B2(_0458_),
    .C(_1584_),
    .ZN(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2914_ (.A1(_0206_),
    .A2(_0451_),
    .B1(_0452_),
    .B2(_0459_),
    .ZN(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _2915_ (.A1(_1431_),
    .A2(_0210_),
    .A3(_0211_),
    .Z(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _2916_ (.A1(_0460_),
    .A2(_0462_),
    .B(_0215_),
    .C(_0213_),
    .ZN(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2917_ (.A1(_0312_),
    .A2(_0337_),
    .A3(_0350_),
    .ZN(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2918_ (.A1(_0445_),
    .A2(_0463_),
    .B(_0464_),
    .ZN(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2919_ (.A1(_0355_),
    .A2(_0357_),
    .ZN(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2920_ (.A1(_0465_),
    .A2(_0466_),
    .B(_0412_),
    .ZN(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2921_ (.A1(_0436_),
    .A2(_0442_),
    .Z(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2922_ (.A1(_0467_),
    .A2(_0419_),
    .A3(_0468_),
    .ZN(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2923_ (.A1(_0465_),
    .A2(_0466_),
    .B(_0388_),
    .ZN(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2924_ (.A1(_0415_),
    .A2(_0411_),
    .ZN(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2925_ (.A1(_0470_),
    .A2(_0471_),
    .B(_0414_),
    .C(_0416_),
    .ZN(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2926_ (.A1(\freeRunCntr[11] ),
    .A2(_0444_),
    .A3(_0469_),
    .B1(\freeRunCntr[10] ),
    .B2(_0473_),
    .ZN(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2927_ (.I(_0388_),
    .ZN(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2928_ (.A1(_0352_),
    .A2(_0358_),
    .A3(_0475_),
    .ZN(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2929_ (.A1(_0470_),
    .A2(_0476_),
    .Z(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2930_ (.A1(\freeRunCntr[10] ),
    .A2(_0473_),
    .B1(_0477_),
    .B2(_0560_),
    .ZN(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2931_ (.I(\freeRunCntr[6] ),
    .ZN(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2932_ (.A1(_0445_),
    .A2(_0463_),
    .ZN(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2933_ (.I(_0346_),
    .ZN(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2934_ (.A1(_0480_),
    .A2(_0481_),
    .B(_0353_),
    .ZN(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2935_ (.A1(_0349_),
    .A2(_0482_),
    .Z(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2936_ (.A1(_1533_),
    .A2(_0217_),
    .B(_0350_),
    .ZN(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2937_ (.A1(_0354_),
    .A2(_0485_),
    .ZN(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2938_ (.A1(_0312_),
    .A2(_0486_),
    .Z(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2939_ (.A1(_0479_),
    .A2(_0484_),
    .B1(_0487_),
    .B2(_0946_),
    .ZN(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2940_ (.A1(_1485_),
    .A2(_0460_),
    .A3(_0211_),
    .B(_1531_),
    .ZN(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2941_ (.A1(_1430_),
    .A2(_0489_),
    .B(_0214_),
    .ZN(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2942_ (.A1(_1375_),
    .A2(_0490_),
    .Z(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2943_ (.A1(_0460_),
    .A2(_0211_),
    .ZN(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2944_ (.A1(_0460_),
    .A2(_0211_),
    .Z(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _2945_ (.A1(\freeRunCntr[2] ),
    .A2(\freeRunCntr[1] ),
    .A3(_0492_),
    .A4(_0493_),
    .ZN(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2946_ (.A1(_1486_),
    .A2(_1529_),
    .ZN(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2947_ (.A1(_0460_),
    .A2(_0211_),
    .B(_0496_),
    .ZN(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2948_ (.A1(_0210_),
    .A2(_0497_),
    .ZN(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2949_ (.A1(\freeRunCntr[1] ),
    .A2(_0492_),
    .A3(_0493_),
    .B(\freeRunCntr[2] ),
    .ZN(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2950_ (.A1(_0495_),
    .A2(_0498_),
    .B(_0499_),
    .ZN(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2951_ (.A1(_1430_),
    .A2(_0489_),
    .ZN(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2952_ (.A1(\freeRunCntr[3] ),
    .A2(_0501_),
    .Z(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2953_ (.A1(\freeRunCntr[3] ),
    .A2(_0501_),
    .Z(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2954_ (.A1(\freeRunCntr[4] ),
    .A2(_0491_),
    .B1(_0500_),
    .B2(_0502_),
    .C(_0503_),
    .ZN(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2955_ (.A1(_0480_),
    .A2(_0346_),
    .Z(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2956_ (.A1(_0882_),
    .A2(_0506_),
    .B1(_0491_),
    .B2(\freeRunCntr[4] ),
    .ZN(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2957_ (.A1(_0882_),
    .A2(_0506_),
    .ZN(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _2958_ (.A1(_0479_),
    .A2(_0484_),
    .B1(_0504_),
    .B2(_0507_),
    .C(_0508_),
    .ZN(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2959_ (.I(_0312_),
    .ZN(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2960_ (.A1(_0354_),
    .A2(_0485_),
    .B(_0510_),
    .ZN(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2961_ (.A1(_0356_),
    .A2(_0337_),
    .A3(_0511_),
    .Z(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2962_ (.A1(_0356_),
    .A2(_0511_),
    .B(_0337_),
    .ZN(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2963_ (.A1(_0512_),
    .A2(_0513_),
    .Z(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2964_ (.A1(_0946_),
    .A2(_0487_),
    .ZN(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2965_ (.A1(_0488_),
    .A2(_0509_),
    .B1(_0514_),
    .B2(\freeRunCntr[8] ),
    .C(_0515_),
    .ZN(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2966_ (.I(\freeRunCntr[10] ),
    .ZN(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2967_ (.A1(_0352_),
    .A2(_0358_),
    .B(_0475_),
    .ZN(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2968_ (.A1(_0415_),
    .A2(_0411_),
    .Z(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2969_ (.I(_0416_),
    .ZN(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2970_ (.A1(_0519_),
    .A2(_0520_),
    .B(_0467_),
    .C(_0521_),
    .ZN(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2971_ (.A1(_0470_),
    .A2(_0476_),
    .B(_0560_),
    .ZN(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2972_ (.A1(_0518_),
    .A2(_0522_),
    .B(_0523_),
    .ZN(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2973_ (.A1(\freeRunCntr[8] ),
    .A2(_0512_),
    .A3(_0513_),
    .B1(_0477_),
    .B2(_0560_),
    .ZN(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _2974_ (.A1(_0474_),
    .A2(_0524_),
    .A3(_0525_),
    .Z(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2975_ (.A1(_0432_),
    .A2(_0429_),
    .Z(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2976_ (.A1(_0424_),
    .A2(_0427_),
    .ZN(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2977_ (.A1(_0431_),
    .A2(_0429_),
    .ZN(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2978_ (.A1(_0972_),
    .A2(_1151_),
    .ZN(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2979_ (.A1(_0425_),
    .A2(_0426_),
    .ZN(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2980_ (.A1(_0969_),
    .A2(_1304_),
    .ZN(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2981_ (.A1(_1378_),
    .A2(_1317_),
    .B1(_1318_),
    .B2(_0472_),
    .ZN(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2982_ (.A1(_0533_),
    .A2(_0534_),
    .Z(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2983_ (.A1(_0532_),
    .A2(_0535_),
    .Z(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2984_ (.A1(_0531_),
    .A2(_0536_),
    .Z(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2985_ (.A1(_0529_),
    .A2(_0530_),
    .B(_0537_),
    .ZN(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2986_ (.A1(_0529_),
    .A2(_0537_),
    .A3(_0530_),
    .Z(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2987_ (.A1(_0539_),
    .A2(_0540_),
    .ZN(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2988_ (.A1(_0528_),
    .A2(_0541_),
    .Z(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2989_ (.A1(_0423_),
    .A2(_0434_),
    .ZN(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2990_ (.A1(_0421_),
    .A2(_0435_),
    .B(_0543_),
    .ZN(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2991_ (.A1(_0542_),
    .A2(_0544_),
    .Z(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2992_ (.I(_0545_),
    .ZN(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2993_ (.A1(_0441_),
    .A2(_0546_),
    .Z(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2994_ (.A1(_0467_),
    .A2(_0419_),
    .B(_0468_),
    .ZN(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2995_ (.I0(_0546_),
    .I1(_0547_),
    .S(_0548_),
    .Z(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2996_ (.A1(_0414_),
    .A2(_0420_),
    .A3(_0443_),
    .ZN(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2997_ (.A1(_0548_),
    .A2(_0551_),
    .B(_0814_),
    .ZN(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2998_ (.A1(\freeRunCntr[12] ),
    .A2(_0550_),
    .B(_0552_),
    .ZN(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _2999_ (.A1(_0474_),
    .A2(_0478_),
    .B1(_0517_),
    .B2(_0526_),
    .C(_0553_),
    .ZN(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3000_ (.I(_0542_),
    .ZN(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3001_ (.A1(_0436_),
    .A2(_0555_),
    .B1(_0545_),
    .B2(_0441_),
    .ZN(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3002_ (.A1(_0468_),
    .A2(_0546_),
    .ZN(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3003_ (.A1(_0420_),
    .A2(_0557_),
    .ZN(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _3004_ (.A1(_0465_),
    .A2(_0466_),
    .B(_0412_),
    .C(_0557_),
    .ZN(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3005_ (.A1(_0425_),
    .A2(_0426_),
    .A3(_0535_),
    .ZN(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _3006_ (.A1(_0972_),
    .A2(_1151_),
    .A3(_0536_),
    .B(_0561_),
    .ZN(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3007_ (.A1(_0533_),
    .A2(_0534_),
    .ZN(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3008_ (.A1(_0417_),
    .A2(_1189_),
    .ZN(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3009_ (.A1(_0972_),
    .A2(_1304_),
    .ZN(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3010_ (.A1(_0563_),
    .A2(_0564_),
    .A3(_0565_),
    .Z(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3011_ (.A1(_0562_),
    .A2(_0566_),
    .Z(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3012_ (.A1(_0539_),
    .A2(_0567_),
    .ZN(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3013_ (.A1(_0528_),
    .A2(_0541_),
    .Z(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3014_ (.A1(_0543_),
    .A2(_0542_),
    .B(_0569_),
    .ZN(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3015_ (.A1(_0568_),
    .A2(_0570_),
    .Z(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _3016_ (.A1(_0556_),
    .A2(_0558_),
    .A3(_0559_),
    .B(_0572_),
    .ZN(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3017_ (.A1(_0568_),
    .A2(_0570_),
    .ZN(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _3018_ (.A1(_0972_),
    .A2(_1304_),
    .A3(_0564_),
    .B(_0563_),
    .ZN(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3019_ (.A1(_0562_),
    .A2(_0566_),
    .B(_0574_),
    .C(_0575_),
    .ZN(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3020_ (.A1(\freeRunCntr[14] ),
    .A2(_0573_),
    .A3(_0576_),
    .Z(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3021_ (.A1(\freeRunCntr[15] ),
    .A2(\freeRunCntr[16] ),
    .ZN(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3022_ (.A1(\freeRunCntr[12] ),
    .A2(_0550_),
    .B(_0578_),
    .ZN(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3023_ (.A1(_0556_),
    .A2(_0558_),
    .A3(_0559_),
    .ZN(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3024_ (.A1(_0580_),
    .A2(_0572_),
    .Z(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3025_ (.A1(\freeRunCntr[13] ),
    .A2(_0581_),
    .ZN(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3026_ (.A1(_0573_),
    .A2(_0576_),
    .Z(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3027_ (.A1(_0580_),
    .A2(_0572_),
    .ZN(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3028_ (.I(\freeRunCntr[13] ),
    .ZN(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3029_ (.A1(\freeRunCntr[14] ),
    .A2(_0584_),
    .B1(_0585_),
    .B2(_0586_),
    .ZN(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _3030_ (.A1(_0577_),
    .A2(_0579_),
    .A3(_0583_),
    .A4(_0587_),
    .ZN(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3031_ (.A1(\freeRunCntr[14] ),
    .A2(_0584_),
    .ZN(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3032_ (.A1(\freeRunCntr[13] ),
    .A2(_0581_),
    .B(_0577_),
    .ZN(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3033_ (.A1(_0589_),
    .A2(_0590_),
    .B(_0578_),
    .ZN(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3034_ (.A1(_0554_),
    .A2(_0588_),
    .B(_0591_),
    .ZN(net6));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3035_ (.I(net4),
    .ZN(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3036_ (.A1(net2),
    .A2(net1),
    .A3(net3),
    .ZN(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3037_ (.A1(_0593_),
    .A2(_0594_),
    .Z(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3038_ (.A1(\freeRunCntr[0] ),
    .A2(_0595_),
    .ZN(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _3039_ (.I(net1),
    .ZN(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _3040_ (.A1(net2),
    .A2(_0597_),
    .A3(net3),
    .A4(net4),
    .ZN(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3041_ (.A1(\freeRunCntr[1] ),
    .A2(_0598_),
    .ZN(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3042_ (.A1(_0596_),
    .A2(_0599_),
    .Z(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3043_ (.I(_0600_),
    .Z(_0011_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3044_ (.I(net4),
    .Z(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3045_ (.A1(net2),
    .A2(_0597_),
    .ZN(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3046_ (.A1(net3),
    .A2(_0601_),
    .A3(_0603_),
    .ZN(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3047_ (.A1(\freeRunCntr[2] ),
    .A2(_0604_),
    .Z(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3048_ (.A1(\freeRunCntr[1] ),
    .A2(_0598_),
    .ZN(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3049_ (.A1(_0596_),
    .A2(_0599_),
    .B(_0606_),
    .ZN(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3050_ (.A1(_0605_),
    .A2(_0607_),
    .Z(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3051_ (.I(_0608_),
    .Z(_0022_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3052_ (.A1(net2),
    .A2(net1),
    .ZN(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3053_ (.A1(net3),
    .A2(_0601_),
    .A3(_0609_),
    .ZN(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3054_ (.A1(\freeRunCntr[2] ),
    .A2(_0604_),
    .Z(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3055_ (.A1(_0605_),
    .A2(_0607_),
    .B(_0611_),
    .ZN(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3056_ (.A1(_0885_),
    .A2(_0610_),
    .A3(_0613_),
    .Z(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3057_ (.I(_0614_),
    .Z(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3058_ (.A1(net2),
    .A2(net1),
    .ZN(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3059_ (.A1(net3),
    .A2(_0615_),
    .ZN(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3060_ (.A1(_0601_),
    .A2(_0616_),
    .ZN(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3061_ (.A1(\freeRunCntr[4] ),
    .A2(_0617_),
    .Z(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3062_ (.A1(\freeRunCntr[3] ),
    .A2(_0610_),
    .ZN(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3063_ (.A1(\freeRunCntr[3] ),
    .A2(_0610_),
    .ZN(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3064_ (.A1(_0619_),
    .A2(_0613_),
    .B(_0620_),
    .ZN(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3065_ (.A1(_0618_),
    .A2(_0621_),
    .Z(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3066_ (.I(_0623_),
    .Z(_0027_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3067_ (.I(net3),
    .Z(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3068_ (.A1(net2),
    .A2(_0597_),
    .ZN(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3069_ (.A1(_0624_),
    .A2(_0593_),
    .A3(_0625_),
    .Z(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3070_ (.A1(_0883_),
    .A2(_0601_),
    .A3(_0616_),
    .ZN(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3071_ (.A1(_0618_),
    .A2(_0621_),
    .B(_0627_),
    .ZN(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _3072_ (.A1(_0882_),
    .A2(_0626_),
    .A3(_0628_),
    .ZN(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3073_ (.I(_0629_),
    .Z(_0028_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3074_ (.A1(net2),
    .A2(_0597_),
    .Z(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3075_ (.A1(_0624_),
    .A2(_0630_),
    .ZN(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3076_ (.A1(_0601_),
    .A2(_0632_),
    .ZN(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3077_ (.A1(\freeRunCntr[6] ),
    .A2(_0633_),
    .Z(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3078_ (.A1(_0882_),
    .A2(_0626_),
    .ZN(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3079_ (.A1(_0882_),
    .A2(_0626_),
    .ZN(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3080_ (.A1(_0635_),
    .A2(_0628_),
    .B(_0636_),
    .ZN(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3081_ (.A1(_0634_),
    .A2(_0637_),
    .Z(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3082_ (.I(_0638_),
    .Z(_0029_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3083_ (.A1(net2),
    .A2(net1),
    .A3(_0624_),
    .ZN(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3084_ (.A1(_0601_),
    .A2(_0639_),
    .ZN(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3085_ (.A1(_0479_),
    .A2(_0601_),
    .A3(_0632_),
    .ZN(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3086_ (.A1(_0634_),
    .A2(_0637_),
    .B(_0642_),
    .ZN(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3087_ (.A1(_0946_),
    .A2(_0640_),
    .A3(_0643_),
    .Z(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3088_ (.I(_0644_),
    .Z(_0030_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3089_ (.A1(_0601_),
    .A2(_0594_),
    .B(\freeRunCntr[8] ),
    .ZN(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3090_ (.A1(\freeRunCntr[8] ),
    .A2(_0601_),
    .A3(_0594_),
    .Z(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3091_ (.A1(_0645_),
    .A2(_0646_),
    .ZN(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3092_ (.A1(\freeRunCntr[7] ),
    .A2(_0640_),
    .ZN(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3093_ (.A1(\freeRunCntr[7] ),
    .A2(_0640_),
    .ZN(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3094_ (.A1(_0648_),
    .A2(_0643_),
    .B(_0649_),
    .ZN(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3095_ (.A1(_0647_),
    .A2(_0650_),
    .Z(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3096_ (.I(_0652_),
    .Z(_0031_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3097_ (.I(_0601_),
    .Z(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3098_ (.A1(net2),
    .A2(_0597_),
    .A3(_0624_),
    .ZN(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3099_ (.A1(_0653_),
    .A2(_0654_),
    .ZN(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3100_ (.A1(_0647_),
    .A2(_0650_),
    .B(_0646_),
    .ZN(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3101_ (.A1(_0560_),
    .A2(_0655_),
    .A3(_0656_),
    .Z(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3102_ (.I(_0657_),
    .Z(_0032_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3103_ (.A1(_0624_),
    .A2(_0603_),
    .ZN(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3104_ (.A1(_0653_),
    .A2(_0658_),
    .B(\freeRunCntr[10] ),
    .ZN(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _3105_ (.A1(_0518_),
    .A2(_0624_),
    .A3(_0593_),
    .A4(_0603_),
    .ZN(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3106_ (.A1(_0659_),
    .A2(_0661_),
    .ZN(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3107_ (.A1(_0653_),
    .A2(_0654_),
    .B(_0560_),
    .ZN(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3108_ (.A1(_0560_),
    .A2(_0653_),
    .A3(_0654_),
    .ZN(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3109_ (.A1(_0663_),
    .A2(_0656_),
    .B(_0664_),
    .ZN(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3110_ (.A1(_0662_),
    .A2(_0665_),
    .Z(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3111_ (.I(_0666_),
    .Z(_0001_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3112_ (.A1(_0624_),
    .A2(_0609_),
    .ZN(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3113_ (.A1(_0653_),
    .A2(_0667_),
    .ZN(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3114_ (.A1(_0662_),
    .A2(_0665_),
    .B(_0661_),
    .ZN(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3115_ (.A1(\freeRunCntr[11] ),
    .A2(_0668_),
    .A3(_0669_),
    .Z(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3116_ (.I(_0671_),
    .Z(_0002_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3117_ (.I(\freeRunCntr[12] ),
    .ZN(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3118_ (.A1(_0624_),
    .A2(_0653_),
    .A3(_0615_),
    .ZN(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3119_ (.A1(_0672_),
    .A2(_0673_),
    .Z(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3120_ (.A1(_0653_),
    .A2(_0667_),
    .B(\freeRunCntr[11] ),
    .ZN(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3121_ (.A1(\freeRunCntr[11] ),
    .A2(_0653_),
    .A3(_0667_),
    .ZN(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3122_ (.A1(_0675_),
    .A2(_0669_),
    .B(_0676_),
    .ZN(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3123_ (.A1(_0674_),
    .A2(_0677_),
    .Z(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3124_ (.I(_0678_),
    .Z(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3125_ (.A1(_0624_),
    .A2(_0653_),
    .A3(_0625_),
    .ZN(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3126_ (.I(_0680_),
    .ZN(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3127_ (.A1(_0672_),
    .A2(_0673_),
    .ZN(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3128_ (.A1(_0674_),
    .A2(_0677_),
    .B(_0682_),
    .ZN(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3129_ (.A1(_0586_),
    .A2(_0681_),
    .A3(_0683_),
    .Z(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3130_ (.I(_0684_),
    .Z(_0004_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3131_ (.I(\freeRunCntr[14] ),
    .ZN(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3132_ (.A1(_0624_),
    .A2(_0653_),
    .A3(_0630_),
    .ZN(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3133_ (.A1(_0685_),
    .A2(_0686_),
    .Z(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3134_ (.A1(\freeRunCntr[13] ),
    .A2(_0681_),
    .ZN(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3135_ (.A1(\freeRunCntr[13] ),
    .A2(_0681_),
    .ZN(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3136_ (.A1(_0688_),
    .A2(_0683_),
    .B(_0690_),
    .ZN(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3137_ (.A1(_0687_),
    .A2(_0691_),
    .Z(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3138_ (.I(_0692_),
    .Z(_0005_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3139_ (.A1(_0593_),
    .A2(_0639_),
    .Z(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3140_ (.A1(_0685_),
    .A2(_0686_),
    .ZN(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3141_ (.A1(_0687_),
    .A2(_0691_),
    .B(_0694_),
    .ZN(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3142_ (.A1(\freeRunCntr[15] ),
    .A2(_0693_),
    .A3(_0695_),
    .Z(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3143_ (.I(_0696_),
    .Z(_0006_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3144_ (.I(_0693_),
    .ZN(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3145_ (.A1(\freeRunCntr[15] ),
    .A2(_0697_),
    .ZN(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3146_ (.A1(\freeRunCntr[15] ),
    .A2(_0697_),
    .ZN(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3147_ (.A1(_0699_),
    .A2(_0695_),
    .B(_0700_),
    .ZN(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3148_ (.A1(\freeRunCntr[16] ),
    .A2(_0701_),
    .Z(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3149_ (.I(_0702_),
    .Z(_0007_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3150_ (.A1(\freeRunCntr[16] ),
    .A2(_0701_),
    .Z(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3151_ (.A1(\freeRunCntr[17] ),
    .A2(_0703_),
    .Z(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3152_ (.I(_0704_),
    .Z(_0008_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3153_ (.A1(\freeRunCntr[17] ),
    .A2(_0703_),
    .ZN(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3154_ (.A1(_1433_),
    .A2(_0705_),
    .ZN(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3155_ (.I(_0706_),
    .Z(_0009_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3156_ (.I(_1466_),
    .ZN(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3157_ (.A1(_1433_),
    .A2(\freeRunCntr[17] ),
    .A3(_0703_),
    .ZN(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3158_ (.A1(_0708_),
    .A2(_0709_),
    .Z(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3159_ (.I(_0710_),
    .Z(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3160_ (.A1(_0708_),
    .A2(_0709_),
    .ZN(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3161_ (.A1(_1411_),
    .A2(_0711_),
    .Z(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3162_ (.I(_0712_),
    .Z(_0012_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3163_ (.A1(_1411_),
    .A2(_0711_),
    .ZN(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3164_ (.A1(\csTable.address[3] ),
    .A2(_0713_),
    .ZN(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3165_ (.I(_0714_),
    .Z(_0013_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3166_ (.A1(\csTable.address[3] ),
    .A2(_1411_),
    .A3(_0711_),
    .ZN(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3167_ (.A1(\csTable.address[4] ),
    .A2(_0716_),
    .ZN(_0717_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3168_ (.I(_0717_),
    .Z(_0014_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3169_ (.A1(\csTable.address[3] ),
    .A2(_1411_),
    .A3(\csTable.address[4] ),
    .A4(_0711_),
    .Z(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3170_ (.A1(\csTable.address[5] ),
    .A2(_0718_),
    .Z(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3171_ (.I(_0719_),
    .Z(_0015_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3172_ (.A1(\csTable.address[5] ),
    .A2(_0718_),
    .ZN(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3173_ (.A1(_1345_),
    .A2(_0720_),
    .ZN(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3174_ (.I(_0721_),
    .Z(_0016_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3175_ (.A1(_0955_),
    .A2(_0720_),
    .ZN(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3176_ (.A1(_0417_),
    .A2(_0720_),
    .B(_0723_),
    .ZN(_0017_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3177_ (.A1(_0955_),
    .A2(_1345_),
    .ZN(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3178_ (.A1(_0724_),
    .A2(_0720_),
    .ZN(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3179_ (.A1(\freeRunCntr[26] ),
    .A2(_0725_),
    .Z(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3180_ (.I(_0726_),
    .Z(_0018_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3181_ (.I(\freeRunCntr[26] ),
    .ZN(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3182_ (.A1(_0727_),
    .A2(_0724_),
    .A3(_0720_),
    .ZN(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3183_ (.A1(\freeRunCntr[27] ),
    .A2(_0728_),
    .Z(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3184_ (.I(_0729_),
    .Z(_0019_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3185_ (.A1(\freeRunCntr[27] ),
    .A2(_0728_),
    .ZN(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3186_ (.A1(\freeRunCntr[28] ),
    .A2(_0731_),
    .ZN(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3187_ (.I(_0732_),
    .Z(_0020_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _3188_ (.A1(\freeRunCntr[27] ),
    .A2(\freeRunCntr[28] ),
    .A3(_0728_),
    .ZN(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3189_ (.A1(_1140_),
    .A2(_0733_),
    .Z(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3190_ (.I(_0734_),
    .Z(_0021_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3191_ (.A1(_1140_),
    .A2(_0733_),
    .ZN(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3192_ (.A1(_1117_),
    .A2(_0735_),
    .Z(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3193_ (.I(_0736_),
    .Z(_0023_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3194_ (.A1(_1117_),
    .A2(_0735_),
    .ZN(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3195_ (.A1(_1116_),
    .A2(_0737_),
    .Z(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3196_ (.I(_0739_),
    .Z(_0024_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3197_ (.A1(_1124_),
    .A2(_0733_),
    .B(_1118_),
    .ZN(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3198_ (.A1(_1144_),
    .A2(_0737_),
    .B(_0740_),
    .ZN(_0025_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3199_ (.A1(\freeRunCntr[0] ),
    .A2(_0595_),
    .Z(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3200_ (.I(_0741_),
    .Z(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3201_ (.D(_0000_),
    .RN(net9),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\freeRunCntr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3202_ (.D(_0011_),
    .RN(net9),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\freeRunCntr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 _3203_ (.D(_0022_),
    .RN(net9),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\freeRunCntr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3204_ (.D(_0026_),
    .RN(net9),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\freeRunCntr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3205_ (.D(_0027_),
    .RN(net10),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\freeRunCntr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3206_ (.D(_0028_),
    .RN(net10),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\freeRunCntr[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3207_ (.D(_0029_),
    .RN(net10),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\freeRunCntr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3208_ (.D(_0030_),
    .RN(net10),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\freeRunCntr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3209_ (.D(_0031_),
    .RN(net9),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\freeRunCntr[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3210_ (.D(_0032_),
    .RN(net12),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\freeRunCntr[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 _3211_ (.D(_0001_),
    .RN(net12),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\freeRunCntr[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 _3212_ (.D(_0002_),
    .RN(net12),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\freeRunCntr[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3213_ (.D(_0003_),
    .RN(net12),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\freeRunCntr[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 _3214_ (.D(_0004_),
    .RN(net10),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\freeRunCntr[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3215_ (.D(_0005_),
    .RN(net10),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\freeRunCntr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3216_ (.D(_0006_),
    .RN(net10),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\freeRunCntr[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3217_ (.D(_0007_),
    .RN(net9),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\freeRunCntr[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3218_ (.D(_0008_),
    .RN(net11),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\freeRunCntr[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3219_ (.D(_0009_),
    .RN(net11),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\csTable.address[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3220_ (.D(_0010_),
    .RN(net9),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\csTable.address[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3221_ (.D(_0012_),
    .RN(net9),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\csTable.address[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3222_ (.D(_0013_),
    .RN(net9),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\csTable.address[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3223_ (.D(_0014_),
    .RN(net9),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\csTable.address[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3224_ (.D(_0015_),
    .RN(net11),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\csTable.address[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3225_ (.D(_0016_),
    .RN(net11),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\csTable.address[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3226_ (.D(_0017_),
    .RN(net10),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\csTable.address[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3227_ (.D(_0018_),
    .RN(net11),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\freeRunCntr[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3228_ (.D(_0019_),
    .RN(net11),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\freeRunCntr[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3229_ (.D(_0020_),
    .RN(net11),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\freeRunCntr[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 _3230_ (.D(_0021_),
    .RN(net10),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\sigRom.address[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3231_ (.D(_0023_),
    .RN(net10),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\sigRom.address[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3232_ (.D(_0024_),
    .RN(net11),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\sigRom.address[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3233_ (.D(_0025_),
    .RN(net11),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\sigRom.address[3] ));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_670 ();
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1 (.I(divSel[0]),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input2 (.I(divSel[1]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input3 (.I(divSel[2]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input4 (.I(divSel[3]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input5 (.I(rst),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output6 (.I(net6),
    .Z(qcomplex));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output7 (.I(net7),
    .Z(qcos));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output8 (.I(net8),
    .Z(qsin));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 fanout9 (.I(net12),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 fanout10 (.I(net11),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 fanout11 (.I(net12),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout12 (.I(net5),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_clk (.I(clk),
    .Z(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_2_0__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_2_1__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_2_2__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_2_3__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3202__D (.I(_0011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3203__D (.I(_0022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3204__D (.I(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3205__D (.I(_0027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3206__D (.I(_0028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3207__D (.I(_0029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2572__A2 (.I(_0042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2571__I1 (.I(_0042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2536__A2 (.I(_0042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2535__S (.I(_0042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2583__A1 (.I(_0049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2544__A1 (.I(_0049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2542__A1 (.I(_0049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2583__A2 (.I(_0050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2544__A2 (.I(_0050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2542__A2 (.I(_0050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1999__I0 (.I(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1930__A2 (.I(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1884__B (.I(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1826__B (.I(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1799__I (.I(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1795__I1 (.I(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1788__A2 (.I(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1776__A1 (.I(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1640__A2 (.I(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1627__I (.I(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1933__A1 (.I(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1856__A2 (.I(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1804__A1 (.I(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1774__A2 (.I(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1771__A1 (.I(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1747__A1 (.I(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1739__A2 (.I(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1703__A2 (.I(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1645__A2 (.I(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1628__B (.I(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2597__A2 (.I(_0083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2593__A2 (.I(_0083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2572__B1 (.I(_0083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2576__A1 (.I(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2574__A1 (.I(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2576__A2 (.I(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2574__A2 (.I(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2014__B (.I(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1988__B (.I(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1794__B (.I(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1789__C (.I(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1787__C (.I(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1695__A2 (.I(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1630__I (.I(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2581__A2 (.I(_0092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2580__A2 (.I(_0092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2010__B (.I(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1991__B2 (.I(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1962__C (.I(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1932__B (.I(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1793__C (.I(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1758__C (.I(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1688__B (.I(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1647__I (.I(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1642__I (.I(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1631__B (.I(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2604__A2 (.I(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2603__A1 (.I(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2608__A1 (.I(_0119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2606__A1 (.I(_0119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2014__A2 (.I(_0120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1795__I0 (.I(_0120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1792__A1 (.I(_0120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1788__A1 (.I(_0120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1756__B (.I(_0120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1746__A2 (.I(_0120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1686__I (.I(_0120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1680__B (.I(_0120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1640__B (.I(_0120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1633__I (.I(_0120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2912__A1 (.I(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2616__A2 (.I(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2043__A2 (.I(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1981__A1 (.I(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1977__A1 (.I(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1942__A1 (.I(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1927__A1 (.I(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1840__B (.I(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1701__C (.I(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1673__I (.I(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1652__A1 (.I(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1641__A1 (.I(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1937__A2 (.I(_0142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1884__A2 (.I(_0142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1826__A2 (.I(_0142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1794__A2 (.I(_0142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1792__A2 (.I(_0142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1789__A2 (.I(_0142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1776__A2 (.I(_0142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1725__A1 (.I(_0142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1638__I (.I(_0142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1636__A2 (.I(_0142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2632__A1 (.I(_0143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2626__I (.I(_0143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2632__A2 (.I(_0145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2628__A2 (.I(_0145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2014__A3 (.I(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1937__B (.I(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1802__A1 (.I(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1794__A1 (.I(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1789__A1 (.I(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1757__A1 (.I(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1752__A1 (.I(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1709__A2 (.I(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1639__A2 (.I(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1636__B (.I(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2642__A1 (.I(_0155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2639__A1 (.I(_0155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1910__A2 (.I(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1783__B1 (.I(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1652__A2 (.I(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1641__A2 (.I(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1887__I0 (.I(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1852__A1 (.I(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1844__A1 (.I(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1782__A1 (.I(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1739__A1 (.I(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1709__A1 (.I(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1703__A1 (.I(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1687__A1 (.I(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1675__I0 (.I(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1639__A1 (.I(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1992__A1 (.I(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1804__A2 (.I(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1782__A2 (.I(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1777__I (.I(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1752__A2 (.I(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1703__A3 (.I(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1690__A3 (.I(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1687__A2 (.I(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1675__S (.I(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1639__A3 (.I(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2681__B (.I(_0199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1837__C (.I(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1811__A1 (.I(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1734__B (.I(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1653__A2 (.I(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1641__B2 (.I(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2693__A1 (.I(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2947__A2 (.I(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2944__A2 (.I(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2943__A2 (.I(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2940__A3 (.I(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2915__A3 (.I(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2688__A3 (.I(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2936__A2 (.I(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2815__A2 (.I(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2720__A1 (.I(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2707__A1 (.I(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2045__A1 (.I(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2044__C (.I(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1979__C (.I(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1888__B (.I(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1883__C (.I(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1759__A1 (.I(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1736__A1 (.I(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1715__B (.I(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1702__C (.I(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1643__B2 (.I(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2727__A1 (.I(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2710__A1 (.I(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2013__A1 (.I(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2010__A1 (.I(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2008__B2 (.I(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2003__A1 (.I(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1960__A1 (.I(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1844__A2 (.I(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1755__B (.I(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1714__I (.I(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1688__A1 (.I(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1646__A1 (.I(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2763__A2 (.I(_0260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2733__A2 (.I(_0260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2767__A2 (.I(_0262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2735__A2 (.I(_0262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2023__A1 (.I(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1654__A2 (.I(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1648__A2 (.I(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2002__B (.I(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1981__C (.I(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1973__C (.I(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1966__A2 (.I(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1934__A1 (.I(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1839__A2 (.I(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1748__B (.I(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1681__I (.I(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1653__A1 (.I(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1648__A3 (.I(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2796__A1 (.I(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2776__A1 (.I(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2091__A2 (.I(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1650__A2 (.I(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2856__B2 (.I(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2832__A1 (.I(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2771__C2 (.I(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2201__A1 (.I(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2163__A1 (.I(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1670__A2 (.I(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1656__A2 (.I(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2011__C (.I(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1965__C (.I(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1960__B (.I(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1867__B (.I(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1846__A2 (.I(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1745__C (.I(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1729__I (.I(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1726__B (.I(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1676__I (.I(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1652__B (.I(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1914__A1 (.I(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1663__A2 (.I(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1654__B1 (.I(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2967__A1 (.I(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2928__A1 (.I(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2872__A1 (.I(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2883__B2 (.I(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2856__A1 (.I(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2790__C1 (.I(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2267__I0 (.I(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2262__A1 (.I(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2117__A1 (.I(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1665__A2 (.I(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1656__B1 (.I(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2376__A1 (.I(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2127__A1 (.I(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2039__A1 (.I(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2017__B (.I(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2016__A1 (.I(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2007__A1 (.I(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1976__A1 (.I(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1958__A1 (.I(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1920__A1 (.I(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1658__A1 (.I(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2886__I (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2857__A2 (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2888__A2 (.I(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2860__A2 (.I(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2193__A1 (.I(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1895__A1 (.I(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1798__A1 (.I(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1719__A1 (.I(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1659__I (.I(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2896__A2 (.I(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2893__A2 (.I(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2875__A2 (.I(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2869__A1 (.I(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2896__A1 (.I(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2893__A1 (.I(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2868__A1 (.I(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2996__A1 (.I(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2925__B (.I(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2899__A1 (.I(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3176__A1 (.I(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3008__A1 (.I(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2091__A1 (.I(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1876__A1 (.I(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1849__B (.I(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1848__A1 (.I(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1814__B (.I(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1813__A1 (.I(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1718__B (.I(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1664__A1 (.I(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3005__A2 (.I(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2979__A2 (.I(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2884__A2 (.I(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2012__C (.I(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1994__A1 (.I(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1991__C (.I(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1846__A1 (.I(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1839__A1 (.I(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1796__B (.I(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1661__I (.I(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2047__A1 (.I(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2046__A1 (.I(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1979__B (.I(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1974__C (.I(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1963__A1 (.I(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1886__B (.I(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1821__B (.I(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1759__C (.I(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1732__B (.I(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1662__I (.I(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1975__A1 (.I(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1946__A1 (.I(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1922__A1 (.I(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1915__A1 (.I(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1912__A1 (.I(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1860__C (.I(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1838__B (.I(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1803__A1 (.I(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1696__A1 (.I(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1663__A1 (.I(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2912__B (.I(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2913__B2 (.I(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2947__A1 (.I(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2944__A1 (.I(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2943__A1 (.I(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2940__A2 (.I(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2916__A1 (.I(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2932__A2 (.I(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2918__A2 (.I(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3004__A1 (.I(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2923__A1 (.I(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2920__A1 (.I(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2981__B2 (.I(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2883__A1 (.I(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2832__C2 (.I(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2306__I1 (.I(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2266__A1 (.I(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2176__A1 (.I(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1666__B1 (.I(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1665__B1 (.I(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3085__A1 (.I(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2958__A1 (.I(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2939__A1 (.I(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2958__A2 (.I(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2939__A2 (.I(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2965__A2 (.I(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2999__B1 (.I(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3105__A1 (.I(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2972__A1 (.I(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3007__A2 (.I(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2982__A2 (.I(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3004__C (.I(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3003__A2 (.I(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3023__A2 (.I(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3016__A2 (.I(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3023__A3 (.I(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3016__A3 (.I(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3108__A1 (.I(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3107__B (.I(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3101__A1 (.I(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2973__B2 (.I(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2971__B (.I(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2930__B2 (.I(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2059__A1 (.I(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2058__B2 (.I(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1900__A1 (.I(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1721__A1 (.I(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3018__A3 (.I(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3010__A2 (.I(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2034__A1 (.I(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2024__A1 (.I(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1868__A1 (.I(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1858__B (.I(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1842__A1 (.I(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1810__B (.I(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1708__C (.I(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1702__A1 (.I(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1694__A1 (.I(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1677__A1 (.I(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2044__A1 (.I(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1959__A1 (.I(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1887__I1 (.I(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1852__A2 (.I(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1840__A2 (.I(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1822__A2 (.I(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1755__A1 (.I(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1692__A1 (.I(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1690__A2 (.I(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1675__I1 (.I(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3129__A1 (.I(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3029__B2 (.I(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3034__A2 (.I(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3034__B (.I(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2045__A2 (.I(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1836__A1 (.I(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1677__A2 (.I(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3139__A1 (.I(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3105__A3 (.I(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3069__A2 (.I(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3037__A1 (.I(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3049__A1 (.I(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3042__A1 (.I(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3098__A2 (.I(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3074__A2 (.I(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3068__A2 (.I(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3045__A2 (.I(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3040__A2 (.I(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3097__I (.I(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3090__A2 (.I(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3089__A1 (.I(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3085__A2 (.I(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3084__A1 (.I(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3076__A1 (.I(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3070__A2 (.I(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3060__A1 (.I(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3053__A2 (.I(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3046__A2 (.I(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2042__B (.I(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2001__B2 (.I(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1950__B (.I(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1941__A1 (.I(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1940__C (.I(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1866__C (.I(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1820__C (.I(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1781__C (.I(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1705__B (.I(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1677__B (.I(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2011__A2 (.I(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1982__B1 (.I(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1682__A1 (.I(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2031__B1 (.I(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1980__A1 (.I(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1856__A3 (.I(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1842__A3 (.I(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1789__B1 (.I(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1775__B1 (.I(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1757__A2 (.I(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1735__A2 (.I(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1710__A1 (.I(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1680__A2 (.I(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3139__A2 (.I(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3084__A2 (.I(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1987__B1 (.I(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1970__A1 (.I(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1965__B1 (.I(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1682__A2 (.I(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3100__A2 (.I(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3095__A2 (.I(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2033__A1 (.I(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2025__B (.I(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1874__A1 (.I(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1873__A1 (.I(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1860__A1 (.I(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1859__A1 (.I(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1853__C (.I(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1816__B (.I(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1710__B (.I(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1682__B (.I(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3132__A2 (.I(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3125__A2 (.I(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3121__A2 (.I(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3120__A1 (.I(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3118__A2 (.I(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3113__A1 (.I(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3108__A2 (.I(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3107__A1 (.I(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3104__A1 (.I(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3099__A1 (.I(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1684__A2 (.I(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2038__A1 (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2027__A1 (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2026__B (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1957__A1 (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1919__A1 (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1875__A1 (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1855__B (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1810__A1 (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1717__C (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1684__B (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1698__A1 (.I(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1697__A2 (.I(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2002__A2 (.I(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1992__B2 (.I(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1980__A2 (.I(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1972__A1 (.I(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1701__B (.I(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1689__A1 (.I(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1980__B (.I(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1938__B (.I(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1856__A1 (.I(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1804__B (.I(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1787__A1 (.I(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1782__B (.I(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1733__I (.I(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1709__B (.I(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1693__A2 (.I(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1687__B (.I(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3150__A2 (.I(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3148__A2 (.I(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2004__A2 (.I(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1859__A2 (.I(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1827__A2 (.I(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1716__A2 (.I(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1689__A2 (.I(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3169__A4 (.I(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3166__A3 (.I(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3163__A2 (.I(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3161__A2 (.I(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1982__C (.I(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1970__A2 (.I(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1827__B (.I(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1689__B (.I(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1872__A1 (.I(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1770__A1 (.I(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1734__A2 (.I(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1708__A1 (.I(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1694__A2 (.I(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3197__A2 (.I(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3191__A2 (.I(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3189__A2 (.I(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2035__B2 (.I(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2013__A2 (.I(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1872__A2 (.I(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1841__A1 (.I(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1770__A2 (.I(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1734__A3 (.I(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1708__A2 (.I(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1694__A3 (.I(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1858__A2 (.I(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1694__B1 (.I(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1950__A2 (.I(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1866__B2 (.I(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1780__A2 (.I(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1694__B2 (.I(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2038__B2 (.I(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1993__A1 (.I(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1945__A1 (.I(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1929__A1 (.I(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1911__A1 (.I(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1696__B2 (.I(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1698__A2 (.I(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1697__A3 (.I(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2711__A1 (.I(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2472__A1 (.I(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2378__I0 (.I(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2332__I1 (.I(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2271__C1 (.I(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2201__A2 (.I(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1900__A2 (.I(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1721__A2 (.I(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2006__A1 (.I(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1954__C (.I(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1890__C (.I(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1874__B (.I(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1828__C (.I(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1809__A1 (.I(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1806__C (.I(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1785__A1 (.I(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1784__A1 (.I(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1706__A1 (.I(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1753__A3 (.I(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1705__A1 (.I(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2045__B1 (.I(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1990__A2 (.I(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1943__A2 (.I(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1932__A2 (.I(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1885__A2 (.I(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1853__B2 (.I(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1837__A2 (.I(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1705__A2 (.I(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2037__A2 (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2024__A3 (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1938__A2 (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1889__B1 (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1872__B (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1845__B1 (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1806__A2 (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1770__B (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1708__B (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1999__I1 (.I(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1959__B (.I(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1792__A3 (.I(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1751__A2 (.I(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1745__B1 (.I(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1730__I1 (.I(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1712__A2 (.I(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2031__A2 (.I(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1871__C (.I(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1716__A1 (.I(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2043__A1 (.I(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2002__A1 (.I(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1853__A1 (.I(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1819__A1 (.I(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1818__A1 (.I(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1805__A1 (.I(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1800__A1 (.I(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1778__A1 (.I(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1726__A1 (.I(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1715__A1 (.I(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1973__A1 (.I(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1969__A1 (.I(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1961__A1 (.I(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1951__A1 (.I(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1885__B2 (.I(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1883__A1 (.I(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1801__B (.I(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1740__A1 (.I(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1727__A1 (.I(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1715__A2 (.I(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2771__B2 (.I(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2428__A1 (.I(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2333__A1 (.I(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2308__C1 (.I(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2114__A1 (.I(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1900__B1 (.I(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1722__A2 (.I(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1721__B1 (.I(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2003__A3 (.I(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1964__A1 (.I(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1933__A2 (.I(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1727__A2 (.I(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1983__A1 (.I(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1939__A2 (.I(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1870__A2 (.I(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1776__B (.I(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1725__A2 (.I(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1964__A2 (.I(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1883__A2 (.I(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1874__A3 (.I(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1857__B (.I(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1837__A1 (.I(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1801__A1 (.I(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1727__A3 (.I(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2036__A1 (.I(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2032__A1 (.I(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2031__A1 (.I(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2025__A1 (.I(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1954__A1 (.I(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1825__A1 (.I(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1816__A1 (.I(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1775__B2 (.I(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1773__A1 (.I(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1731__A1 (.I(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2004__B (.I(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1972__B (.I(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1889__C (.I(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1885__C (.I(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1807__I (.I(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1783__C (.I(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1775__C (.I(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1772__B (.I(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1738__A1 (.I(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1731__A2 (.I(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1977__A2 (.I(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1787__A2 (.I(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1731__A3 (.I(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1743__A2 (.I(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1742__A1 (.I(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2041__A1 (.I(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1965__A1 (.I(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1940__B2 (.I(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1910__A1 (.I(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1907__A1 (.I(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1888__A1 (.I(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1819__B (.I(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1783__A1 (.I(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1779__A1 (.I(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1734__A1 (.I(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2036__A2 (.I(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1990__A1 (.I(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1989__B (.I(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1962__A1 (.I(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1940__A1 (.I(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1931__A1 (.I(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1820__B1 (.I(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1738__A2 (.I(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2003__A4 (.I(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1866__A2 (.I(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1740__A2 (.I(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1743__A3 (.I(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1742__A2 (.I(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2790__B2 (.I(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2771__A1 (.I(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2711__C2 (.I(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2152__A1 (.I(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1763__A2 (.I(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2021__A1 (.I(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2011__A1 (.I(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1953__A1 (.I(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1748__A1 (.I(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2021__A2 (.I(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2020__A1 (.I(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1825__A2 (.I(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1748__A2 (.I(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2709__A1 (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1761__A1 (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1760__A2 (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2025__A2 (.I(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1966__A3 (.I(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1962__B2 (.I(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1943__A1 (.I(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1932__A1 (.I(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1787__B1 (.I(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1753__A2 (.I(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1992__B1 (.I(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1955__B1 (.I(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1753__B1 (.I(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2003__A2 (.I(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1883__B2 (.I(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1866__A1 (.I(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1816__A2 (.I(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1753__B2 (.I(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1942__A2 (.I(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1788__A3 (.I(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1755__A2 (.I(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1992__A2 (.I(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1962__B1 (.I(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1940__A2 (.I(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1933__B (.I(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1931__B2 (.I(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1787__B2 (.I(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1758__B1 (.I(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2020__A3 (.I(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1931__B1 (.I(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1809__A3 (.I(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1758__B2 (.I(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2709__A2 (.I(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1761__A2 (.I(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1760__A3 (.I(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2832__B2 (.I(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2790__A1 (.I(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2150__A1 (.I(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1766__A2 (.I(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1763__B1 (.I(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2997__B (.I(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1767__A1 (.I(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2704__A1 (.I(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2113__A1 (.I(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1767__A2 (.I(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2031__B2 (.I(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1978__A1 (.I(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1868__A2 (.I(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1783__A2 (.I(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1780__A1 (.I(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1772__A2 (.I(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1982__A2 (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1954__A2 (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1889__A2 (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1775__A2 (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1981__A2 (.I(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1793__A1 (.I(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1781__A1 (.I(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2043__A3 (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1973__A2 (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1955__B2 (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1949__A2 (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1882__A2 (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1870__A1 (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1853__A2 (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1843__A2 (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1840__A3 (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1778__A2 (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1811__A2 (.I(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1779__A2 (.I(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1895__A2 (.I(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1786__A2 (.I(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2483__A1 (.I(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2442__A1 (.I(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2308__B2 (.I(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2271__A1 (.I(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2152__A2 (.I(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1899__A2 (.I(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2000__A2 (.I(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1928__A2 (.I(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1793__A2 (.I(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1797__B1 (.I(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2711__B2 (.I(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2308__A1 (.I(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2205__A1 (.I(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2189__A1 (.I(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2166__A1 (.I(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1901__A2 (.I(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1899__B1 (.I(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2045__B2 (.I(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2035__A1 (.I(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1998__A2 (.I(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1997__A1 (.I(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1928__A1 (.I(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1907__A2 (.I(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1843__A1 (.I(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1842__A2 (.I(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1818__A2 (.I(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1800__A2 (.I(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1890__A1 (.I(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1808__A1 (.I(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2008__A1 (.I(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1803__A2 (.I(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2037__B1 (.I(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1889__B2 (.I(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1872__C (.I(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1806__B1 (.I(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1808__B (.I(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2022__B2 (.I(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2019__A1 (.I(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1953__B2 (.I(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1918__A1 (.I(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1909__A1 (.I(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1854__C (.I(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1837__B (.I(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1828__A1 (.I(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1811__B (.I(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1808__C (.I(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1814__A1 (.I(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1813__A2 (.I(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1814__A2 (.I(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1813__A3 (.I(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2534__A2 (.I(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1834__A2 (.I(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1815__A2 (.I(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2011__B (.I(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1988__A1 (.I(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1973__B1 (.I(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1874__A2 (.I(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1820__A1 (.I(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1830__A1 (.I(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1829__A2 (.I(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2013__A3 (.I(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1931__A3 (.I(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1871__A1 (.I(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1854__A1 (.I(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1841__A2 (.I(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1825__B1 (.I(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1994__A3 (.I(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1871__A2 (.I(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1854__A2 (.I(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1825__B2 (.I(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2024__A2 (.I(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2008__A2 (.I(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1827__A1 (.I(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1830__A2 (.I(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1829__A3 (.I(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2535__I1 (.I(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2487__A2 (.I(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1894__A2 (.I(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1881__B1 (.I(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3079__A1 (.I(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3078__A1 (.I(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3072__A1 (.I(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2957__A1 (.I(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2956__A1 (.I(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2053__A1 (.I(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2052__B2 (.I(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1894__A1 (.I(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1881__B2 (.I(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2349__C2 (.I(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2346__A1 (.I(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2169__C2 (.I(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2154__A1 (.I(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1880__A2 (.I(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1838__A1 (.I(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2037__C (.I(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1944__A2 (.I(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1935__A1 (.I(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1847__A1 (.I(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1978__A2 (.I(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1972__A2 (.I(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1845__A2 (.I(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1847__B1 (.I(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2009__A1 (.I(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1956__A1 (.I(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1915__B2 (.I(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1847__B2 (.I(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1849__A2 (.I(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1848__A3 (.I(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2596__A1 (.I(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2572__A1 (.I(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2397__A1 (.I(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2348__B2 (.I(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2154__B2 (.I(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2147__A1 (.I(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1878__A2 (.I(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1851__A2 (.I(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2396__A1 (.I(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2142__A1 (.I(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1863__A1 (.I(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2396__A2 (.I(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2142__A2 (.I(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1863__A2 (.I(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2625__A1 (.I(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2595__I0 (.I(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2594__A1 (.I(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2442__B2 (.I(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2440__A1 (.I(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1877__A2 (.I(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1864__A2 (.I(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1987__A2 (.I(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1955__A1 (.I(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1950__A1 (.I(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1866__B1 (.I(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2032__C (.I(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1994__A4 (.I(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1983__B (.I(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1868__C (.I(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1875__A2 (.I(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2021__B2 (.I(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1871__B (.I(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1873__A3 (.I(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2347__A2 (.I(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1876__A2 (.I(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2647__I1 (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2644__A1 (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2487__A1 (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2486__A1 (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2440__B2 (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1877__B (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1988__A2 (.I(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1973__B2 (.I(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1885__B1 (.I(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1892__A1 (.I(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1891__A2 (.I(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2034__A2 (.I(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1969__A2 (.I(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1888__A2 (.I(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1892__A2 (.I(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1891__A3 (.I(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2271__B2 (.I(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1897__A2 (.I(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1894__B1 (.I(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2471__A1 (.I(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2397__C (.I(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2173__A1 (.I(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2169__B2 (.I(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2151__A1 (.I(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1898__B1 (.I(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3087__A1 (.I(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2964__A1 (.I(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2939__B2 (.I(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2057__A1 (.I(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2054__B2 (.I(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1898__B2 (.I(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1902__A2 (.I(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1905__I (.I(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3177__A1 (.I(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3175__A1 (.I(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2375__A1 (.I(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2240__A1 (.I(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2028__A1 (.I(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1968__A1 (.I(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1947__A1 (.I(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1923__A1 (.I(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1916__A1 (.I(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1913__A1 (.I(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2854__B2 (.I(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2833__A1 (.I(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2764__A1 (.I(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2216__A1 (.I(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2124__A1 (.I(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2062__A2 (.I(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1917__A2 (.I(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2882__A1 (.I(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2854__A1 (.I(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2785__A1 (.I(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2462__A1 (.I(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2243__A1 (.I(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2215__A1 (.I(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1921__B1 (.I(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1917__B1 (.I(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2980__A1 (.I(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2881__A1 (.I(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2829__A1 (.I(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1924__B1 (.I(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1921__A2 (.I(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3018__A1 (.I(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3009__A1 (.I(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3006__A1 (.I(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2978__A1 (.I(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2853__A1 (.I(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2290__A1 (.I(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1926__A2 (.I(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1924__A2 (.I(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2020__A2 (.I(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1962__A2 (.I(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1931__A2 (.I(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2834__A1 (.I(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2787__A1 (.I(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2725__A1 (.I(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2217__A1 (.I(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2072__A1 (.I(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2064__A2 (.I(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1948__A2 (.I(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2015__A3 (.I(_0987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1941__A3 (.I(_0987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2041__A2 (.I(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1961__A2 (.I(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1951__A2 (.I(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1940__B1 (.I(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2035__A2 (.I(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2032__B (.I(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1952__A1 (.I(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1943__B (.I(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2788__A1 (.I(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2768__A1 (.I(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2705__B2 (.I(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2125__A1 (.I(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2081__A1 (.I(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2061__A2 (.I(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1948__B1 (.I(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2769__A1 (.I(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2731__A1 (.I(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2301__A1 (.I(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2243__A2 (.I(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2073__A1 (.I(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2061__B1 (.I(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2059__B1 (.I(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2127__A2 (.I(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1968__A2 (.I(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2710__B2 (.I(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2386__I0 (.I(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2385__A1 (.I(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2220__A1 (.I(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2058__A2 (.I(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2056__A2 (.I(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1976__A2 (.I(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2732__A1 (.I(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2705__A1 (.I(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2324__A1 (.I(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2258__B2 (.I(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2219__A1 (.I(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2059__A2 (.I(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2058__B1 (.I(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1986__A2 (.I(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2424__A2 (.I(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2302__B2 (.I(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2259__A1 (.I(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2129__B2 (.I(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2084__A1 (.I(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2057__A2 (.I(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2054__B1 (.I(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2005__A1 (.I(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1991__A1 (.I(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2523__A1 (.I(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2466__A1 (.I(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2258__A1 (.I(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2192__A1 (.I(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2085__A1 (.I(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2079__A1 (.I(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2055__A2 (.I(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2053__B1 (.I(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2008__B1 (.I(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2000__B1 (.I(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2007__A2 (.I(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2607__A1 (.I(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2600__A1 (.I(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2562__A1 (.I(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2374__A1 (.I(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2326__A1 (.I(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2177__A1 (.I(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2115__A1 (.I(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2052__A2 (.I(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2050__B1 (.I(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2045__C (.I(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2015__A4 (.I(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2325__A1 (.I(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2018__A1 (.I(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2325__A2 (.I(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2018__A2 (.I(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2194__A1 (.I(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2175__A1 (.I(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2079__B2 (.I(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2053__A2 (.I(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2052__B1 (.I(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2468__A1 (.I(_1077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2380__A1 (.I(_1077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2098__A1 (.I(_1077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2029__I (.I(_1077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2662__A1 (.I(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2661__A1 (.I(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2660__A1 (.I(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2630__A1 (.I(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2629__A1 (.I(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2520__I1 (.I(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2470__A1 (.I(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2439__A1 (.I(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2340__A1 (.I(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2030__I (.I(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2651__A1 (.I(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2636__A1 (.I(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2049__A2 (.I(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2040__A2 (.I(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2375__A2 (.I(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2039__A2 (.I(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2485__A1 (.I(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2339__A1 (.I(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2040__B (.I(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2376__A2 (.I(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2048__A2 (.I(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2425__A1 (.I(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2335__A1 (.I(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2118__A1 (.I(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2104__B (.I(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2050__A2 (.I(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2049__B1 (.I(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3195__A1 (.I(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2110__A1 (.I(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2071__A1 (.I(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3194__A1 (.I(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3192__A1 (.I(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2143__A2 (.I(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2140__A2 (.I(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2116__A1 (.I(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2097__A1 (.I(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2082__A1 (.I(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2076__A3 (.I(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2074__A3 (.I(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2071__A2 (.I(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3197__B (.I(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2139__A1 (.I(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2110__A3 (.I(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2099__A2 (.I(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2082__A2 (.I(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2075__I (.I(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2074__B (.I(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2071__A3 (.I(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2219__A2 (.I(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2217__A2 (.I(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2216__A2 (.I(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2125__A2 (.I(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2123__I (.I(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2081__A2 (.I(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2079__A2 (.I(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2073__A2 (.I(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2072__A2 (.I(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2906__A1 (.I(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2903__A1 (.I(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2759__A1 (.I(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2724__A1 (.I(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2342__A1 (.I(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2130__A1 (.I(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2090__A1 (.I(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2530__A1 (.I(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2528__B (.I(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2434__A1 (.I(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2391__A1 (.I(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2329__A1 (.I(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2328__A1 (.I(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2244__A1 (.I(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2080__A1 (.I(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2128__A2 (.I(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2078__A2 (.I(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2257__I (.I(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2220__A2 (.I(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2085__A2 (.I(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2079__B1 (.I(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2384__A1 (.I(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2330__B2 (.I(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2291__A1 (.I(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2087__A1 (.I(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2241__I (.I(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2129__A2 (.I(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2084__A2 (.I(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2575__A1 (.I(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2564__A1 (.I(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2521__A1 (.I(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2474__A1 (.I(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2470__B1 (.I(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2426__A1 (.I(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2126__A1 (.I(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2086__A1 (.I(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3191__A1 (.I(_1140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3189__A1 (.I(_1140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2099__A1 (.I(_1140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2093__A2 (.I(_1140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2193__A2 (.I(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2165__B (.I(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2108__A3 (.I(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2094__I (.I(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2623__A2 (.I(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2471__A2 (.I(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2441__A3 (.I(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2397__B (.I(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2346__A2 (.I(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2253__B (.I(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2173__A2 (.I(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2113__A2 (.I(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2107__A2 (.I(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2095__A2 (.I(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2732__B (.I(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2336__A1 (.I(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2104__A1 (.I(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3198__A1 (.I(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2116__A2 (.I(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2097__A2 (.I(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2302__B1 (.I(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2098__A2 (.I(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2335__A2 (.I(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2192__A2 (.I(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2175__A2 (.I(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2115__A2 (.I(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2103__I (.I(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3006__A2 (.I(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2978__A2 (.I(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2881__A2 (.I(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2854__A2 (.I(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2833__A2 (.I(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2787__A2 (.I(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2768__A2 (.I(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2731__A2 (.I(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2705__A2 (.I(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2104__C (.I(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2489__A1 (.I(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2114__A2 (.I(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2438__A1 (.I(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2267__S (.I(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2112__I0 (.I(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2734__A1 (.I(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2437__A1 (.I(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2300__A1 (.I(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2112__I1 (.I(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2166__A2 (.I(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2163__A2 (.I(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2149__I (.I(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2136__B (.I(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2117__A2 (.I(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2111__B (.I(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2597__A1 (.I(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2593__A1 (.I(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2572__B2 (.I(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2533__B (.I(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2532__A1 (.I(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2493__A1 (.I(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2488__B2 (.I(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2444__A1 (.I(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2443__A1 (.I(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2112__S (.I(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2732__A2 (.I(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2339__A2 (.I(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2256__I (.I(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2194__A2 (.I(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2177__A2 (.I(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2118__A2 (.I(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2769__B (.I(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2254__A1 (.I(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2207__A1 (.I(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2118__B (.I(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2134__A1 (.I(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2133__A1 (.I(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2466__A2 (.I(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2462__A2 (.I(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2425__A2 (.I(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2385__A2 (.I(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2374__A2 (.I(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2324__A2 (.I(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2290__A2 (.I(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2243__A3 (.I(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2215__A2 (.I(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2124__A2 (.I(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2901__A1 (.I(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2726__A1 (.I(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2558__A1 (.I(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2512__A1 (.I(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2285__A1 (.I(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2239__A1 (.I(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2211__A1 (.I(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2132__A1 (.I(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2695__A2 (.I(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2479__A1 (.I(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2387__B2 (.I(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2292__A2 (.I(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2126__B (.I(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2473__A1 (.I(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2387__A1 (.I(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2302__A1 (.I(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2129__A1 (.I(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2439__A2 (.I(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2377__B1 (.I(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2129__B1 (.I(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2218__A2 (.I(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2130__A2 (.I(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2379__B2 (.I(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2306__S (.I(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2173__B (.I(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2151__A2 (.I(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2137__A1 (.I(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2734__A2 (.I(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2349__A2 (.I(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2348__A2 (.I(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2206__A2 (.I(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2169__A2 (.I(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2154__A2 (.I(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2147__A2 (.I(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3008__A2 (.I(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2734__B1 (.I(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2349__B1 (.I(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2206__B1 (.I(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2169__C1 (.I(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2154__B1 (.I(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2147__B1 (.I(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2734__C2 (.I(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2349__C1 (.I(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2348__B1 (.I(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2169__B1 (.I(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2154__C1 (.I(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2147__C1 (.I(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2536__A1 (.I(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2488__A1 (.I(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2206__B2 (.I(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2169__A1 (.I(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2147__C2 (.I(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2158__A1 (.I(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2156__A1 (.I(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2534__B (.I(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2331__B (.I(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2266__A2 (.I(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2262__A2 (.I(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2200__I (.I(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2198__A3 (.I(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2189__A2 (.I(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2176__A2 (.I(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2152__B (.I(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2150__A2 (.I(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2161__A2 (.I(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2160__A3 (.I(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2153__A2 (.I(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2158__A2 (.I(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2156__A2 (.I(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2183__A1 (.I(_1207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2181__A1 (.I(_1207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2185__A1 (.I(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2171__A1 (.I(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2734__C1 (.I(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2191__A1 (.I(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2167__I0 (.I(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2339__B (.I(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2190__A1 (.I(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2174__A1 (.I(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2167__I1 (.I(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2438__A2 (.I(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2428__A2 (.I(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2378__S (.I(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2190__A2 (.I(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2167__S (.I(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2187__A1 (.I(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2170__A1 (.I(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2187__A2 (.I(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2170__A2 (.I(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2213__A1 (.I(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2212__A1 (.I(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2179__A2 (.I(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2788__B (.I(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2177__B (.I(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2188__A2 (.I(_1225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2178__A2 (.I(_1225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2183__A2 (.I(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2181__A2 (.I(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2518__A1 (.I(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2516__A2 (.I(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2437__A2 (.I(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2379__A2 (.I(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2191__A2 (.I(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2237__A1 (.I(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2196__A1 (.I(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2834__B (.I(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2194__B (.I(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2251__A2 (.I(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2195__A2 (.I(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2484__A2 (.I(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2378__I1 (.I(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2332__I0 (.I(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2199__A2 (.I(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2710__A2 (.I(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2594__A2 (.I(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2487__B (.I(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2486__A2 (.I(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2483__A2 (.I(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2442__A2 (.I(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2440__A2 (.I(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2333__A2 (.I(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2305__A2 (.I(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2201__B (.I(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2856__C2 (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2832__C1 (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2790__C2 (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2771__C1 (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2711__C1 (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2442__B1 (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2440__B1 (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2308__C2 (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2271__C2 (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2205__A2 (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2265__A3 (.I(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2207__A3 (.I(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2249__A2 (.I(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2248__A2 (.I(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2208__A3 (.I(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2229__A1 (.I(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2223__A1 (.I(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2765__A1 (.I(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2682__A1 (.I(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2511__A1 (.I(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2244__A2 (.I(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2235__A1 (.I(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2222__A1 (.I(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2904__A1 (.I(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2683__A1 (.I(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2515__A1 (.I(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2233__A1 (.I(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2221__A1 (.I(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2706__A1 (.I(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2561__A1 (.I(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2557__A1 (.I(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2218__A1 (.I(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2568__A1 (.I(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2567__A1 (.I(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2388__A1 (.I(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2386__S (.I(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2220__B (.I(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2285__A2 (.I(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2239__A2 (.I(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2233__A2 (.I(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2221__A3 (.I(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2695__A1 (.I(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2292__A1 (.I(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2242__A1 (.I(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2662__A2 (.I(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2629__B (.I(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2598__A2 (.I(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2517__A2 (.I(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2516__A3 (.I(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2473__A2 (.I(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2468__A2 (.I(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2424__A3 (.I(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2325__A3 (.I(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2242__A2 (.I(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2785__B (.I(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2423__A1 (.I(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2420__A1 (.I(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2291__A2 (.I(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2289__A1 (.I(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2284__A1 (.I(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2245__A2 (.I(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2734__B2 (.I(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2379__A1 (.I(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2334__A1 (.I(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2253__A2 (.I(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2380__A2 (.I(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2377__A2 (.I(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2340__A2 (.I(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2302__A2 (.I(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2259__A2 (.I(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3018__A2 (.I(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3009__A2 (.I(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2980__A2 (.I(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2882__A2 (.I(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2854__B1 (.I(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2834__A2 (.I(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2788__A2 (.I(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2769__A2 (.I(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2710__B1 (.I(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2258__A2 (.I(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2853__A2 (.I(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2829__A2 (.I(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2785__A2 (.I(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2764__A2 (.I(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2725__A2 (.I(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2705__B1 (.I(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2485__A2 (.I(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2326__A2 (.I(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2301__A2 (.I(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2258__B1 (.I(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2297__A1 (.I(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2273__A1 (.I(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2981__A2 (.I(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2883__A2 (.I(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2856__A2 (.I(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2832__A2 (.I(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2790__A2 (.I(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2771__A2 (.I(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2711__A2 (.I(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2308__A2 (.I(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2271__A2 (.I(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2981__B1 (.I(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2883__B1 (.I(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2856__B1 (.I(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2832__B1 (.I(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2790__B1 (.I(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2771__B1 (.I(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2711__B1 (.I(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2308__B1 (.I(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2271__B1 (.I(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2048__A1 (.I(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1996__A1 (.I(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1986__A1 (.I(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1936__A1 (.I(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1906__I (.I(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1657__I (.I(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1602__A1 (.I(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2689__A1 (.I(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2322__A1 (.I(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1625__A1 (.I(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1619__A1 (.I(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1614__A1 (.I(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1613__A1 (.I(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1610__A1 (.I(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1608__A1 (.I(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1601__I (.I(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2741__A1 (.I(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2295__A1 (.I(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2829__B (.I(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2697__A1 (.I(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2696__A1 (.I(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2421__A1 (.I(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2371__A1 (.I(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2293__A1 (.I(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3177__A2 (.I(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3173__A1 (.I(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1660__A1 (.I(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1658__A2 (.I(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1651__A1 (.I(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1632__A1 (.I(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1629__A1 (.I(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1622__A1 (.I(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1605__A1 (.I(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1602__A2 (.I(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2694__A2 (.I(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2303__A2 (.I(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1760__A1 (.I(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1655__A1 (.I(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1650__A1 (.I(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1603__I (.I(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2727__A2 (.I(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2704__B1 (.I(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2307__A1 (.I(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2347__A1 (.I(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1892__B (.I(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1891__A1 (.I(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1830__B (.I(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1829__A1 (.I(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1786__A1 (.I(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1761__B (.I(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1743__A1 (.I(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1742__B (.I(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1604__I (.I(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2805__A2 (.I(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2321__A2 (.I(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2981__A1 (.I(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2856__C1 (.I(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2305__A1 (.I(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1862__B (.I(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1861__A1 (.I(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1698__B (.I(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1697__A1 (.I(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1669__A2 (.I(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1668__A2 (.I(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1666__A2 (.I(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2636__B2 (.I(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2631__A1 (.I(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2563__A1 (.I(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2562__A2 (.I(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2538__A1 (.I(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2525__A1 (.I(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2519__A1 (.I(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2326__B (.I(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2627__A1 (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2596__B2 (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2535__I0 (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2531__A2 (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2334__A2 (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2332__S (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2341__A2 (.I(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2338__A3 (.I(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2015__A1 (.I(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1983__C (.I(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1934__C (.I(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1790__B (.I(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1695__A1 (.I(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1606__I (.I(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2361__A2 (.I(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2344__A1 (.I(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2343__A1 (.I(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2005__C (.I(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1984__A1 (.I(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1966__B (.I(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1749__B (.I(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1741__C (.I(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1700__I (.I(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1683__I (.I(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1654__A1 (.I(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1649__A1 (.I(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1648__A1 (.I(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2648__A1 (.I(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2625__B2 (.I(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2399__A1 (.I(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2398__A1 (.I(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2395__A1 (.I(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2352__A1 (.I(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2350__A1 (.I(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2623__A1 (.I(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2531__A1 (.I(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2349__B2 (.I(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2348__A1 (.I(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2408__A1 (.I(_1409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2357__A1 (.I(_1409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2355__A1 (.I(_1409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3169__A2 (.I(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3166__A2 (.I(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3163__A1 (.I(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3161__A1 (.I(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1737__A2 (.I(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1724__A2 (.I(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1711__A2 (.I(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1685__A2 (.I(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1625__A2 (.I(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1608__A2 (.I(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2362__A1 (.I(_1415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2360__A1 (.I(_1415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2362__A2 (.I(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2360__A2 (.I(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1971__A2 (.I(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1824__A1 (.I(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1817__A1 (.I(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1750__B (.I(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1730__I0 (.I(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1678__A1 (.I(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1674__I (.I(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1635__I (.I(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1615__A2 (.I(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1611__A1 (.I(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2659__A1 (.I(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2652__A1 (.I(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2599__A1 (.I(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2563__A2 (.I(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2429__A1 (.I(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2404__A1 (.I(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2383__A1 (.I(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3157__A1 (.I(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3154__A1 (.I(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1754__A2 (.I(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1737__A1 (.I(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1685__A1 (.I(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1679__A2 (.I(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1622__A2 (.I(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1610__A2 (.I(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2517__A1 (.I(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2516__A1 (.I(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2377__A1 (.I(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2629__A2 (.I(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2598__A1 (.I(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2424__A1 (.I(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2377__B2 (.I(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2383__B2 (.I(_1438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2382__A1 (.I(_1438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2394__A1 (.I(_1442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2392__A1 (.I(_1442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1965__B2 (.I(_1455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1745__A1 (.I(_1455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1616__A1 (.I(_1455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2494__A1 (.I(_1458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2444__A2 (.I(_1458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2443__B2 (.I(_1458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2401__A2 (.I(_1458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2399__A3 (.I(_1458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3156__I (.I(_1466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1754__A1 (.I(_1466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1724__A1 (.I(_1466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1711__A1 (.I(_1466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1679__A1 (.I(_1466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1619__A2 (.I(_1466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1613__A2 (.I(_1466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1989__A1 (.I(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1971__A1 (.I(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1826__A1 (.I(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1823__A1 (.I(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1756__A1 (.I(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1713__I (.I(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1691__A1 (.I(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1637__I (.I(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1636__A1 (.I(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1615__A1 (.I(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2419__A1 (.I(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2418__A1 (.I(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1817__B (.I(_1488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1751__A1 (.I(_1488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1704__B (.I(_1488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1617__I (.I(_1488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1615__B (.I(_1488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2630__A2 (.I(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2474__A2 (.I(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2426__A2 (.I(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2432__A1 (.I(_1492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2430__A1 (.I(_1492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1982__A1 (.I(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1945__B2 (.I(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1889__A1 (.I(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1827__C (.I(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1806__A1 (.I(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1775__A1 (.I(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1745__A2 (.I(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1682__C (.I(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1616__A2 (.I(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2495__A3 (.I(_1504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2445__A1 (.I(_1504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2645__A1 (.I(_1506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2644__A2 (.I(_1506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2595__S (.I(_1506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2571__S (.I(_1506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2442__C (.I(_1506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1994__A2 (.I(_1510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1648__A4 (.I(_1510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1643__A1 (.I(_1510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2500__A1 (.I(_1511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2449__A1 (.I(_1511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2447__A1 (.I(_1511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2500__A2 (.I(_1512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2449__A2 (.I(_1512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2447__A2 (.I(_1512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2453__A2 (.I(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2452__A2 (.I(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1990__B2 (.I(_1521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1987__A1 (.I(_1521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1930__B (.I(_1521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1867__A2 (.I(_1521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1824__B (.I(_1521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1802__B (.I(_1521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1791__A1 (.I(_1521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1789__B2 (.I(_1521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1644__I (.I(_1521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1618__I (.I(_1521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2462__A3 (.I(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2462__B (.I(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2000__B2 (.I(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1966__A1 (.I(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1882__B (.I(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1772__A1 (.I(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1753__A1 (.I(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1745__B2 (.I(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1735__A1 (.I(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1728__I (.I(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1726__A2 (.I(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1631__A1 (.I(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2936__A1 (.I(_1533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2900__I (.I(_1533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2815__A1 (.I(_1533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2601__A1 (.I(_1534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2520__S (.I(_1534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2470__A2 (.I(_1534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2467__I (.I(_1534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2607__B2 (.I(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2565__A1 (.I(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2469__A1 (.I(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2485__B1 (.I(_1540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2477__A1 (.I(_1540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2476__A1 (.I(_1540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2014__A1 (.I(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1937__A1 (.I(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1930__A1 (.I(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1884__A1 (.I(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1867__A1 (.I(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1746__A1 (.I(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1723__A1 (.I(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1645__A1 (.I(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1640__A1 (.I(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1621__I (.I(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2541__A1 (.I(_1555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2492__A1 (.I(_1555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1998__A1 (.I(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1949__A1 (.I(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1882__A1 (.I(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1840__A1 (.I(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1822__A1 (.I(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1774__A1 (.I(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1701__A1 (.I(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1693__A1 (.I(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1690__A1 (.I(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1628__A1 (.I(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1959__A2 (.I(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1939__A1 (.I(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1824__A2 (.I(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1802__A2 (.I(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1791__A2 (.I(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1774__A3 (.I(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1771__A2 (.I(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1723__A2 (.I(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1688__A2 (.I(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1624__I (.I(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1887__S (.I(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1819__A2 (.I(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1805__A2 (.I(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1800__B (.I(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1747__A2 (.I(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1712__A1 (.I(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1702__A2 (.I(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1701__A2 (.I(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1692__A2 (.I(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1628__A2 (.I(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_0_clk_I (.I(clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3169__A1 (.I(\csTable.address[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3166__A1 (.I(\csTable.address[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3164__A1 (.I(\csTable.address[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1632__A2 (.I(\csTable.address[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1614__A2 (.I(\csTable.address[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3169__A3 (.I(\csTable.address[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3167__A1 (.I(\csTable.address[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1651__A2 (.I(\csTable.address[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1629__A2 (.I(\csTable.address[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3172__A1 (.I(\csTable.address[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3170__A1 (.I(\csTable.address[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1660__A2 (.I(\csTable.address[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1605__A2 (.I(\csTable.address[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(divSel[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(divSel[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(divSel[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(divSel[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3104__B (.I(\freeRunCntr[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2966__I (.I(\freeRunCntr[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2930__A1 (.I(\freeRunCntr[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2926__B1 (.I(\freeRunCntr[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2061__B2 (.I(\freeRunCntr[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2059__B2 (.I(\freeRunCntr[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1900__B2 (.I(\freeRunCntr[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1722__A1 (.I(\freeRunCntr[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1721__B2 (.I(\freeRunCntr[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3121__A1 (.I(\freeRunCntr[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3120__B (.I(\freeRunCntr[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3115__A1 (.I(\freeRunCntr[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2926__A1 (.I(\freeRunCntr[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2061__A1 (.I(\freeRunCntr[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1948__B2 (.I(\freeRunCntr[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1764__I (.I(\freeRunCntr[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1763__A1 (.I(\freeRunCntr[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3117__I (.I(\freeRunCntr[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3022__A1 (.I(\freeRunCntr[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2998__A1 (.I(\freeRunCntr[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2064__A1 (.I(\freeRunCntr[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1948__A1 (.I(\freeRunCntr[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1766__A1 (.I(\freeRunCntr[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1763__B2 (.I(\freeRunCntr[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3135__A1 (.I(\freeRunCntr[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3134__A1 (.I(\freeRunCntr[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3032__A1 (.I(\freeRunCntr[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3028__I (.I(\freeRunCntr[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3025__A1 (.I(\freeRunCntr[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2062__A1 (.I(\freeRunCntr[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1917__A1 (.I(\freeRunCntr[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1670__A1 (.I(\freeRunCntr[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1656__A1 (.I(\freeRunCntr[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3131__I (.I(\freeRunCntr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3031__A1 (.I(\freeRunCntr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3029__A1 (.I(\freeRunCntr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3020__A1 (.I(\freeRunCntr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1921__B2 (.I(\freeRunCntr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1917__B2 (.I(\freeRunCntr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1665__A1 (.I(\freeRunCntr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1656__B2 (.I(\freeRunCntr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3146__A1 (.I(\freeRunCntr[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3145__A1 (.I(\freeRunCntr[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3142__A1 (.I(\freeRunCntr[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3021__A1 (.I(\freeRunCntr[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1924__B2 (.I(\freeRunCntr[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1921__A1 (.I(\freeRunCntr[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1666__B2 (.I(\freeRunCntr[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1665__B2 (.I(\freeRunCntr[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3150__A1 (.I(\freeRunCntr[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3148__A1 (.I(\freeRunCntr[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3021__A2 (.I(\freeRunCntr[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1926__A1 (.I(\freeRunCntr[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1924__A1 (.I(\freeRunCntr[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1669__A1 (.I(\freeRunCntr[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1668__A1 (.I(\freeRunCntr[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1666__A1 (.I(\freeRunCntr[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3048__A1 (.I(\freeRunCntr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3041__A1 (.I(\freeRunCntr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2949__A1 (.I(\freeRunCntr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2945__A2 (.I(\freeRunCntr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2040__C (.I(\freeRunCntr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1877__C (.I(\freeRunCntr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3054__A1 (.I(\freeRunCntr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3047__A1 (.I(\freeRunCntr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2949__B (.I(\freeRunCntr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2945__A1 (.I(\freeRunCntr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2049__A1 (.I(\freeRunCntr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2040__A1 (.I(\freeRunCntr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1877__A1 (.I(\freeRunCntr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1864__A1 (.I(\freeRunCntr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3063__A1 (.I(\freeRunCntr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3062__A1 (.I(\freeRunCntr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2953__A1 (.I(\freeRunCntr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2952__A1 (.I(\freeRunCntr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2050__A1 (.I(\freeRunCntr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2049__B2 (.I(\freeRunCntr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1835__I (.I(\freeRunCntr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3061__A1 (.I(\freeRunCntr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2956__B2 (.I(\freeRunCntr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2954__A1 (.I(\freeRunCntr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2052__A1 (.I(\freeRunCntr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2050__B2 (.I(\freeRunCntr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1881__A1 (.I(\freeRunCntr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1833__I (.I(\freeRunCntr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1832__I (.I(\freeRunCntr[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3077__A1 (.I(\freeRunCntr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2931__I (.I(\freeRunCntr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2055__A1 (.I(\freeRunCntr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2053__B2 (.I(\freeRunCntr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1897__A1 (.I(\freeRunCntr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1894__B2 (.I(\freeRunCntr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3093__A1 (.I(\freeRunCntr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3092__A1 (.I(\freeRunCntr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1899__A1 (.I(\freeRunCntr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1896__I (.I(\freeRunCntr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3090__A1 (.I(\freeRunCntr[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3089__B (.I(\freeRunCntr[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2973__A1 (.I(\freeRunCntr[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2965__B2 (.I(\freeRunCntr[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2058__A1 (.I(\freeRunCntr[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2056__A1 (.I(\freeRunCntr[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1901__A1 (.I(\freeRunCntr[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1899__B2 (.I(\freeRunCntr[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(rst));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2144__A1 (.I(\sigRom.address[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2138__A2 (.I(\sigRom.address[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2110__A2 (.I(\sigRom.address[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2092__I (.I(\sigRom.address[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2076__A2 (.I(\sigRom.address[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2074__A2 (.I(\sigRom.address[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2101__A1 (.I(\sigRom.address[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2100__A1 (.I(\sigRom.address[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2069__I (.I(\sigRom.address[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3083__A2 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3058__A2 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3052__A2 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3039__I (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3036__A2 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3098__A1 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3083__A1 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3074__A1 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3068__A1 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3058__A1 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3052__A1 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3045__A1 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3040__A1 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3036__A1 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3067__I (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3059__A1 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3053__A1 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3046__A1 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3040__A3 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3036__A3 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3044__I (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3040__A4 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3035__I (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output6_I (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output8_I (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3209__RN (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3204__RN (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3202__RN (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3201__RN (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3223__RN (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3222__RN (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3221__RN (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3220__RN (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3217__RN (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3203__RN (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3231__RN (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3230__RN (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3226__RN (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3216__RN (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3208__RN (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3215__RN (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3214__RN (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3207__RN (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3206__RN (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3205__RN (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3232__RN (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3233__RN (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout10_I (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3229__RN (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3228__RN (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3227__RN (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3225__RN (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3224__RN (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3219__RN (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3218__RN (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout11_I (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3210__RN (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3211__RN (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3212__RN (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3213__RN (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout9_I (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_2_3__f_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_2_2__f_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_2_1__f_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_2_0__f_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3202__CLK (.I(clknet_2_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3203__CLK (.I(clknet_2_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3205__CLK (.I(clknet_2_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3217__CLK (.I(clknet_2_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3220__CLK (.I(clknet_2_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3221__CLK (.I(clknet_2_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3222__CLK (.I(clknet_2_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3223__CLK (.I(clknet_2_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3201__CLK (.I(clknet_2_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3204__CLK (.I(clknet_2_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3209__CLK (.I(clknet_2_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3210__CLK (.I(clknet_2_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3211__CLK (.I(clknet_2_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3212__CLK (.I(clknet_2_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3213__CLK (.I(clknet_2_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3214__CLK (.I(clknet_2_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3207__CLK (.I(clknet_2_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3218__CLK (.I(clknet_2_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3219__CLK (.I(clknet_2_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3224__CLK (.I(clknet_2_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3225__CLK (.I(clknet_2_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3226__CLK (.I(clknet_2_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3227__CLK (.I(clknet_2_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3228__CLK (.I(clknet_2_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3229__CLK (.I(clknet_2_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3206__CLK (.I(clknet_2_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3208__CLK (.I(clknet_2_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3215__CLK (.I(clknet_2_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3216__CLK (.I(clknet_2_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3230__CLK (.I(clknet_2_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3231__CLK (.I(clknet_2_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3232__CLK (.I(clknet_2_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3233__CLK (.I(clknet_2_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_512 ();
endmodule

