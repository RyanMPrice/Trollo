VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO DiffDigota
  CLASS BLOCK ;
  FOREIGN DiffDigota ;
  ORIGIN 0.000 0.000 ;
  SIZE 80.000 BY 80.000 ;
  PIN INmb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 24.080 0.000 24.640 4.000 ;
    END
  END INmb
  PIN INpb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 8.400 0.000 8.960 4.000 ;
    END
  END INpb
  PIN OUTm
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 55.440 0.000 56.000 4.000 ;
    END
  END OUTm
  PIN OUTp
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 39.760 0.000 40.320 4.000 ;
    END
  END OUTp
  PIN cmnmos
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 59.360 4.000 59.920 ;
    END
  END cmnmos
  PIN cmpmos
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 19.600 4.000 20.160 ;
    END
  END cmpmos
  PIN oe
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 71.120 0.000 71.680 4.000 ;
    END
  END oe
  PIN omnmos
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 68.880 76.000 69.440 80.000 ;
    END
  END omnmos
  PIN ompmos
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 49.280 76.000 49.840 80.000 ;
    END
  END ompmos
  PIN opnmos
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 29.680 76.000 30.240 80.000 ;
    END
  END opnmos
  PIN oppmos
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 10.080 76.000 10.640 80.000 ;
    END
  END oppmos
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 14.180 15.380 15.780 63.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 30.700 15.380 32.300 63.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 47.220 15.380 48.820 63.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 63.740 15.380 65.340 63.020 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 22.440 15.380 24.040 63.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 38.960 15.380 40.560 63.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 55.480 15.380 57.080 63.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 72.000 15.380 73.600 63.020 ;
    END
  END vss
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 73.600 63.020 ;
      LAYER Metal2 ;
        RECT 8.540 75.700 9.780 76.000 ;
        RECT 10.940 75.700 29.380 76.000 ;
        RECT 30.540 75.700 48.980 76.000 ;
        RECT 50.140 75.700 68.580 76.000 ;
        RECT 69.740 75.700 73.460 76.000 ;
        RECT 8.540 4.300 73.460 75.700 ;
        RECT 9.260 3.500 23.780 4.300 ;
        RECT 24.940 3.500 39.460 4.300 ;
        RECT 40.620 3.500 55.140 4.300 ;
        RECT 56.300 3.500 70.820 4.300 ;
        RECT 71.980 3.500 73.460 4.300 ;
      LAYER Metal3 ;
        RECT 4.000 60.220 73.510 62.860 ;
        RECT 4.300 59.060 73.510 60.220 ;
        RECT 4.000 20.460 73.510 59.060 ;
        RECT 4.300 19.300 73.510 20.460 ;
        RECT 4.000 15.540 73.510 19.300 ;
  END
END DiffDigota
END LIBRARY

