magic
tech gf180mcuC
magscale 1 5
timestamp 1670260475
<< metal1 >>
rect 672 4325 5320 4342
rect 672 4299 1188 4325
rect 1214 4299 1240 4325
rect 1266 4299 1292 4325
rect 1318 4299 2350 4325
rect 2376 4299 2402 4325
rect 2428 4299 2454 4325
rect 2480 4299 3512 4325
rect 3538 4299 3564 4325
rect 3590 4299 3616 4325
rect 3642 4299 4674 4325
rect 4700 4299 4726 4325
rect 4752 4299 4778 4325
rect 4804 4299 5320 4325
rect 672 4282 5320 4299
rect 3425 4159 3431 4185
rect 3457 4159 3463 4185
rect 3089 4103 3095 4129
rect 3121 4103 3127 4129
rect 672 3933 5400 3950
rect 672 3907 1769 3933
rect 1795 3907 1821 3933
rect 1847 3907 1873 3933
rect 1899 3907 2931 3933
rect 2957 3907 2983 3933
rect 3009 3907 3035 3933
rect 3061 3907 4093 3933
rect 4119 3907 4145 3933
rect 4171 3907 4197 3933
rect 4223 3907 5255 3933
rect 5281 3907 5307 3933
rect 5333 3907 5359 3933
rect 5385 3907 5400 3933
rect 672 3890 5400 3907
rect 672 3541 5320 3558
rect 672 3515 1188 3541
rect 1214 3515 1240 3541
rect 1266 3515 1292 3541
rect 1318 3515 2350 3541
rect 2376 3515 2402 3541
rect 2428 3515 2454 3541
rect 2480 3515 3512 3541
rect 3538 3515 3564 3541
rect 3590 3515 3616 3541
rect 3642 3515 4674 3541
rect 4700 3515 4726 3541
rect 4752 3515 4778 3541
rect 4804 3515 5320 3541
rect 672 3498 5320 3515
rect 1633 3375 1639 3401
rect 1665 3375 1671 3401
rect 2871 3289 2897 3295
rect 961 3263 967 3289
rect 993 3263 999 3289
rect 2871 3257 2897 3263
rect 3039 3289 3065 3295
rect 3039 3257 3065 3263
rect 672 3149 5400 3166
rect 672 3123 1769 3149
rect 1795 3123 1821 3149
rect 1847 3123 1873 3149
rect 1899 3123 2931 3149
rect 2957 3123 2983 3149
rect 3009 3123 3035 3149
rect 3061 3123 4093 3149
rect 4119 3123 4145 3149
rect 4171 3123 4197 3149
rect 4223 3123 5255 3149
rect 5281 3123 5307 3149
rect 5333 3123 5359 3149
rect 5385 3123 5400 3149
rect 672 3106 5400 3123
rect 3313 3039 3319 3065
rect 3345 3039 3351 3065
rect 911 3009 937 3015
rect 2703 3009 2729 3015
rect 2081 2983 2087 3009
rect 2113 2983 2119 3009
rect 911 2977 937 2983
rect 2703 2977 2729 2983
rect 3151 2953 3177 2959
rect 3151 2921 3177 2927
rect 3039 2897 3065 2903
rect 1913 2871 1919 2897
rect 1945 2871 1951 2897
rect 3039 2865 3065 2871
rect 672 2757 5320 2774
rect 672 2731 1188 2757
rect 1214 2731 1240 2757
rect 1266 2731 1292 2757
rect 1318 2731 2350 2757
rect 2376 2731 2402 2757
rect 2428 2731 2454 2757
rect 2480 2731 3512 2757
rect 3538 2731 3564 2757
rect 3590 2731 3616 2757
rect 3642 2731 4674 2757
rect 4700 2731 4726 2757
rect 4752 2731 4778 2757
rect 4804 2731 5320 2757
rect 672 2714 5320 2731
rect 2311 2673 2337 2679
rect 2311 2641 2337 2647
rect 2367 2561 2393 2567
rect 2367 2529 2393 2535
rect 672 2365 5400 2382
rect 672 2339 1769 2365
rect 1795 2339 1821 2365
rect 1847 2339 1873 2365
rect 1899 2339 2931 2365
rect 2957 2339 2983 2365
rect 3009 2339 3035 2365
rect 3061 2339 4093 2365
rect 4119 2339 4145 2365
rect 4171 2339 4197 2365
rect 4223 2339 5255 2365
rect 5281 2339 5307 2365
rect 5333 2339 5359 2365
rect 5385 2339 5400 2365
rect 672 2322 5400 2339
rect 672 1973 5320 1990
rect 672 1947 1188 1973
rect 1214 1947 1240 1973
rect 1266 1947 1292 1973
rect 1318 1947 2350 1973
rect 2376 1947 2402 1973
rect 2428 1947 2454 1973
rect 2480 1947 3512 1973
rect 3538 1947 3564 1973
rect 3590 1947 3616 1973
rect 3642 1947 4674 1973
rect 4700 1947 4726 1973
rect 4752 1947 4778 1973
rect 4804 1947 5320 1973
rect 672 1930 5320 1947
rect 3089 1807 3095 1833
rect 3121 1807 3127 1833
rect 2871 1721 2897 1727
rect 3593 1695 3599 1721
rect 3625 1695 3631 1721
rect 2871 1689 2897 1695
rect 672 1581 5400 1598
rect 672 1555 1769 1581
rect 1795 1555 1821 1581
rect 1847 1555 1873 1581
rect 1899 1555 2931 1581
rect 2957 1555 2983 1581
rect 3009 1555 3035 1581
rect 3061 1555 4093 1581
rect 4119 1555 4145 1581
rect 4171 1555 4197 1581
rect 4223 1555 5255 1581
rect 5281 1555 5307 1581
rect 5333 1555 5359 1581
rect 5385 1555 5400 1581
rect 672 1538 5400 1555
<< via1 >>
rect 1188 4299 1214 4325
rect 1240 4299 1266 4325
rect 1292 4299 1318 4325
rect 2350 4299 2376 4325
rect 2402 4299 2428 4325
rect 2454 4299 2480 4325
rect 3512 4299 3538 4325
rect 3564 4299 3590 4325
rect 3616 4299 3642 4325
rect 4674 4299 4700 4325
rect 4726 4299 4752 4325
rect 4778 4299 4804 4325
rect 3431 4159 3457 4185
rect 3095 4103 3121 4129
rect 1769 3907 1795 3933
rect 1821 3907 1847 3933
rect 1873 3907 1899 3933
rect 2931 3907 2957 3933
rect 2983 3907 3009 3933
rect 3035 3907 3061 3933
rect 4093 3907 4119 3933
rect 4145 3907 4171 3933
rect 4197 3907 4223 3933
rect 5255 3907 5281 3933
rect 5307 3907 5333 3933
rect 5359 3907 5385 3933
rect 1188 3515 1214 3541
rect 1240 3515 1266 3541
rect 1292 3515 1318 3541
rect 2350 3515 2376 3541
rect 2402 3515 2428 3541
rect 2454 3515 2480 3541
rect 3512 3515 3538 3541
rect 3564 3515 3590 3541
rect 3616 3515 3642 3541
rect 4674 3515 4700 3541
rect 4726 3515 4752 3541
rect 4778 3515 4804 3541
rect 1639 3375 1665 3401
rect 967 3263 993 3289
rect 2871 3263 2897 3289
rect 3039 3263 3065 3289
rect 1769 3123 1795 3149
rect 1821 3123 1847 3149
rect 1873 3123 1899 3149
rect 2931 3123 2957 3149
rect 2983 3123 3009 3149
rect 3035 3123 3061 3149
rect 4093 3123 4119 3149
rect 4145 3123 4171 3149
rect 4197 3123 4223 3149
rect 5255 3123 5281 3149
rect 5307 3123 5333 3149
rect 5359 3123 5385 3149
rect 3319 3039 3345 3065
rect 911 2983 937 3009
rect 2087 2983 2113 3009
rect 2703 2983 2729 3009
rect 3151 2927 3177 2953
rect 1919 2871 1945 2897
rect 3039 2871 3065 2897
rect 1188 2731 1214 2757
rect 1240 2731 1266 2757
rect 1292 2731 1318 2757
rect 2350 2731 2376 2757
rect 2402 2731 2428 2757
rect 2454 2731 2480 2757
rect 3512 2731 3538 2757
rect 3564 2731 3590 2757
rect 3616 2731 3642 2757
rect 4674 2731 4700 2757
rect 4726 2731 4752 2757
rect 4778 2731 4804 2757
rect 2311 2647 2337 2673
rect 2367 2535 2393 2561
rect 1769 2339 1795 2365
rect 1821 2339 1847 2365
rect 1873 2339 1899 2365
rect 2931 2339 2957 2365
rect 2983 2339 3009 2365
rect 3035 2339 3061 2365
rect 4093 2339 4119 2365
rect 4145 2339 4171 2365
rect 4197 2339 4223 2365
rect 5255 2339 5281 2365
rect 5307 2339 5333 2365
rect 5359 2339 5385 2365
rect 1188 1947 1214 1973
rect 1240 1947 1266 1973
rect 1292 1947 1318 1973
rect 2350 1947 2376 1973
rect 2402 1947 2428 1973
rect 2454 1947 2480 1973
rect 3512 1947 3538 1973
rect 3564 1947 3590 1973
rect 3616 1947 3642 1973
rect 4674 1947 4700 1973
rect 4726 1947 4752 1973
rect 4778 1947 4804 1973
rect 3095 1807 3121 1833
rect 2871 1695 2897 1721
rect 3599 1695 3625 1721
rect 1769 1555 1795 1581
rect 1821 1555 1847 1581
rect 1873 1555 1899 1581
rect 2931 1555 2957 1581
rect 2983 1555 3009 1581
rect 3035 1555 3061 1581
rect 4093 1555 4119 1581
rect 4145 1555 4171 1581
rect 4197 1555 4223 1581
rect 5255 1555 5281 1581
rect 5307 1555 5333 1581
rect 5359 1555 5385 1581
<< metal2 >>
rect 2968 5600 3024 6000
rect 1187 4326 1319 4331
rect 1215 4298 1239 4326
rect 1267 4298 1291 4326
rect 1187 4293 1319 4298
rect 2349 4326 2481 4331
rect 2377 4298 2401 4326
rect 2429 4298 2453 4326
rect 2349 4293 2481 4298
rect 2982 4186 3010 5600
rect 3511 4326 3643 4331
rect 3539 4298 3563 4326
rect 3591 4298 3615 4326
rect 3511 4293 3643 4298
rect 4673 4326 4805 4331
rect 4701 4298 4725 4326
rect 4753 4298 4777 4326
rect 4673 4293 4805 4298
rect 2982 4153 3010 4158
rect 3430 4186 3458 4191
rect 3430 4139 3458 4158
rect 3094 4129 3122 4135
rect 3094 4103 3095 4129
rect 3121 4103 3122 4129
rect 1768 3934 1900 3939
rect 1796 3906 1820 3934
rect 1848 3906 1872 3934
rect 1768 3901 1900 3906
rect 2930 3934 3062 3939
rect 2958 3906 2982 3934
rect 3010 3906 3034 3934
rect 2930 3901 3062 3906
rect 1187 3542 1319 3547
rect 1215 3514 1239 3542
rect 1267 3514 1291 3542
rect 1187 3509 1319 3514
rect 2349 3542 2481 3547
rect 2377 3514 2401 3542
rect 2429 3514 2453 3542
rect 2349 3509 2481 3514
rect 1638 3402 1666 3407
rect 1638 3401 1722 3402
rect 1638 3375 1639 3401
rect 1665 3375 1722 3401
rect 1638 3374 1722 3375
rect 1638 3369 1666 3374
rect 966 3290 994 3295
rect 910 3289 994 3290
rect 910 3263 967 3289
rect 993 3263 994 3289
rect 910 3262 994 3263
rect 910 3010 938 3262
rect 966 3257 994 3262
rect 1694 3234 1722 3374
rect 2870 3289 2898 3295
rect 2870 3263 2871 3289
rect 2897 3263 2898 3289
rect 1694 3206 2114 3234
rect 1768 3150 1900 3155
rect 1796 3122 1820 3150
rect 1848 3122 1872 3150
rect 1768 3117 1900 3122
rect 910 2963 938 2982
rect 2086 3009 2114 3206
rect 2870 3066 2898 3263
rect 3038 3290 3066 3295
rect 3094 3290 3122 4103
rect 4092 3934 4224 3939
rect 4120 3906 4144 3934
rect 4172 3906 4196 3934
rect 4092 3901 4224 3906
rect 5254 3934 5386 3939
rect 5282 3906 5306 3934
rect 5334 3906 5358 3934
rect 5254 3901 5386 3906
rect 3511 3542 3643 3547
rect 3539 3514 3563 3542
rect 3591 3514 3615 3542
rect 3511 3509 3643 3514
rect 4673 3542 4805 3547
rect 4701 3514 4725 3542
rect 4753 3514 4777 3542
rect 4673 3509 4805 3514
rect 3038 3289 3122 3290
rect 3038 3263 3039 3289
rect 3065 3263 3122 3289
rect 3038 3262 3122 3263
rect 3038 3257 3066 3262
rect 2930 3150 3062 3155
rect 2958 3122 2982 3150
rect 3010 3122 3034 3150
rect 2930 3117 3062 3122
rect 4092 3150 4224 3155
rect 4120 3122 4144 3150
rect 4172 3122 4196 3150
rect 4092 3117 4224 3122
rect 5254 3150 5386 3155
rect 5282 3122 5306 3150
rect 5334 3122 5358 3150
rect 5254 3117 5386 3122
rect 3318 3066 3346 3071
rect 2870 3065 3346 3066
rect 2870 3039 3319 3065
rect 3345 3039 3346 3065
rect 2870 3038 3346 3039
rect 3318 3033 3346 3038
rect 2086 2983 2087 3009
rect 2113 2983 2114 3009
rect 2086 2977 2114 2983
rect 2702 3010 2730 3015
rect 2702 3009 3178 3010
rect 2702 2983 2703 3009
rect 2729 2983 3178 3009
rect 2702 2982 3178 2983
rect 2702 2977 2730 2982
rect 3150 2953 3178 2982
rect 3150 2927 3151 2953
rect 3177 2927 3178 2953
rect 3150 2921 3178 2927
rect 1918 2898 1946 2903
rect 3038 2898 3066 2903
rect 1918 2897 2282 2898
rect 1918 2871 1919 2897
rect 1945 2871 2282 2897
rect 1918 2870 2282 2871
rect 1918 2865 1946 2870
rect 1187 2758 1319 2763
rect 1215 2730 1239 2758
rect 1267 2730 1291 2758
rect 1187 2725 1319 2730
rect 2254 2674 2282 2870
rect 3038 2897 3122 2898
rect 3038 2871 3039 2897
rect 3065 2871 3122 2897
rect 3038 2870 3122 2871
rect 3038 2865 3066 2870
rect 2349 2758 2481 2763
rect 2377 2730 2401 2758
rect 2429 2730 2453 2758
rect 2349 2725 2481 2730
rect 2310 2674 2338 2679
rect 2254 2673 2338 2674
rect 2254 2647 2311 2673
rect 2337 2647 2338 2673
rect 2254 2646 2338 2647
rect 2310 2641 2338 2646
rect 2366 2562 2394 2567
rect 2366 2515 2394 2534
rect 3094 2562 3122 2870
rect 3511 2758 3643 2763
rect 3539 2730 3563 2758
rect 3591 2730 3615 2758
rect 3511 2725 3643 2730
rect 4673 2758 4805 2763
rect 4701 2730 4725 2758
rect 4753 2730 4777 2758
rect 4673 2725 4805 2730
rect 1768 2366 1900 2371
rect 1796 2338 1820 2366
rect 1848 2338 1872 2366
rect 1768 2333 1900 2338
rect 2930 2366 3062 2371
rect 2958 2338 2982 2366
rect 3010 2338 3034 2366
rect 2930 2333 3062 2338
rect 1187 1974 1319 1979
rect 1215 1946 1239 1974
rect 1267 1946 1291 1974
rect 1187 1941 1319 1946
rect 2349 1974 2481 1979
rect 2377 1946 2401 1974
rect 2429 1946 2453 1974
rect 2349 1941 2481 1946
rect 3094 1833 3122 2534
rect 4092 2366 4224 2371
rect 4120 2338 4144 2366
rect 4172 2338 4196 2366
rect 4092 2333 4224 2338
rect 5254 2366 5386 2371
rect 5282 2338 5306 2366
rect 5334 2338 5358 2366
rect 5254 2333 5386 2338
rect 3511 1974 3643 1979
rect 3539 1946 3563 1974
rect 3591 1946 3615 1974
rect 3511 1941 3643 1946
rect 4673 1974 4805 1979
rect 4701 1946 4725 1974
rect 4753 1946 4777 1974
rect 4673 1941 4805 1946
rect 3094 1807 3095 1833
rect 3121 1807 3122 1833
rect 3094 1801 3122 1807
rect 2870 1722 2898 1727
rect 1768 1582 1900 1587
rect 1796 1554 1820 1582
rect 1848 1554 1872 1582
rect 1768 1549 1900 1554
rect 2870 1162 2898 1694
rect 3598 1722 3626 1727
rect 3598 1675 3626 1694
rect 2930 1582 3062 1587
rect 2958 1554 2982 1582
rect 3010 1554 3034 1582
rect 2930 1549 3062 1554
rect 4092 1582 4224 1587
rect 4120 1554 4144 1582
rect 4172 1554 4196 1582
rect 4092 1549 4224 1554
rect 5254 1582 5386 1587
rect 5282 1554 5306 1582
rect 5334 1554 5358 1582
rect 5254 1549 5386 1554
rect 2870 1134 3010 1162
rect 2982 400 3010 1134
rect 2968 0 3024 400
<< via2 >>
rect 1187 4325 1215 4326
rect 1187 4299 1188 4325
rect 1188 4299 1214 4325
rect 1214 4299 1215 4325
rect 1187 4298 1215 4299
rect 1239 4325 1267 4326
rect 1239 4299 1240 4325
rect 1240 4299 1266 4325
rect 1266 4299 1267 4325
rect 1239 4298 1267 4299
rect 1291 4325 1319 4326
rect 1291 4299 1292 4325
rect 1292 4299 1318 4325
rect 1318 4299 1319 4325
rect 1291 4298 1319 4299
rect 2349 4325 2377 4326
rect 2349 4299 2350 4325
rect 2350 4299 2376 4325
rect 2376 4299 2377 4325
rect 2349 4298 2377 4299
rect 2401 4325 2429 4326
rect 2401 4299 2402 4325
rect 2402 4299 2428 4325
rect 2428 4299 2429 4325
rect 2401 4298 2429 4299
rect 2453 4325 2481 4326
rect 2453 4299 2454 4325
rect 2454 4299 2480 4325
rect 2480 4299 2481 4325
rect 2453 4298 2481 4299
rect 3511 4325 3539 4326
rect 3511 4299 3512 4325
rect 3512 4299 3538 4325
rect 3538 4299 3539 4325
rect 3511 4298 3539 4299
rect 3563 4325 3591 4326
rect 3563 4299 3564 4325
rect 3564 4299 3590 4325
rect 3590 4299 3591 4325
rect 3563 4298 3591 4299
rect 3615 4325 3643 4326
rect 3615 4299 3616 4325
rect 3616 4299 3642 4325
rect 3642 4299 3643 4325
rect 3615 4298 3643 4299
rect 4673 4325 4701 4326
rect 4673 4299 4674 4325
rect 4674 4299 4700 4325
rect 4700 4299 4701 4325
rect 4673 4298 4701 4299
rect 4725 4325 4753 4326
rect 4725 4299 4726 4325
rect 4726 4299 4752 4325
rect 4752 4299 4753 4325
rect 4725 4298 4753 4299
rect 4777 4325 4805 4326
rect 4777 4299 4778 4325
rect 4778 4299 4804 4325
rect 4804 4299 4805 4325
rect 4777 4298 4805 4299
rect 2982 4158 3010 4186
rect 3430 4185 3458 4186
rect 3430 4159 3431 4185
rect 3431 4159 3457 4185
rect 3457 4159 3458 4185
rect 3430 4158 3458 4159
rect 1768 3933 1796 3934
rect 1768 3907 1769 3933
rect 1769 3907 1795 3933
rect 1795 3907 1796 3933
rect 1768 3906 1796 3907
rect 1820 3933 1848 3934
rect 1820 3907 1821 3933
rect 1821 3907 1847 3933
rect 1847 3907 1848 3933
rect 1820 3906 1848 3907
rect 1872 3933 1900 3934
rect 1872 3907 1873 3933
rect 1873 3907 1899 3933
rect 1899 3907 1900 3933
rect 1872 3906 1900 3907
rect 2930 3933 2958 3934
rect 2930 3907 2931 3933
rect 2931 3907 2957 3933
rect 2957 3907 2958 3933
rect 2930 3906 2958 3907
rect 2982 3933 3010 3934
rect 2982 3907 2983 3933
rect 2983 3907 3009 3933
rect 3009 3907 3010 3933
rect 2982 3906 3010 3907
rect 3034 3933 3062 3934
rect 3034 3907 3035 3933
rect 3035 3907 3061 3933
rect 3061 3907 3062 3933
rect 3034 3906 3062 3907
rect 1187 3541 1215 3542
rect 1187 3515 1188 3541
rect 1188 3515 1214 3541
rect 1214 3515 1215 3541
rect 1187 3514 1215 3515
rect 1239 3541 1267 3542
rect 1239 3515 1240 3541
rect 1240 3515 1266 3541
rect 1266 3515 1267 3541
rect 1239 3514 1267 3515
rect 1291 3541 1319 3542
rect 1291 3515 1292 3541
rect 1292 3515 1318 3541
rect 1318 3515 1319 3541
rect 1291 3514 1319 3515
rect 2349 3541 2377 3542
rect 2349 3515 2350 3541
rect 2350 3515 2376 3541
rect 2376 3515 2377 3541
rect 2349 3514 2377 3515
rect 2401 3541 2429 3542
rect 2401 3515 2402 3541
rect 2402 3515 2428 3541
rect 2428 3515 2429 3541
rect 2401 3514 2429 3515
rect 2453 3541 2481 3542
rect 2453 3515 2454 3541
rect 2454 3515 2480 3541
rect 2480 3515 2481 3541
rect 2453 3514 2481 3515
rect 1768 3149 1796 3150
rect 1768 3123 1769 3149
rect 1769 3123 1795 3149
rect 1795 3123 1796 3149
rect 1768 3122 1796 3123
rect 1820 3149 1848 3150
rect 1820 3123 1821 3149
rect 1821 3123 1847 3149
rect 1847 3123 1848 3149
rect 1820 3122 1848 3123
rect 1872 3149 1900 3150
rect 1872 3123 1873 3149
rect 1873 3123 1899 3149
rect 1899 3123 1900 3149
rect 1872 3122 1900 3123
rect 910 3009 938 3010
rect 910 2983 911 3009
rect 911 2983 937 3009
rect 937 2983 938 3009
rect 910 2982 938 2983
rect 4092 3933 4120 3934
rect 4092 3907 4093 3933
rect 4093 3907 4119 3933
rect 4119 3907 4120 3933
rect 4092 3906 4120 3907
rect 4144 3933 4172 3934
rect 4144 3907 4145 3933
rect 4145 3907 4171 3933
rect 4171 3907 4172 3933
rect 4144 3906 4172 3907
rect 4196 3933 4224 3934
rect 4196 3907 4197 3933
rect 4197 3907 4223 3933
rect 4223 3907 4224 3933
rect 4196 3906 4224 3907
rect 5254 3933 5282 3934
rect 5254 3907 5255 3933
rect 5255 3907 5281 3933
rect 5281 3907 5282 3933
rect 5254 3906 5282 3907
rect 5306 3933 5334 3934
rect 5306 3907 5307 3933
rect 5307 3907 5333 3933
rect 5333 3907 5334 3933
rect 5306 3906 5334 3907
rect 5358 3933 5386 3934
rect 5358 3907 5359 3933
rect 5359 3907 5385 3933
rect 5385 3907 5386 3933
rect 5358 3906 5386 3907
rect 3511 3541 3539 3542
rect 3511 3515 3512 3541
rect 3512 3515 3538 3541
rect 3538 3515 3539 3541
rect 3511 3514 3539 3515
rect 3563 3541 3591 3542
rect 3563 3515 3564 3541
rect 3564 3515 3590 3541
rect 3590 3515 3591 3541
rect 3563 3514 3591 3515
rect 3615 3541 3643 3542
rect 3615 3515 3616 3541
rect 3616 3515 3642 3541
rect 3642 3515 3643 3541
rect 3615 3514 3643 3515
rect 4673 3541 4701 3542
rect 4673 3515 4674 3541
rect 4674 3515 4700 3541
rect 4700 3515 4701 3541
rect 4673 3514 4701 3515
rect 4725 3541 4753 3542
rect 4725 3515 4726 3541
rect 4726 3515 4752 3541
rect 4752 3515 4753 3541
rect 4725 3514 4753 3515
rect 4777 3541 4805 3542
rect 4777 3515 4778 3541
rect 4778 3515 4804 3541
rect 4804 3515 4805 3541
rect 4777 3514 4805 3515
rect 2930 3149 2958 3150
rect 2930 3123 2931 3149
rect 2931 3123 2957 3149
rect 2957 3123 2958 3149
rect 2930 3122 2958 3123
rect 2982 3149 3010 3150
rect 2982 3123 2983 3149
rect 2983 3123 3009 3149
rect 3009 3123 3010 3149
rect 2982 3122 3010 3123
rect 3034 3149 3062 3150
rect 3034 3123 3035 3149
rect 3035 3123 3061 3149
rect 3061 3123 3062 3149
rect 3034 3122 3062 3123
rect 4092 3149 4120 3150
rect 4092 3123 4093 3149
rect 4093 3123 4119 3149
rect 4119 3123 4120 3149
rect 4092 3122 4120 3123
rect 4144 3149 4172 3150
rect 4144 3123 4145 3149
rect 4145 3123 4171 3149
rect 4171 3123 4172 3149
rect 4144 3122 4172 3123
rect 4196 3149 4224 3150
rect 4196 3123 4197 3149
rect 4197 3123 4223 3149
rect 4223 3123 4224 3149
rect 4196 3122 4224 3123
rect 5254 3149 5282 3150
rect 5254 3123 5255 3149
rect 5255 3123 5281 3149
rect 5281 3123 5282 3149
rect 5254 3122 5282 3123
rect 5306 3149 5334 3150
rect 5306 3123 5307 3149
rect 5307 3123 5333 3149
rect 5333 3123 5334 3149
rect 5306 3122 5334 3123
rect 5358 3149 5386 3150
rect 5358 3123 5359 3149
rect 5359 3123 5385 3149
rect 5385 3123 5386 3149
rect 5358 3122 5386 3123
rect 1187 2757 1215 2758
rect 1187 2731 1188 2757
rect 1188 2731 1214 2757
rect 1214 2731 1215 2757
rect 1187 2730 1215 2731
rect 1239 2757 1267 2758
rect 1239 2731 1240 2757
rect 1240 2731 1266 2757
rect 1266 2731 1267 2757
rect 1239 2730 1267 2731
rect 1291 2757 1319 2758
rect 1291 2731 1292 2757
rect 1292 2731 1318 2757
rect 1318 2731 1319 2757
rect 1291 2730 1319 2731
rect 2349 2757 2377 2758
rect 2349 2731 2350 2757
rect 2350 2731 2376 2757
rect 2376 2731 2377 2757
rect 2349 2730 2377 2731
rect 2401 2757 2429 2758
rect 2401 2731 2402 2757
rect 2402 2731 2428 2757
rect 2428 2731 2429 2757
rect 2401 2730 2429 2731
rect 2453 2757 2481 2758
rect 2453 2731 2454 2757
rect 2454 2731 2480 2757
rect 2480 2731 2481 2757
rect 2453 2730 2481 2731
rect 2366 2561 2394 2562
rect 2366 2535 2367 2561
rect 2367 2535 2393 2561
rect 2393 2535 2394 2561
rect 2366 2534 2394 2535
rect 3511 2757 3539 2758
rect 3511 2731 3512 2757
rect 3512 2731 3538 2757
rect 3538 2731 3539 2757
rect 3511 2730 3539 2731
rect 3563 2757 3591 2758
rect 3563 2731 3564 2757
rect 3564 2731 3590 2757
rect 3590 2731 3591 2757
rect 3563 2730 3591 2731
rect 3615 2757 3643 2758
rect 3615 2731 3616 2757
rect 3616 2731 3642 2757
rect 3642 2731 3643 2757
rect 3615 2730 3643 2731
rect 4673 2757 4701 2758
rect 4673 2731 4674 2757
rect 4674 2731 4700 2757
rect 4700 2731 4701 2757
rect 4673 2730 4701 2731
rect 4725 2757 4753 2758
rect 4725 2731 4726 2757
rect 4726 2731 4752 2757
rect 4752 2731 4753 2757
rect 4725 2730 4753 2731
rect 4777 2757 4805 2758
rect 4777 2731 4778 2757
rect 4778 2731 4804 2757
rect 4804 2731 4805 2757
rect 4777 2730 4805 2731
rect 3094 2534 3122 2562
rect 1768 2365 1796 2366
rect 1768 2339 1769 2365
rect 1769 2339 1795 2365
rect 1795 2339 1796 2365
rect 1768 2338 1796 2339
rect 1820 2365 1848 2366
rect 1820 2339 1821 2365
rect 1821 2339 1847 2365
rect 1847 2339 1848 2365
rect 1820 2338 1848 2339
rect 1872 2365 1900 2366
rect 1872 2339 1873 2365
rect 1873 2339 1899 2365
rect 1899 2339 1900 2365
rect 1872 2338 1900 2339
rect 2930 2365 2958 2366
rect 2930 2339 2931 2365
rect 2931 2339 2957 2365
rect 2957 2339 2958 2365
rect 2930 2338 2958 2339
rect 2982 2365 3010 2366
rect 2982 2339 2983 2365
rect 2983 2339 3009 2365
rect 3009 2339 3010 2365
rect 2982 2338 3010 2339
rect 3034 2365 3062 2366
rect 3034 2339 3035 2365
rect 3035 2339 3061 2365
rect 3061 2339 3062 2365
rect 3034 2338 3062 2339
rect 1187 1973 1215 1974
rect 1187 1947 1188 1973
rect 1188 1947 1214 1973
rect 1214 1947 1215 1973
rect 1187 1946 1215 1947
rect 1239 1973 1267 1974
rect 1239 1947 1240 1973
rect 1240 1947 1266 1973
rect 1266 1947 1267 1973
rect 1239 1946 1267 1947
rect 1291 1973 1319 1974
rect 1291 1947 1292 1973
rect 1292 1947 1318 1973
rect 1318 1947 1319 1973
rect 1291 1946 1319 1947
rect 2349 1973 2377 1974
rect 2349 1947 2350 1973
rect 2350 1947 2376 1973
rect 2376 1947 2377 1973
rect 2349 1946 2377 1947
rect 2401 1973 2429 1974
rect 2401 1947 2402 1973
rect 2402 1947 2428 1973
rect 2428 1947 2429 1973
rect 2401 1946 2429 1947
rect 2453 1973 2481 1974
rect 2453 1947 2454 1973
rect 2454 1947 2480 1973
rect 2480 1947 2481 1973
rect 2453 1946 2481 1947
rect 4092 2365 4120 2366
rect 4092 2339 4093 2365
rect 4093 2339 4119 2365
rect 4119 2339 4120 2365
rect 4092 2338 4120 2339
rect 4144 2365 4172 2366
rect 4144 2339 4145 2365
rect 4145 2339 4171 2365
rect 4171 2339 4172 2365
rect 4144 2338 4172 2339
rect 4196 2365 4224 2366
rect 4196 2339 4197 2365
rect 4197 2339 4223 2365
rect 4223 2339 4224 2365
rect 4196 2338 4224 2339
rect 5254 2365 5282 2366
rect 5254 2339 5255 2365
rect 5255 2339 5281 2365
rect 5281 2339 5282 2365
rect 5254 2338 5282 2339
rect 5306 2365 5334 2366
rect 5306 2339 5307 2365
rect 5307 2339 5333 2365
rect 5333 2339 5334 2365
rect 5306 2338 5334 2339
rect 5358 2365 5386 2366
rect 5358 2339 5359 2365
rect 5359 2339 5385 2365
rect 5385 2339 5386 2365
rect 5358 2338 5386 2339
rect 3511 1973 3539 1974
rect 3511 1947 3512 1973
rect 3512 1947 3538 1973
rect 3538 1947 3539 1973
rect 3511 1946 3539 1947
rect 3563 1973 3591 1974
rect 3563 1947 3564 1973
rect 3564 1947 3590 1973
rect 3590 1947 3591 1973
rect 3563 1946 3591 1947
rect 3615 1973 3643 1974
rect 3615 1947 3616 1973
rect 3616 1947 3642 1973
rect 3642 1947 3643 1973
rect 3615 1946 3643 1947
rect 4673 1973 4701 1974
rect 4673 1947 4674 1973
rect 4674 1947 4700 1973
rect 4700 1947 4701 1973
rect 4673 1946 4701 1947
rect 4725 1973 4753 1974
rect 4725 1947 4726 1973
rect 4726 1947 4752 1973
rect 4752 1947 4753 1973
rect 4725 1946 4753 1947
rect 4777 1973 4805 1974
rect 4777 1947 4778 1973
rect 4778 1947 4804 1973
rect 4804 1947 4805 1973
rect 4777 1946 4805 1947
rect 2870 1721 2898 1722
rect 2870 1695 2871 1721
rect 2871 1695 2897 1721
rect 2897 1695 2898 1721
rect 2870 1694 2898 1695
rect 1768 1581 1796 1582
rect 1768 1555 1769 1581
rect 1769 1555 1795 1581
rect 1795 1555 1796 1581
rect 1768 1554 1796 1555
rect 1820 1581 1848 1582
rect 1820 1555 1821 1581
rect 1821 1555 1847 1581
rect 1847 1555 1848 1581
rect 1820 1554 1848 1555
rect 1872 1581 1900 1582
rect 1872 1555 1873 1581
rect 1873 1555 1899 1581
rect 1899 1555 1900 1581
rect 1872 1554 1900 1555
rect 3598 1721 3626 1722
rect 3598 1695 3599 1721
rect 3599 1695 3625 1721
rect 3625 1695 3626 1721
rect 3598 1694 3626 1695
rect 2930 1581 2958 1582
rect 2930 1555 2931 1581
rect 2931 1555 2957 1581
rect 2957 1555 2958 1581
rect 2930 1554 2958 1555
rect 2982 1581 3010 1582
rect 2982 1555 2983 1581
rect 2983 1555 3009 1581
rect 3009 1555 3010 1581
rect 2982 1554 3010 1555
rect 3034 1581 3062 1582
rect 3034 1555 3035 1581
rect 3035 1555 3061 1581
rect 3061 1555 3062 1581
rect 3034 1554 3062 1555
rect 4092 1581 4120 1582
rect 4092 1555 4093 1581
rect 4093 1555 4119 1581
rect 4119 1555 4120 1581
rect 4092 1554 4120 1555
rect 4144 1581 4172 1582
rect 4144 1555 4145 1581
rect 4145 1555 4171 1581
rect 4171 1555 4172 1581
rect 4144 1554 4172 1555
rect 4196 1581 4224 1582
rect 4196 1555 4197 1581
rect 4197 1555 4223 1581
rect 4223 1555 4224 1581
rect 4196 1554 4224 1555
rect 5254 1581 5282 1582
rect 5254 1555 5255 1581
rect 5255 1555 5281 1581
rect 5281 1555 5282 1581
rect 5254 1554 5282 1555
rect 5306 1581 5334 1582
rect 5306 1555 5307 1581
rect 5307 1555 5333 1581
rect 5333 1555 5334 1581
rect 5306 1554 5334 1555
rect 5358 1581 5386 1582
rect 5358 1555 5359 1581
rect 5359 1555 5385 1581
rect 5385 1555 5386 1581
rect 5358 1554 5386 1555
<< metal3 >>
rect 1182 4298 1187 4326
rect 1215 4298 1239 4326
rect 1267 4298 1291 4326
rect 1319 4298 1324 4326
rect 2344 4298 2349 4326
rect 2377 4298 2401 4326
rect 2429 4298 2453 4326
rect 2481 4298 2486 4326
rect 3506 4298 3511 4326
rect 3539 4298 3563 4326
rect 3591 4298 3615 4326
rect 3643 4298 3648 4326
rect 4668 4298 4673 4326
rect 4701 4298 4725 4326
rect 4753 4298 4777 4326
rect 4805 4298 4810 4326
rect 2977 4158 2982 4186
rect 3010 4158 3430 4186
rect 3458 4158 3463 4186
rect 1763 3906 1768 3934
rect 1796 3906 1820 3934
rect 1848 3906 1872 3934
rect 1900 3906 1905 3934
rect 2925 3906 2930 3934
rect 2958 3906 2982 3934
rect 3010 3906 3034 3934
rect 3062 3906 3067 3934
rect 4087 3906 4092 3934
rect 4120 3906 4144 3934
rect 4172 3906 4196 3934
rect 4224 3906 4229 3934
rect 5249 3906 5254 3934
rect 5282 3906 5306 3934
rect 5334 3906 5358 3934
rect 5386 3906 5391 3934
rect 1182 3514 1187 3542
rect 1215 3514 1239 3542
rect 1267 3514 1291 3542
rect 1319 3514 1324 3542
rect 2344 3514 2349 3542
rect 2377 3514 2401 3542
rect 2429 3514 2453 3542
rect 2481 3514 2486 3542
rect 3506 3514 3511 3542
rect 3539 3514 3563 3542
rect 3591 3514 3615 3542
rect 3643 3514 3648 3542
rect 4668 3514 4673 3542
rect 4701 3514 4725 3542
rect 4753 3514 4777 3542
rect 4805 3514 4810 3542
rect 1763 3122 1768 3150
rect 1796 3122 1820 3150
rect 1848 3122 1872 3150
rect 1900 3122 1905 3150
rect 2925 3122 2930 3150
rect 2958 3122 2982 3150
rect 3010 3122 3034 3150
rect 3062 3122 3067 3150
rect 4087 3122 4092 3150
rect 4120 3122 4144 3150
rect 4172 3122 4196 3150
rect 4224 3122 4229 3150
rect 5249 3122 5254 3150
rect 5282 3122 5306 3150
rect 5334 3122 5358 3150
rect 5386 3122 5391 3150
rect 0 3010 400 3024
rect 0 2982 910 3010
rect 938 2982 943 3010
rect 0 2968 400 2982
rect 1182 2730 1187 2758
rect 1215 2730 1239 2758
rect 1267 2730 1291 2758
rect 1319 2730 1324 2758
rect 2344 2730 2349 2758
rect 2377 2730 2401 2758
rect 2429 2730 2453 2758
rect 2481 2730 2486 2758
rect 3506 2730 3511 2758
rect 3539 2730 3563 2758
rect 3591 2730 3615 2758
rect 3643 2730 3648 2758
rect 4668 2730 4673 2758
rect 4701 2730 4725 2758
rect 4753 2730 4777 2758
rect 4805 2730 4810 2758
rect 2361 2534 2366 2562
rect 2394 2534 3094 2562
rect 3122 2534 3127 2562
rect 1763 2338 1768 2366
rect 1796 2338 1820 2366
rect 1848 2338 1872 2366
rect 1900 2338 1905 2366
rect 2925 2338 2930 2366
rect 2958 2338 2982 2366
rect 3010 2338 3034 2366
rect 3062 2338 3067 2366
rect 4087 2338 4092 2366
rect 4120 2338 4144 2366
rect 4172 2338 4196 2366
rect 4224 2338 4229 2366
rect 5249 2338 5254 2366
rect 5282 2338 5306 2366
rect 5334 2338 5358 2366
rect 5386 2338 5391 2366
rect 1182 1946 1187 1974
rect 1215 1946 1239 1974
rect 1267 1946 1291 1974
rect 1319 1946 1324 1974
rect 2344 1946 2349 1974
rect 2377 1946 2401 1974
rect 2429 1946 2453 1974
rect 2481 1946 2486 1974
rect 3506 1946 3511 1974
rect 3539 1946 3563 1974
rect 3591 1946 3615 1974
rect 3643 1946 3648 1974
rect 4668 1946 4673 1974
rect 4701 1946 4725 1974
rect 4753 1946 4777 1974
rect 4805 1946 4810 1974
rect 2865 1694 2870 1722
rect 2898 1694 3598 1722
rect 3626 1694 3631 1722
rect 1763 1554 1768 1582
rect 1796 1554 1820 1582
rect 1848 1554 1872 1582
rect 1900 1554 1905 1582
rect 2925 1554 2930 1582
rect 2958 1554 2982 1582
rect 3010 1554 3034 1582
rect 3062 1554 3067 1582
rect 4087 1554 4092 1582
rect 4120 1554 4144 1582
rect 4172 1554 4196 1582
rect 4224 1554 4229 1582
rect 5249 1554 5254 1582
rect 5282 1554 5306 1582
rect 5334 1554 5358 1582
rect 5386 1554 5391 1582
<< via3 >>
rect 1187 4298 1215 4326
rect 1239 4298 1267 4326
rect 1291 4298 1319 4326
rect 2349 4298 2377 4326
rect 2401 4298 2429 4326
rect 2453 4298 2481 4326
rect 3511 4298 3539 4326
rect 3563 4298 3591 4326
rect 3615 4298 3643 4326
rect 4673 4298 4701 4326
rect 4725 4298 4753 4326
rect 4777 4298 4805 4326
rect 1768 3906 1796 3934
rect 1820 3906 1848 3934
rect 1872 3906 1900 3934
rect 2930 3906 2958 3934
rect 2982 3906 3010 3934
rect 3034 3906 3062 3934
rect 4092 3906 4120 3934
rect 4144 3906 4172 3934
rect 4196 3906 4224 3934
rect 5254 3906 5282 3934
rect 5306 3906 5334 3934
rect 5358 3906 5386 3934
rect 1187 3514 1215 3542
rect 1239 3514 1267 3542
rect 1291 3514 1319 3542
rect 2349 3514 2377 3542
rect 2401 3514 2429 3542
rect 2453 3514 2481 3542
rect 3511 3514 3539 3542
rect 3563 3514 3591 3542
rect 3615 3514 3643 3542
rect 4673 3514 4701 3542
rect 4725 3514 4753 3542
rect 4777 3514 4805 3542
rect 1768 3122 1796 3150
rect 1820 3122 1848 3150
rect 1872 3122 1900 3150
rect 2930 3122 2958 3150
rect 2982 3122 3010 3150
rect 3034 3122 3062 3150
rect 4092 3122 4120 3150
rect 4144 3122 4172 3150
rect 4196 3122 4224 3150
rect 5254 3122 5282 3150
rect 5306 3122 5334 3150
rect 5358 3122 5386 3150
rect 1187 2730 1215 2758
rect 1239 2730 1267 2758
rect 1291 2730 1319 2758
rect 2349 2730 2377 2758
rect 2401 2730 2429 2758
rect 2453 2730 2481 2758
rect 3511 2730 3539 2758
rect 3563 2730 3591 2758
rect 3615 2730 3643 2758
rect 4673 2730 4701 2758
rect 4725 2730 4753 2758
rect 4777 2730 4805 2758
rect 1768 2338 1796 2366
rect 1820 2338 1848 2366
rect 1872 2338 1900 2366
rect 2930 2338 2958 2366
rect 2982 2338 3010 2366
rect 3034 2338 3062 2366
rect 4092 2338 4120 2366
rect 4144 2338 4172 2366
rect 4196 2338 4224 2366
rect 5254 2338 5282 2366
rect 5306 2338 5334 2366
rect 5358 2338 5386 2366
rect 1187 1946 1215 1974
rect 1239 1946 1267 1974
rect 1291 1946 1319 1974
rect 2349 1946 2377 1974
rect 2401 1946 2429 1974
rect 2453 1946 2481 1974
rect 3511 1946 3539 1974
rect 3563 1946 3591 1974
rect 3615 1946 3643 1974
rect 4673 1946 4701 1974
rect 4725 1946 4753 1974
rect 4777 1946 4805 1974
rect 1768 1554 1796 1582
rect 1820 1554 1848 1582
rect 1872 1554 1900 1582
rect 2930 1554 2958 1582
rect 2982 1554 3010 1582
rect 3034 1554 3062 1582
rect 4092 1554 4120 1582
rect 4144 1554 4172 1582
rect 4196 1554 4224 1582
rect 5254 1554 5282 1582
rect 5306 1554 5334 1582
rect 5358 1554 5386 1582
<< metal4 >>
rect 1173 4326 1333 4342
rect 1173 4298 1187 4326
rect 1215 4298 1239 4326
rect 1267 4298 1291 4326
rect 1319 4298 1333 4326
rect 1173 3542 1333 4298
rect 1173 3514 1187 3542
rect 1215 3514 1239 3542
rect 1267 3514 1291 3542
rect 1319 3514 1333 3542
rect 1173 2758 1333 3514
rect 1173 2730 1187 2758
rect 1215 2730 1239 2758
rect 1267 2730 1291 2758
rect 1319 2730 1333 2758
rect 1173 1974 1333 2730
rect 1173 1946 1187 1974
rect 1215 1946 1239 1974
rect 1267 1946 1291 1974
rect 1319 1946 1333 1974
rect 1173 1538 1333 1946
rect 1754 3934 1914 4342
rect 1754 3906 1768 3934
rect 1796 3906 1820 3934
rect 1848 3906 1872 3934
rect 1900 3906 1914 3934
rect 1754 3150 1914 3906
rect 1754 3122 1768 3150
rect 1796 3122 1820 3150
rect 1848 3122 1872 3150
rect 1900 3122 1914 3150
rect 1754 2366 1914 3122
rect 1754 2338 1768 2366
rect 1796 2338 1820 2366
rect 1848 2338 1872 2366
rect 1900 2338 1914 2366
rect 1754 1582 1914 2338
rect 1754 1554 1768 1582
rect 1796 1554 1820 1582
rect 1848 1554 1872 1582
rect 1900 1554 1914 1582
rect 1754 1538 1914 1554
rect 2335 4326 2495 4342
rect 2335 4298 2349 4326
rect 2377 4298 2401 4326
rect 2429 4298 2453 4326
rect 2481 4298 2495 4326
rect 2335 3542 2495 4298
rect 2335 3514 2349 3542
rect 2377 3514 2401 3542
rect 2429 3514 2453 3542
rect 2481 3514 2495 3542
rect 2335 2758 2495 3514
rect 2335 2730 2349 2758
rect 2377 2730 2401 2758
rect 2429 2730 2453 2758
rect 2481 2730 2495 2758
rect 2335 1974 2495 2730
rect 2335 1946 2349 1974
rect 2377 1946 2401 1974
rect 2429 1946 2453 1974
rect 2481 1946 2495 1974
rect 2335 1538 2495 1946
rect 2916 3934 3076 4342
rect 2916 3906 2930 3934
rect 2958 3906 2982 3934
rect 3010 3906 3034 3934
rect 3062 3906 3076 3934
rect 2916 3150 3076 3906
rect 2916 3122 2930 3150
rect 2958 3122 2982 3150
rect 3010 3122 3034 3150
rect 3062 3122 3076 3150
rect 2916 2366 3076 3122
rect 2916 2338 2930 2366
rect 2958 2338 2982 2366
rect 3010 2338 3034 2366
rect 3062 2338 3076 2366
rect 2916 1582 3076 2338
rect 2916 1554 2930 1582
rect 2958 1554 2982 1582
rect 3010 1554 3034 1582
rect 3062 1554 3076 1582
rect 2916 1538 3076 1554
rect 3497 4326 3657 4342
rect 3497 4298 3511 4326
rect 3539 4298 3563 4326
rect 3591 4298 3615 4326
rect 3643 4298 3657 4326
rect 3497 3542 3657 4298
rect 3497 3514 3511 3542
rect 3539 3514 3563 3542
rect 3591 3514 3615 3542
rect 3643 3514 3657 3542
rect 3497 2758 3657 3514
rect 3497 2730 3511 2758
rect 3539 2730 3563 2758
rect 3591 2730 3615 2758
rect 3643 2730 3657 2758
rect 3497 1974 3657 2730
rect 3497 1946 3511 1974
rect 3539 1946 3563 1974
rect 3591 1946 3615 1974
rect 3643 1946 3657 1974
rect 3497 1538 3657 1946
rect 4078 3934 4238 4342
rect 4078 3906 4092 3934
rect 4120 3906 4144 3934
rect 4172 3906 4196 3934
rect 4224 3906 4238 3934
rect 4078 3150 4238 3906
rect 4078 3122 4092 3150
rect 4120 3122 4144 3150
rect 4172 3122 4196 3150
rect 4224 3122 4238 3150
rect 4078 2366 4238 3122
rect 4078 2338 4092 2366
rect 4120 2338 4144 2366
rect 4172 2338 4196 2366
rect 4224 2338 4238 2366
rect 4078 1582 4238 2338
rect 4078 1554 4092 1582
rect 4120 1554 4144 1582
rect 4172 1554 4196 1582
rect 4224 1554 4238 1582
rect 4078 1538 4238 1554
rect 4659 4326 4819 4342
rect 4659 4298 4673 4326
rect 4701 4298 4725 4326
rect 4753 4298 4777 4326
rect 4805 4298 4819 4326
rect 4659 3542 4819 4298
rect 4659 3514 4673 3542
rect 4701 3514 4725 3542
rect 4753 3514 4777 3542
rect 4805 3514 4819 3542
rect 4659 2758 4819 3514
rect 4659 2730 4673 2758
rect 4701 2730 4725 2758
rect 4753 2730 4777 2758
rect 4805 2730 4819 2758
rect 4659 1974 4819 2730
rect 4659 1946 4673 1974
rect 4701 1946 4725 1974
rect 4753 1946 4777 1974
rect 4805 1946 4819 1974
rect 4659 1538 4819 1946
rect 5240 3934 5400 4342
rect 5240 3906 5254 3934
rect 5282 3906 5306 3934
rect 5334 3906 5358 3934
rect 5386 3906 5400 3934
rect 5240 3150 5400 3906
rect 5240 3122 5254 3150
rect 5282 3122 5306 3150
rect 5334 3122 5358 3150
rect 5386 3122 5400 3150
rect 5240 2366 5400 3122
rect 5240 2338 5254 2366
rect 5282 2338 5306 2366
rect 5334 2338 5358 2366
rect 5386 2338 5400 2366
rect 5240 1582 5400 2338
rect 5240 1554 5254 1582
rect 5282 1554 5306 1582
rect 5334 1554 5358 1582
rect 5386 1554 5400 1582
rect 5240 1538 5400 1554
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 2912 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1669390400
transform -1 0 952 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2 Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 784 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34 Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 2576 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37
timestamp 1669390400
transform 1 0 2744 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40 Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 2912 0 1 1568
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58 Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 3920 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66 Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 4368 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_72
timestamp 1669390400
transform 1 0 4704 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80
timestamp 1669390400
transform 1 0 5152 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_2 Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 784 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_66
timestamp 1669390400
transform 1 0 4368 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_70
timestamp 1669390400
transform 1 0 4592 0 -1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_73
timestamp 1669390400
transform 1 0 4760 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_2 Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 784 0 1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_18
timestamp 1669390400
transform 1 0 1680 0 1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_26
timestamp 1669390400
transform 1 0 2128 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_32
timestamp 1669390400
transform 1 0 2464 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_34
timestamp 1669390400
transform 1 0 2576 0 1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_37
timestamp 1669390400
transform 1 0 2744 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_69
timestamp 1669390400
transform 1 0 4536 0 1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_77
timestamp 1669390400
transform 1 0 4984 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_2
timestamp 1669390400
transform 1 0 784 0 -1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_5
timestamp 1669390400
transform 1 0 952 0 -1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_13
timestamp 1669390400
transform 1 0 1400 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_17
timestamp 1669390400
transform 1 0 1624 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_39
timestamp 1669390400
transform 1 0 2856 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_49
timestamp 1669390400
transform 1 0 3416 0 -1 3136
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_65
timestamp 1669390400
transform 1 0 4312 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_69
timestamp 1669390400
transform 1 0 4536 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_73
timestamp 1669390400
transform 1 0 4760 0 -1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_2
timestamp 1669390400
transform 1 0 784 0 1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_19
timestamp 1669390400
transform 1 0 1736 0 1 3136
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_37
timestamp 1669390400
transform 1 0 2744 0 1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_44
timestamp 1669390400
transform 1 0 3136 0 1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_76
timestamp 1669390400
transform 1 0 4928 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_80
timestamp 1669390400
transform 1 0 5152 0 1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_2
timestamp 1669390400
transform 1 0 784 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_66
timestamp 1669390400
transform 1 0 4368 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_70
timestamp 1669390400
transform 1 0 4592 0 -1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_73
timestamp 1669390400
transform 1 0 4760 0 -1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_2
timestamp 1669390400
transform 1 0 784 0 1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_34
timestamp 1669390400
transform 1 0 2576 0 1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_37
timestamp 1669390400
transform 1 0 2744 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_41
timestamp 1669390400
transform 1 0 2968 0 1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_56
timestamp 1669390400
transform 1 0 3808 0 1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_64
timestamp 1669390400
transform 1 0 4256 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_68
timestamp 1669390400
transform 1 0 4480 0 1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_72
timestamp 1669390400
transform 1 0 4704 0 1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_80
timestamp 1669390400
transform 1 0 5152 0 1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_0 Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 672 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_1
timestamp 1669390400
transform -1 0 5320 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_2
timestamp 1669390400
transform 1 0 672 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_3
timestamp 1669390400
transform -1 0 5320 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_4
timestamp 1669390400
transform 1 0 672 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_5
timestamp 1669390400
transform -1 0 5320 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_6
timestamp 1669390400
transform 1 0 672 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_7
timestamp 1669390400
transform -1 0 5320 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_8
timestamp 1669390400
transform 1 0 672 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_9
timestamp 1669390400
transform -1 0 5320 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_10
timestamp 1669390400
transform 1 0 672 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_11
timestamp 1669390400
transform -1 0 5320 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_12
timestamp 1669390400
transform 1 0 672 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_13
timestamp 1669390400
transform -1 0 5320 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_14 Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 2632 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_15
timestamp 1669390400
transform 1 0 4592 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_16
timestamp 1669390400
transform 1 0 4648 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_17
timestamp 1669390400
transform 1 0 2632 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_18
timestamp 1669390400
transform 1 0 4648 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_19
timestamp 1669390400
transform 1 0 2632 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_20
timestamp 1669390400
transform 1 0 4648 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_21
timestamp 1669390400
transform 1 0 2632 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_22
timestamp 1669390400
transform 1 0 4592 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 2464 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _3_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 2968 0 -1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _4_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 2800 0 1 3136
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _5_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 1736 0 -1 3136
box -43 -43 1163 435
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input1 Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 3920 0 1 1568
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input2
timestamp 1669390400
transform 1 0 840 0 1 3136
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output3 Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 3024 0 1 3920
box -43 -43 827 435
<< labels >>
flabel metal2 s 2968 0 3024 400 0 FreeSans 224 90 0 0 clk
port 0 nsew signal input
flabel metal3 s 0 2968 400 3024 0 FreeSans 224 0 0 0 gate
port 1 nsew signal input
flabel metal2 s 2968 5600 3024 6000 0 FreeSans 224 90 0 0 gclk
port 2 nsew signal tristate
flabel metal4 s 1173 1538 1333 4342 0 FreeSans 640 90 0 0 vdd
port 3 nsew power bidirectional
flabel metal4 s 2335 1538 2495 4342 0 FreeSans 640 90 0 0 vdd
port 3 nsew power bidirectional
flabel metal4 s 3497 1538 3657 4342 0 FreeSans 640 90 0 0 vdd
port 3 nsew power bidirectional
flabel metal4 s 4659 1538 4819 4342 0 FreeSans 640 90 0 0 vdd
port 3 nsew power bidirectional
flabel metal4 s 1754 1538 1914 4342 0 FreeSans 640 90 0 0 vss
port 4 nsew ground bidirectional
flabel metal4 s 2916 1538 3076 4342 0 FreeSans 640 90 0 0 vss
port 4 nsew ground bidirectional
flabel metal4 s 4078 1538 4238 4342 0 FreeSans 640 90 0 0 vss
port 4 nsew ground bidirectional
flabel metal4 s 5240 1538 5400 4342 0 FreeSans 640 90 0 0 vss
port 4 nsew ground bidirectional
rlabel metal1 2996 4312 2996 4312 0 vdd
rlabel via1 3036 3920 3036 3920 0 vss
rlabel metal2 3108 3052 3108 3052 0 _0_
rlabel metal2 2296 2660 2296 2660 0 _1_
rlabel metal2 2884 1428 2884 1428 0 clk
rlabel metal2 3164 2968 3164 2968 0 clkp
rlabel metal3 651 2996 651 2996 0 gate
rlabel metal3 3220 4172 3220 4172 0 gclk
rlabel metal2 3080 2884 3080 2884 0 net1
rlabel metal2 2100 3108 2100 3108 0 net2
rlabel metal2 3080 3276 3080 3276 0 net3
<< properties >>
string FIXED_BBOX 0 0 6000 6000
<< end >>
