magic
tech gf180mcuC
magscale 1 5
timestamp 1670260635
<< metal1 >>
rect 672 3149 4392 3166
rect 672 3123 1517 3149
rect 1543 3123 1569 3149
rect 1595 3123 1621 3149
rect 1647 3123 2427 3149
rect 2453 3123 2479 3149
rect 2505 3123 2531 3149
rect 2557 3123 3337 3149
rect 3363 3123 3389 3149
rect 3415 3123 3441 3149
rect 3467 3123 4247 3149
rect 4273 3123 4299 3149
rect 4325 3123 4351 3149
rect 4377 3123 4392 3149
rect 672 3106 4392 3123
rect 2255 3009 2281 3015
rect 1409 2983 1415 3009
rect 1441 2983 1447 3009
rect 3425 2983 3431 3009
rect 3457 2983 3463 3009
rect 2255 2977 2281 2983
rect 1969 2927 1975 2953
rect 2001 2927 2007 2953
rect 2361 2927 2367 2953
rect 2393 2927 2399 2953
rect 2473 2927 2479 2953
rect 2505 2927 2511 2953
rect 2865 2927 2871 2953
rect 2897 2927 2903 2953
rect 1023 2897 1049 2903
rect 1023 2865 1049 2871
rect 1079 2897 1105 2903
rect 1079 2865 1105 2871
rect 2199 2841 2225 2847
rect 2199 2809 2225 2815
rect 672 2757 4312 2774
rect 672 2731 1062 2757
rect 1088 2731 1114 2757
rect 1140 2731 1166 2757
rect 1192 2731 1972 2757
rect 1998 2731 2024 2757
rect 2050 2731 2076 2757
rect 2102 2731 2882 2757
rect 2908 2731 2934 2757
rect 2960 2731 2986 2757
rect 3012 2731 3792 2757
rect 3818 2731 3844 2757
rect 3870 2731 3896 2757
rect 3922 2731 4312 2757
rect 672 2714 4312 2731
rect 2423 2617 2449 2623
rect 961 2591 967 2617
rect 993 2591 999 2617
rect 2423 2585 2449 2591
rect 1807 2561 1833 2567
rect 1521 2535 1527 2561
rect 1553 2535 1559 2561
rect 1807 2529 1833 2535
rect 1863 2561 1889 2567
rect 1863 2529 1889 2535
rect 1975 2561 2001 2567
rect 2081 2535 2087 2561
rect 2113 2535 2119 2561
rect 1975 2529 2001 2535
rect 2367 2449 2393 2455
rect 2367 2417 2393 2423
rect 672 2365 4392 2382
rect 672 2339 1517 2365
rect 1543 2339 1569 2365
rect 1595 2339 1621 2365
rect 1647 2339 2427 2365
rect 2453 2339 2479 2365
rect 2505 2339 2531 2365
rect 2557 2339 3337 2365
rect 3363 2339 3389 2365
rect 3415 2339 3441 2365
rect 3467 2339 4247 2365
rect 4273 2339 4299 2365
rect 4325 2339 4351 2365
rect 4377 2339 4392 2365
rect 672 2322 4392 2339
rect 2423 2225 2449 2231
rect 3481 2199 3487 2225
rect 3513 2199 3519 2225
rect 2423 2193 2449 2199
rect 1975 2169 2001 2175
rect 1409 2143 1415 2169
rect 1441 2143 1447 2169
rect 1975 2137 2001 2143
rect 2143 2169 2169 2175
rect 2143 2137 2169 2143
rect 3935 2169 3961 2175
rect 3935 2137 3961 2143
rect 2031 2113 2057 2119
rect 961 2087 967 2113
rect 993 2087 999 2113
rect 2031 2081 2057 2087
rect 2199 2113 2225 2119
rect 2199 2081 2225 2087
rect 672 1973 4312 1990
rect 672 1947 1062 1973
rect 1088 1947 1114 1973
rect 1140 1947 1166 1973
rect 1192 1947 1972 1973
rect 1998 1947 2024 1973
rect 2050 1947 2076 1973
rect 2102 1947 2882 1973
rect 2908 1947 2934 1973
rect 2960 1947 2986 1973
rect 3012 1947 3792 1973
rect 3818 1947 3844 1973
rect 3870 1947 3896 1973
rect 3922 1947 4312 1973
rect 672 1930 4312 1947
rect 2255 1889 2281 1895
rect 2255 1857 2281 1863
rect 1689 1807 1695 1833
rect 1721 1807 1727 1833
rect 2865 1807 2871 1833
rect 2897 1807 2903 1833
rect 1919 1777 1945 1783
rect 2081 1751 2087 1777
rect 2113 1751 2119 1777
rect 1919 1745 1945 1751
rect 2199 1721 2225 1727
rect 1017 1695 1023 1721
rect 1049 1695 1055 1721
rect 2199 1689 2225 1695
rect 2423 1721 2449 1727
rect 3879 1721 3905 1727
rect 3537 1695 3543 1721
rect 3569 1695 3575 1721
rect 2423 1689 2449 1695
rect 3879 1689 3905 1695
rect 672 1581 4392 1598
rect 672 1555 1517 1581
rect 1543 1555 1569 1581
rect 1595 1555 1621 1581
rect 1647 1555 2427 1581
rect 2453 1555 2479 1581
rect 2505 1555 2531 1581
rect 2557 1555 3337 1581
rect 3363 1555 3389 1581
rect 3415 1555 3441 1581
rect 3467 1555 4247 1581
rect 4273 1555 4299 1581
rect 4325 1555 4351 1581
rect 4377 1555 4392 1581
rect 672 1538 4392 1555
<< via1 >>
rect 1517 3123 1543 3149
rect 1569 3123 1595 3149
rect 1621 3123 1647 3149
rect 2427 3123 2453 3149
rect 2479 3123 2505 3149
rect 2531 3123 2557 3149
rect 3337 3123 3363 3149
rect 3389 3123 3415 3149
rect 3441 3123 3467 3149
rect 4247 3123 4273 3149
rect 4299 3123 4325 3149
rect 4351 3123 4377 3149
rect 1415 2983 1441 3009
rect 2255 2983 2281 3009
rect 3431 2983 3457 3009
rect 1975 2927 2001 2953
rect 2367 2927 2393 2953
rect 2479 2927 2505 2953
rect 2871 2927 2897 2953
rect 1023 2871 1049 2897
rect 1079 2871 1105 2897
rect 2199 2815 2225 2841
rect 1062 2731 1088 2757
rect 1114 2731 1140 2757
rect 1166 2731 1192 2757
rect 1972 2731 1998 2757
rect 2024 2731 2050 2757
rect 2076 2731 2102 2757
rect 2882 2731 2908 2757
rect 2934 2731 2960 2757
rect 2986 2731 3012 2757
rect 3792 2731 3818 2757
rect 3844 2731 3870 2757
rect 3896 2731 3922 2757
rect 967 2591 993 2617
rect 2423 2591 2449 2617
rect 1527 2535 1553 2561
rect 1807 2535 1833 2561
rect 1863 2535 1889 2561
rect 1975 2535 2001 2561
rect 2087 2535 2113 2561
rect 2367 2423 2393 2449
rect 1517 2339 1543 2365
rect 1569 2339 1595 2365
rect 1621 2339 1647 2365
rect 2427 2339 2453 2365
rect 2479 2339 2505 2365
rect 2531 2339 2557 2365
rect 3337 2339 3363 2365
rect 3389 2339 3415 2365
rect 3441 2339 3467 2365
rect 4247 2339 4273 2365
rect 4299 2339 4325 2365
rect 4351 2339 4377 2365
rect 2423 2199 2449 2225
rect 3487 2199 3513 2225
rect 1415 2143 1441 2169
rect 1975 2143 2001 2169
rect 2143 2143 2169 2169
rect 3935 2143 3961 2169
rect 967 2087 993 2113
rect 2031 2087 2057 2113
rect 2199 2087 2225 2113
rect 1062 1947 1088 1973
rect 1114 1947 1140 1973
rect 1166 1947 1192 1973
rect 1972 1947 1998 1973
rect 2024 1947 2050 1973
rect 2076 1947 2102 1973
rect 2882 1947 2908 1973
rect 2934 1947 2960 1973
rect 2986 1947 3012 1973
rect 3792 1947 3818 1973
rect 3844 1947 3870 1973
rect 3896 1947 3922 1973
rect 2255 1863 2281 1889
rect 1695 1807 1721 1833
rect 2871 1807 2897 1833
rect 1919 1751 1945 1777
rect 2087 1751 2113 1777
rect 1023 1695 1049 1721
rect 2199 1695 2225 1721
rect 2423 1695 2449 1721
rect 3543 1695 3569 1721
rect 3879 1695 3905 1721
rect 1517 1555 1543 1581
rect 1569 1555 1595 1581
rect 1621 1555 1647 1581
rect 2427 1555 2453 1581
rect 2479 1555 2505 1581
rect 2531 1555 2557 1581
rect 3337 1555 3363 1581
rect 3389 1555 3415 1581
rect 3441 1555 3467 1581
rect 4247 1555 4273 1581
rect 4299 1555 4325 1581
rect 4351 1555 4377 1581
<< metal2 >>
rect 1232 4600 1288 5000
rect 3696 4600 3752 5000
rect 966 3738 994 3743
rect 966 2617 994 3710
rect 1246 3010 1274 4600
rect 1516 3150 1648 3155
rect 1544 3122 1568 3150
rect 1596 3122 1620 3150
rect 1516 3117 1648 3122
rect 2426 3150 2558 3155
rect 2454 3122 2478 3150
rect 2506 3122 2530 3150
rect 2426 3117 2558 3122
rect 3336 3150 3468 3155
rect 3364 3122 3388 3150
rect 3416 3122 3440 3150
rect 3336 3117 3468 3122
rect 1414 3010 1442 3015
rect 1246 3009 1442 3010
rect 1246 2983 1415 3009
rect 1441 2983 1442 3009
rect 1246 2982 1442 2983
rect 1414 2977 1442 2982
rect 2254 3010 2282 3015
rect 3430 3010 3458 3015
rect 2254 3009 2338 3010
rect 2254 2983 2255 3009
rect 2281 2983 2338 3009
rect 2254 2982 2338 2983
rect 2254 2977 2282 2982
rect 1974 2954 2002 2959
rect 1974 2953 2170 2954
rect 1974 2927 1975 2953
rect 2001 2927 2170 2953
rect 1974 2926 2170 2927
rect 1974 2921 2002 2926
rect 1022 2897 1050 2903
rect 1022 2871 1023 2897
rect 1049 2871 1050 2897
rect 1022 2842 1050 2871
rect 1078 2898 1106 2903
rect 1078 2851 1106 2870
rect 1750 2898 1778 2903
rect 1022 2809 1050 2814
rect 1414 2842 1442 2847
rect 1061 2758 1193 2763
rect 1089 2730 1113 2758
rect 1141 2730 1165 2758
rect 1061 2725 1193 2730
rect 966 2591 967 2617
rect 993 2591 994 2617
rect 966 2585 994 2591
rect 1414 2169 1442 2814
rect 1694 2618 1722 2623
rect 1526 2562 1554 2567
rect 1526 2515 1554 2534
rect 1516 2366 1648 2371
rect 1544 2338 1568 2366
rect 1596 2338 1620 2366
rect 1516 2333 1648 2338
rect 1414 2143 1415 2169
rect 1441 2143 1442 2169
rect 1414 2137 1442 2143
rect 966 2113 994 2119
rect 966 2087 967 2113
rect 993 2087 994 2113
rect 966 1274 994 2087
rect 1061 1974 1193 1979
rect 1089 1946 1113 1974
rect 1141 1946 1165 1974
rect 1061 1941 1193 1946
rect 1694 1833 1722 2590
rect 1750 2114 1778 2870
rect 1971 2758 2103 2763
rect 1999 2730 2023 2758
rect 2051 2730 2075 2758
rect 1971 2725 2103 2730
rect 1806 2562 1834 2567
rect 1806 2515 1834 2534
rect 1862 2561 1890 2567
rect 1862 2535 1863 2561
rect 1889 2535 1890 2561
rect 1862 2282 1890 2535
rect 1974 2562 2002 2567
rect 1974 2515 2002 2534
rect 2086 2562 2114 2567
rect 1862 2249 1890 2254
rect 2086 2226 2114 2534
rect 2142 2394 2170 2926
rect 2198 2842 2226 2847
rect 2198 2795 2226 2814
rect 2310 2786 2338 2982
rect 3430 2963 3458 2982
rect 3710 3010 3738 4600
rect 4246 3150 4378 3155
rect 4274 3122 4298 3150
rect 4326 3122 4350 3150
rect 4246 3117 4378 3122
rect 3710 2977 3738 2982
rect 2366 2953 2394 2959
rect 2366 2927 2367 2953
rect 2393 2927 2394 2953
rect 2366 2898 2394 2927
rect 2366 2865 2394 2870
rect 2478 2953 2506 2959
rect 2870 2954 2898 2959
rect 2478 2927 2479 2953
rect 2505 2927 2506 2953
rect 2310 2758 2450 2786
rect 2422 2617 2450 2758
rect 2422 2591 2423 2617
rect 2449 2591 2450 2617
rect 2310 2506 2338 2511
rect 2142 2366 2282 2394
rect 1974 2198 2086 2226
rect 1974 2170 2002 2198
rect 1750 2081 1778 2086
rect 1862 2169 2002 2170
rect 1862 2143 1975 2169
rect 2001 2143 2002 2169
rect 2086 2160 2114 2198
rect 2142 2282 2170 2287
rect 2142 2169 2170 2254
rect 1862 2142 2002 2143
rect 1694 1807 1695 1833
rect 1721 1807 1722 1833
rect 1694 1801 1722 1807
rect 1862 1778 1890 2142
rect 1974 2137 2002 2142
rect 2142 2143 2143 2169
rect 2169 2143 2170 2169
rect 2142 2137 2170 2143
rect 2030 2114 2058 2119
rect 2030 2058 2058 2086
rect 2198 2114 2226 2119
rect 2198 2067 2226 2086
rect 2030 2030 2170 2058
rect 1971 1974 2103 1979
rect 1999 1946 2023 1974
rect 2051 1946 2075 1974
rect 1971 1941 2103 1946
rect 1918 1778 1946 1783
rect 1862 1777 1946 1778
rect 1862 1751 1919 1777
rect 1945 1751 1946 1777
rect 1862 1750 1946 1751
rect 1918 1745 1946 1750
rect 2086 1778 2114 1783
rect 2142 1778 2170 2030
rect 2254 1889 2282 2366
rect 2254 1863 2255 1889
rect 2281 1863 2282 1889
rect 2254 1857 2282 1863
rect 2086 1777 2170 1778
rect 2086 1751 2087 1777
rect 2113 1751 2170 1777
rect 2086 1750 2170 1751
rect 2310 1834 2338 2478
rect 2422 2506 2450 2591
rect 2478 2562 2506 2927
rect 2478 2529 2506 2534
rect 2814 2953 2898 2954
rect 2814 2927 2871 2953
rect 2897 2927 2898 2953
rect 2814 2926 2898 2927
rect 2422 2473 2450 2478
rect 2366 2449 2394 2455
rect 2366 2423 2367 2449
rect 2393 2423 2394 2449
rect 2366 2282 2394 2423
rect 2426 2366 2558 2371
rect 2454 2338 2478 2366
rect 2506 2338 2530 2366
rect 2426 2333 2558 2338
rect 2366 2249 2394 2254
rect 2422 2226 2450 2231
rect 2422 2179 2450 2198
rect 2086 1745 2114 1750
rect 966 1241 994 1246
rect 1022 1722 1050 1727
rect 1022 1106 1050 1694
rect 2198 1722 2226 1727
rect 2310 1722 2338 1806
rect 2198 1721 2338 1722
rect 2198 1695 2199 1721
rect 2225 1695 2338 1721
rect 2198 1694 2338 1695
rect 2366 2170 2394 2175
rect 2198 1689 2226 1694
rect 1516 1582 1648 1587
rect 1544 1554 1568 1582
rect 1596 1554 1620 1582
rect 1516 1549 1648 1554
rect 2366 1442 2394 2142
rect 2814 2114 2842 2926
rect 2870 2921 2898 2926
rect 2881 2758 3013 2763
rect 2909 2730 2933 2758
rect 2961 2730 2985 2758
rect 2881 2725 3013 2730
rect 3791 2758 3923 2763
rect 3819 2730 3843 2758
rect 3871 2730 3895 2758
rect 3791 2725 3923 2730
rect 3336 2366 3468 2371
rect 3364 2338 3388 2366
rect 3416 2338 3440 2366
rect 3336 2333 3468 2338
rect 4246 2366 4378 2371
rect 4274 2338 4298 2366
rect 4326 2338 4350 2366
rect 4246 2333 4378 2338
rect 3486 2225 3514 2231
rect 3486 2199 3487 2225
rect 3513 2199 3514 2225
rect 3486 2170 3514 2199
rect 3486 2137 3514 2142
rect 3934 2170 3962 2175
rect 3934 2123 3962 2142
rect 2814 2081 2842 2086
rect 2881 1974 3013 1979
rect 2909 1946 2933 1974
rect 2961 1946 2985 1974
rect 2881 1941 3013 1946
rect 3791 1974 3923 1979
rect 3819 1946 3843 1974
rect 3871 1946 3895 1974
rect 3791 1941 3923 1946
rect 2870 1834 2898 1839
rect 2870 1787 2898 1806
rect 2422 1722 2450 1727
rect 2422 1675 2450 1694
rect 3542 1722 3570 1727
rect 3542 1675 3570 1694
rect 3878 1722 3906 1727
rect 2426 1582 2558 1587
rect 2454 1554 2478 1582
rect 2506 1554 2530 1582
rect 2426 1549 2558 1554
rect 3336 1582 3468 1587
rect 3364 1554 3388 1582
rect 3416 1554 3440 1582
rect 3336 1549 3468 1554
rect 2366 1414 2506 1442
rect 854 1078 1050 1106
rect 854 400 882 1078
rect 2478 400 2506 1414
rect 3878 1106 3906 1694
rect 4246 1582 4378 1587
rect 4274 1554 4298 1582
rect 4326 1554 4350 1582
rect 4246 1549 4378 1554
rect 3878 1078 4130 1106
rect 4102 400 4130 1078
rect 840 0 896 400
rect 2464 0 2520 400
rect 4088 0 4144 400
<< via2 >>
rect 966 3710 994 3738
rect 1516 3149 1544 3150
rect 1516 3123 1517 3149
rect 1517 3123 1543 3149
rect 1543 3123 1544 3149
rect 1516 3122 1544 3123
rect 1568 3149 1596 3150
rect 1568 3123 1569 3149
rect 1569 3123 1595 3149
rect 1595 3123 1596 3149
rect 1568 3122 1596 3123
rect 1620 3149 1648 3150
rect 1620 3123 1621 3149
rect 1621 3123 1647 3149
rect 1647 3123 1648 3149
rect 1620 3122 1648 3123
rect 2426 3149 2454 3150
rect 2426 3123 2427 3149
rect 2427 3123 2453 3149
rect 2453 3123 2454 3149
rect 2426 3122 2454 3123
rect 2478 3149 2506 3150
rect 2478 3123 2479 3149
rect 2479 3123 2505 3149
rect 2505 3123 2506 3149
rect 2478 3122 2506 3123
rect 2530 3149 2558 3150
rect 2530 3123 2531 3149
rect 2531 3123 2557 3149
rect 2557 3123 2558 3149
rect 2530 3122 2558 3123
rect 3336 3149 3364 3150
rect 3336 3123 3337 3149
rect 3337 3123 3363 3149
rect 3363 3123 3364 3149
rect 3336 3122 3364 3123
rect 3388 3149 3416 3150
rect 3388 3123 3389 3149
rect 3389 3123 3415 3149
rect 3415 3123 3416 3149
rect 3388 3122 3416 3123
rect 3440 3149 3468 3150
rect 3440 3123 3441 3149
rect 3441 3123 3467 3149
rect 3467 3123 3468 3149
rect 3440 3122 3468 3123
rect 1078 2897 1106 2898
rect 1078 2871 1079 2897
rect 1079 2871 1105 2897
rect 1105 2871 1106 2897
rect 1078 2870 1106 2871
rect 1750 2870 1778 2898
rect 1022 2814 1050 2842
rect 1414 2814 1442 2842
rect 1061 2757 1089 2758
rect 1061 2731 1062 2757
rect 1062 2731 1088 2757
rect 1088 2731 1089 2757
rect 1061 2730 1089 2731
rect 1113 2757 1141 2758
rect 1113 2731 1114 2757
rect 1114 2731 1140 2757
rect 1140 2731 1141 2757
rect 1113 2730 1141 2731
rect 1165 2757 1193 2758
rect 1165 2731 1166 2757
rect 1166 2731 1192 2757
rect 1192 2731 1193 2757
rect 1165 2730 1193 2731
rect 1694 2590 1722 2618
rect 1526 2561 1554 2562
rect 1526 2535 1527 2561
rect 1527 2535 1553 2561
rect 1553 2535 1554 2561
rect 1526 2534 1554 2535
rect 1516 2365 1544 2366
rect 1516 2339 1517 2365
rect 1517 2339 1543 2365
rect 1543 2339 1544 2365
rect 1516 2338 1544 2339
rect 1568 2365 1596 2366
rect 1568 2339 1569 2365
rect 1569 2339 1595 2365
rect 1595 2339 1596 2365
rect 1568 2338 1596 2339
rect 1620 2365 1648 2366
rect 1620 2339 1621 2365
rect 1621 2339 1647 2365
rect 1647 2339 1648 2365
rect 1620 2338 1648 2339
rect 1061 1973 1089 1974
rect 1061 1947 1062 1973
rect 1062 1947 1088 1973
rect 1088 1947 1089 1973
rect 1061 1946 1089 1947
rect 1113 1973 1141 1974
rect 1113 1947 1114 1973
rect 1114 1947 1140 1973
rect 1140 1947 1141 1973
rect 1113 1946 1141 1947
rect 1165 1973 1193 1974
rect 1165 1947 1166 1973
rect 1166 1947 1192 1973
rect 1192 1947 1193 1973
rect 1165 1946 1193 1947
rect 1971 2757 1999 2758
rect 1971 2731 1972 2757
rect 1972 2731 1998 2757
rect 1998 2731 1999 2757
rect 1971 2730 1999 2731
rect 2023 2757 2051 2758
rect 2023 2731 2024 2757
rect 2024 2731 2050 2757
rect 2050 2731 2051 2757
rect 2023 2730 2051 2731
rect 2075 2757 2103 2758
rect 2075 2731 2076 2757
rect 2076 2731 2102 2757
rect 2102 2731 2103 2757
rect 2075 2730 2103 2731
rect 1806 2561 1834 2562
rect 1806 2535 1807 2561
rect 1807 2535 1833 2561
rect 1833 2535 1834 2561
rect 1806 2534 1834 2535
rect 1974 2561 2002 2562
rect 1974 2535 1975 2561
rect 1975 2535 2001 2561
rect 2001 2535 2002 2561
rect 1974 2534 2002 2535
rect 2086 2561 2114 2562
rect 2086 2535 2087 2561
rect 2087 2535 2113 2561
rect 2113 2535 2114 2561
rect 2086 2534 2114 2535
rect 1862 2254 1890 2282
rect 2198 2841 2226 2842
rect 2198 2815 2199 2841
rect 2199 2815 2225 2841
rect 2225 2815 2226 2841
rect 2198 2814 2226 2815
rect 3430 3009 3458 3010
rect 3430 2983 3431 3009
rect 3431 2983 3457 3009
rect 3457 2983 3458 3009
rect 3430 2982 3458 2983
rect 4246 3149 4274 3150
rect 4246 3123 4247 3149
rect 4247 3123 4273 3149
rect 4273 3123 4274 3149
rect 4246 3122 4274 3123
rect 4298 3149 4326 3150
rect 4298 3123 4299 3149
rect 4299 3123 4325 3149
rect 4325 3123 4326 3149
rect 4298 3122 4326 3123
rect 4350 3149 4378 3150
rect 4350 3123 4351 3149
rect 4351 3123 4377 3149
rect 4377 3123 4378 3149
rect 4350 3122 4378 3123
rect 3710 2982 3738 3010
rect 2366 2870 2394 2898
rect 2310 2478 2338 2506
rect 2086 2198 2114 2226
rect 1750 2086 1778 2114
rect 2142 2254 2170 2282
rect 2030 2113 2058 2114
rect 2030 2087 2031 2113
rect 2031 2087 2057 2113
rect 2057 2087 2058 2113
rect 2030 2086 2058 2087
rect 2198 2113 2226 2114
rect 2198 2087 2199 2113
rect 2199 2087 2225 2113
rect 2225 2087 2226 2113
rect 2198 2086 2226 2087
rect 1971 1973 1999 1974
rect 1971 1947 1972 1973
rect 1972 1947 1998 1973
rect 1998 1947 1999 1973
rect 1971 1946 1999 1947
rect 2023 1973 2051 1974
rect 2023 1947 2024 1973
rect 2024 1947 2050 1973
rect 2050 1947 2051 1973
rect 2023 1946 2051 1947
rect 2075 1973 2103 1974
rect 2075 1947 2076 1973
rect 2076 1947 2102 1973
rect 2102 1947 2103 1973
rect 2075 1946 2103 1947
rect 2478 2534 2506 2562
rect 2422 2478 2450 2506
rect 2426 2365 2454 2366
rect 2426 2339 2427 2365
rect 2427 2339 2453 2365
rect 2453 2339 2454 2365
rect 2426 2338 2454 2339
rect 2478 2365 2506 2366
rect 2478 2339 2479 2365
rect 2479 2339 2505 2365
rect 2505 2339 2506 2365
rect 2478 2338 2506 2339
rect 2530 2365 2558 2366
rect 2530 2339 2531 2365
rect 2531 2339 2557 2365
rect 2557 2339 2558 2365
rect 2530 2338 2558 2339
rect 2366 2254 2394 2282
rect 2422 2225 2450 2226
rect 2422 2199 2423 2225
rect 2423 2199 2449 2225
rect 2449 2199 2450 2225
rect 2422 2198 2450 2199
rect 2310 1806 2338 1834
rect 966 1246 994 1274
rect 1022 1721 1050 1722
rect 1022 1695 1023 1721
rect 1023 1695 1049 1721
rect 1049 1695 1050 1721
rect 1022 1694 1050 1695
rect 2366 2142 2394 2170
rect 1516 1581 1544 1582
rect 1516 1555 1517 1581
rect 1517 1555 1543 1581
rect 1543 1555 1544 1581
rect 1516 1554 1544 1555
rect 1568 1581 1596 1582
rect 1568 1555 1569 1581
rect 1569 1555 1595 1581
rect 1595 1555 1596 1581
rect 1568 1554 1596 1555
rect 1620 1581 1648 1582
rect 1620 1555 1621 1581
rect 1621 1555 1647 1581
rect 1647 1555 1648 1581
rect 1620 1554 1648 1555
rect 2881 2757 2909 2758
rect 2881 2731 2882 2757
rect 2882 2731 2908 2757
rect 2908 2731 2909 2757
rect 2881 2730 2909 2731
rect 2933 2757 2961 2758
rect 2933 2731 2934 2757
rect 2934 2731 2960 2757
rect 2960 2731 2961 2757
rect 2933 2730 2961 2731
rect 2985 2757 3013 2758
rect 2985 2731 2986 2757
rect 2986 2731 3012 2757
rect 3012 2731 3013 2757
rect 2985 2730 3013 2731
rect 3791 2757 3819 2758
rect 3791 2731 3792 2757
rect 3792 2731 3818 2757
rect 3818 2731 3819 2757
rect 3791 2730 3819 2731
rect 3843 2757 3871 2758
rect 3843 2731 3844 2757
rect 3844 2731 3870 2757
rect 3870 2731 3871 2757
rect 3843 2730 3871 2731
rect 3895 2757 3923 2758
rect 3895 2731 3896 2757
rect 3896 2731 3922 2757
rect 3922 2731 3923 2757
rect 3895 2730 3923 2731
rect 3336 2365 3364 2366
rect 3336 2339 3337 2365
rect 3337 2339 3363 2365
rect 3363 2339 3364 2365
rect 3336 2338 3364 2339
rect 3388 2365 3416 2366
rect 3388 2339 3389 2365
rect 3389 2339 3415 2365
rect 3415 2339 3416 2365
rect 3388 2338 3416 2339
rect 3440 2365 3468 2366
rect 3440 2339 3441 2365
rect 3441 2339 3467 2365
rect 3467 2339 3468 2365
rect 3440 2338 3468 2339
rect 4246 2365 4274 2366
rect 4246 2339 4247 2365
rect 4247 2339 4273 2365
rect 4273 2339 4274 2365
rect 4246 2338 4274 2339
rect 4298 2365 4326 2366
rect 4298 2339 4299 2365
rect 4299 2339 4325 2365
rect 4325 2339 4326 2365
rect 4298 2338 4326 2339
rect 4350 2365 4378 2366
rect 4350 2339 4351 2365
rect 4351 2339 4377 2365
rect 4377 2339 4378 2365
rect 4350 2338 4378 2339
rect 3486 2142 3514 2170
rect 3934 2169 3962 2170
rect 3934 2143 3935 2169
rect 3935 2143 3961 2169
rect 3961 2143 3962 2169
rect 3934 2142 3962 2143
rect 2814 2086 2842 2114
rect 2881 1973 2909 1974
rect 2881 1947 2882 1973
rect 2882 1947 2908 1973
rect 2908 1947 2909 1973
rect 2881 1946 2909 1947
rect 2933 1973 2961 1974
rect 2933 1947 2934 1973
rect 2934 1947 2960 1973
rect 2960 1947 2961 1973
rect 2933 1946 2961 1947
rect 2985 1973 3013 1974
rect 2985 1947 2986 1973
rect 2986 1947 3012 1973
rect 3012 1947 3013 1973
rect 2985 1946 3013 1947
rect 3791 1973 3819 1974
rect 3791 1947 3792 1973
rect 3792 1947 3818 1973
rect 3818 1947 3819 1973
rect 3791 1946 3819 1947
rect 3843 1973 3871 1974
rect 3843 1947 3844 1973
rect 3844 1947 3870 1973
rect 3870 1947 3871 1973
rect 3843 1946 3871 1947
rect 3895 1973 3923 1974
rect 3895 1947 3896 1973
rect 3896 1947 3922 1973
rect 3922 1947 3923 1973
rect 3895 1946 3923 1947
rect 2870 1833 2898 1834
rect 2870 1807 2871 1833
rect 2871 1807 2897 1833
rect 2897 1807 2898 1833
rect 2870 1806 2898 1807
rect 2422 1721 2450 1722
rect 2422 1695 2423 1721
rect 2423 1695 2449 1721
rect 2449 1695 2450 1721
rect 2422 1694 2450 1695
rect 3542 1721 3570 1722
rect 3542 1695 3543 1721
rect 3543 1695 3569 1721
rect 3569 1695 3570 1721
rect 3542 1694 3570 1695
rect 3878 1721 3906 1722
rect 3878 1695 3879 1721
rect 3879 1695 3905 1721
rect 3905 1695 3906 1721
rect 3878 1694 3906 1695
rect 2426 1581 2454 1582
rect 2426 1555 2427 1581
rect 2427 1555 2453 1581
rect 2453 1555 2454 1581
rect 2426 1554 2454 1555
rect 2478 1581 2506 1582
rect 2478 1555 2479 1581
rect 2479 1555 2505 1581
rect 2505 1555 2506 1581
rect 2478 1554 2506 1555
rect 2530 1581 2558 1582
rect 2530 1555 2531 1581
rect 2531 1555 2557 1581
rect 2557 1555 2558 1581
rect 2530 1554 2558 1555
rect 3336 1581 3364 1582
rect 3336 1555 3337 1581
rect 3337 1555 3363 1581
rect 3363 1555 3364 1581
rect 3336 1554 3364 1555
rect 3388 1581 3416 1582
rect 3388 1555 3389 1581
rect 3389 1555 3415 1581
rect 3415 1555 3416 1581
rect 3388 1554 3416 1555
rect 3440 1581 3468 1582
rect 3440 1555 3441 1581
rect 3441 1555 3467 1581
rect 3467 1555 3468 1581
rect 3440 1554 3468 1555
rect 4246 1581 4274 1582
rect 4246 1555 4247 1581
rect 4247 1555 4273 1581
rect 4273 1555 4274 1581
rect 4246 1554 4274 1555
rect 4298 1581 4326 1582
rect 4298 1555 4299 1581
rect 4299 1555 4325 1581
rect 4325 1555 4326 1581
rect 4298 1554 4326 1555
rect 4350 1581 4378 1582
rect 4350 1555 4351 1581
rect 4351 1555 4377 1581
rect 4377 1555 4378 1581
rect 4350 1554 4378 1555
<< metal3 >>
rect 0 3738 400 3752
rect 0 3710 966 3738
rect 994 3710 999 3738
rect 0 3696 400 3710
rect 1511 3122 1516 3150
rect 1544 3122 1568 3150
rect 1596 3122 1620 3150
rect 1648 3122 1653 3150
rect 2421 3122 2426 3150
rect 2454 3122 2478 3150
rect 2506 3122 2530 3150
rect 2558 3122 2563 3150
rect 3331 3122 3336 3150
rect 3364 3122 3388 3150
rect 3416 3122 3440 3150
rect 3468 3122 3473 3150
rect 4241 3122 4246 3150
rect 4274 3122 4298 3150
rect 4326 3122 4350 3150
rect 4378 3122 4383 3150
rect 3425 2982 3430 3010
rect 3458 2982 3710 3010
rect 3738 2982 3743 3010
rect 1073 2870 1078 2898
rect 1106 2870 1750 2898
rect 1778 2870 1783 2898
rect 2361 2870 2366 2898
rect 2394 2870 2399 2898
rect 1017 2814 1022 2842
rect 1050 2814 1330 2842
rect 1409 2814 1414 2842
rect 1442 2814 2198 2842
rect 2226 2814 2231 2842
rect 1056 2730 1061 2758
rect 1089 2730 1113 2758
rect 1141 2730 1165 2758
rect 1193 2730 1198 2758
rect 1302 2618 1330 2814
rect 1966 2730 1971 2758
rect 1999 2730 2023 2758
rect 2051 2730 2075 2758
rect 2103 2730 2108 2758
rect 2366 2618 2394 2870
rect 2876 2730 2881 2758
rect 2909 2730 2933 2758
rect 2961 2730 2985 2758
rect 3013 2730 3018 2758
rect 3786 2730 3791 2758
rect 3819 2730 3843 2758
rect 3871 2730 3895 2758
rect 3923 2730 3928 2758
rect 1302 2590 1694 2618
rect 1722 2590 2394 2618
rect 1974 2562 2002 2590
rect 1521 2534 1526 2562
rect 1554 2534 1806 2562
rect 1834 2534 1839 2562
rect 1969 2534 1974 2562
rect 2002 2534 2007 2562
rect 2081 2534 2086 2562
rect 2114 2534 2478 2562
rect 2506 2534 2511 2562
rect 2305 2478 2310 2506
rect 2338 2478 2422 2506
rect 2450 2478 2455 2506
rect 1511 2338 1516 2366
rect 1544 2338 1568 2366
rect 1596 2338 1620 2366
rect 1648 2338 1653 2366
rect 2421 2338 2426 2366
rect 2454 2338 2478 2366
rect 2506 2338 2530 2366
rect 2558 2338 2563 2366
rect 3331 2338 3336 2366
rect 3364 2338 3388 2366
rect 3416 2338 3440 2366
rect 3468 2338 3473 2366
rect 4241 2338 4246 2366
rect 4274 2338 4298 2366
rect 4326 2338 4350 2366
rect 4378 2338 4383 2366
rect 1857 2254 1862 2282
rect 1890 2254 2142 2282
rect 2170 2254 2366 2282
rect 2394 2254 2399 2282
rect 2081 2198 2086 2226
rect 2114 2198 2422 2226
rect 2450 2198 2455 2226
rect 2361 2142 2366 2170
rect 2394 2142 3486 2170
rect 3514 2142 3934 2170
rect 3962 2142 3967 2170
rect 1745 2086 1750 2114
rect 1778 2086 2030 2114
rect 2058 2086 2063 2114
rect 2193 2086 2198 2114
rect 2226 2086 2814 2114
rect 2842 2086 2847 2114
rect 1056 1946 1061 1974
rect 1089 1946 1113 1974
rect 1141 1946 1165 1974
rect 1193 1946 1198 1974
rect 1966 1946 1971 1974
rect 1999 1946 2023 1974
rect 2051 1946 2075 1974
rect 2103 1946 2108 1974
rect 2876 1946 2881 1974
rect 2909 1946 2933 1974
rect 2961 1946 2985 1974
rect 3013 1946 3018 1974
rect 3786 1946 3791 1974
rect 3819 1946 3843 1974
rect 3871 1946 3895 1974
rect 3923 1946 3928 1974
rect 2305 1806 2310 1834
rect 2338 1806 2870 1834
rect 2898 1806 2903 1834
rect 1017 1694 1022 1722
rect 1050 1694 2422 1722
rect 2450 1694 2455 1722
rect 3537 1694 3542 1722
rect 3570 1694 3878 1722
rect 3906 1694 3911 1722
rect 1511 1554 1516 1582
rect 1544 1554 1568 1582
rect 1596 1554 1620 1582
rect 1648 1554 1653 1582
rect 2421 1554 2426 1582
rect 2454 1554 2478 1582
rect 2506 1554 2530 1582
rect 2558 1554 2563 1582
rect 3331 1554 3336 1582
rect 3364 1554 3388 1582
rect 3416 1554 3440 1582
rect 3468 1554 3473 1582
rect 4241 1554 4246 1582
rect 4274 1554 4298 1582
rect 4326 1554 4350 1582
rect 4378 1554 4383 1582
rect 0 1274 400 1288
rect 0 1246 966 1274
rect 994 1246 999 1274
rect 0 1232 400 1246
<< via3 >>
rect 1516 3122 1544 3150
rect 1568 3122 1596 3150
rect 1620 3122 1648 3150
rect 2426 3122 2454 3150
rect 2478 3122 2506 3150
rect 2530 3122 2558 3150
rect 3336 3122 3364 3150
rect 3388 3122 3416 3150
rect 3440 3122 3468 3150
rect 4246 3122 4274 3150
rect 4298 3122 4326 3150
rect 4350 3122 4378 3150
rect 1061 2730 1089 2758
rect 1113 2730 1141 2758
rect 1165 2730 1193 2758
rect 1971 2730 1999 2758
rect 2023 2730 2051 2758
rect 2075 2730 2103 2758
rect 2881 2730 2909 2758
rect 2933 2730 2961 2758
rect 2985 2730 3013 2758
rect 3791 2730 3819 2758
rect 3843 2730 3871 2758
rect 3895 2730 3923 2758
rect 1516 2338 1544 2366
rect 1568 2338 1596 2366
rect 1620 2338 1648 2366
rect 2426 2338 2454 2366
rect 2478 2338 2506 2366
rect 2530 2338 2558 2366
rect 3336 2338 3364 2366
rect 3388 2338 3416 2366
rect 3440 2338 3468 2366
rect 4246 2338 4274 2366
rect 4298 2338 4326 2366
rect 4350 2338 4378 2366
rect 1061 1946 1089 1974
rect 1113 1946 1141 1974
rect 1165 1946 1193 1974
rect 1971 1946 1999 1974
rect 2023 1946 2051 1974
rect 2075 1946 2103 1974
rect 2881 1946 2909 1974
rect 2933 1946 2961 1974
rect 2985 1946 3013 1974
rect 3791 1946 3819 1974
rect 3843 1946 3871 1974
rect 3895 1946 3923 1974
rect 1516 1554 1544 1582
rect 1568 1554 1596 1582
rect 1620 1554 1648 1582
rect 2426 1554 2454 1582
rect 2478 1554 2506 1582
rect 2530 1554 2558 1582
rect 3336 1554 3364 1582
rect 3388 1554 3416 1582
rect 3440 1554 3468 1582
rect 4246 1554 4274 1582
rect 4298 1554 4326 1582
rect 4350 1554 4378 1582
<< metal4 >>
rect 1047 2758 1207 3166
rect 1047 2730 1061 2758
rect 1089 2730 1113 2758
rect 1141 2730 1165 2758
rect 1193 2730 1207 2758
rect 1047 1974 1207 2730
rect 1047 1946 1061 1974
rect 1089 1946 1113 1974
rect 1141 1946 1165 1974
rect 1193 1946 1207 1974
rect 1047 1538 1207 1946
rect 1502 3150 1662 3166
rect 1502 3122 1516 3150
rect 1544 3122 1568 3150
rect 1596 3122 1620 3150
rect 1648 3122 1662 3150
rect 1502 2366 1662 3122
rect 1502 2338 1516 2366
rect 1544 2338 1568 2366
rect 1596 2338 1620 2366
rect 1648 2338 1662 2366
rect 1502 1582 1662 2338
rect 1502 1554 1516 1582
rect 1544 1554 1568 1582
rect 1596 1554 1620 1582
rect 1648 1554 1662 1582
rect 1502 1538 1662 1554
rect 1957 2758 2117 3166
rect 1957 2730 1971 2758
rect 1999 2730 2023 2758
rect 2051 2730 2075 2758
rect 2103 2730 2117 2758
rect 1957 1974 2117 2730
rect 1957 1946 1971 1974
rect 1999 1946 2023 1974
rect 2051 1946 2075 1974
rect 2103 1946 2117 1974
rect 1957 1538 2117 1946
rect 2412 3150 2572 3166
rect 2412 3122 2426 3150
rect 2454 3122 2478 3150
rect 2506 3122 2530 3150
rect 2558 3122 2572 3150
rect 2412 2366 2572 3122
rect 2412 2338 2426 2366
rect 2454 2338 2478 2366
rect 2506 2338 2530 2366
rect 2558 2338 2572 2366
rect 2412 1582 2572 2338
rect 2412 1554 2426 1582
rect 2454 1554 2478 1582
rect 2506 1554 2530 1582
rect 2558 1554 2572 1582
rect 2412 1538 2572 1554
rect 2867 2758 3027 3166
rect 2867 2730 2881 2758
rect 2909 2730 2933 2758
rect 2961 2730 2985 2758
rect 3013 2730 3027 2758
rect 2867 1974 3027 2730
rect 2867 1946 2881 1974
rect 2909 1946 2933 1974
rect 2961 1946 2985 1974
rect 3013 1946 3027 1974
rect 2867 1538 3027 1946
rect 3322 3150 3482 3166
rect 3322 3122 3336 3150
rect 3364 3122 3388 3150
rect 3416 3122 3440 3150
rect 3468 3122 3482 3150
rect 3322 2366 3482 3122
rect 3322 2338 3336 2366
rect 3364 2338 3388 2366
rect 3416 2338 3440 2366
rect 3468 2338 3482 2366
rect 3322 1582 3482 2338
rect 3322 1554 3336 1582
rect 3364 1554 3388 1582
rect 3416 1554 3440 1582
rect 3468 1554 3482 1582
rect 3322 1538 3482 1554
rect 3777 2758 3937 3166
rect 3777 2730 3791 2758
rect 3819 2730 3843 2758
rect 3871 2730 3895 2758
rect 3923 2730 3937 2758
rect 3777 1974 3937 2730
rect 3777 1946 3791 1974
rect 3819 1946 3843 1974
rect 3871 1946 3895 1974
rect 3923 1946 3937 1974
rect 3777 1538 3937 1946
rect 4232 3150 4392 3166
rect 4232 3122 4246 3150
rect 4274 3122 4298 3150
rect 4326 3122 4350 3150
rect 4378 3122 4392 3150
rect 4232 2366 4392 3122
rect 4232 2338 4246 2366
rect 4274 2338 4298 2366
rect 4326 2338 4350 2366
rect 4378 2338 4392 2366
rect 4232 1582 4392 2338
rect 4232 1554 4246 1582
rect 4274 1554 4298 1582
rect 4326 1554 4350 1582
rect 4378 1554 4392 1582
rect 4232 1538 4392 1554
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 3920 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1669390400
transform 1 0 2408 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1669390400
transform -1 0 3920 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2 Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 784 0 1 1568
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20
timestamp 1669390400
transform 1 0 1792 0 1 1568
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29
timestamp 1669390400
transform 1 0 2296 0 1 1568
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33
timestamp 1669390400
transform 1 0 2520 0 1 1568
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37 Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 2744 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54
timestamp 1669390400
transform 1 0 3696 0 1 1568
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58 Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 3920 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62
timestamp 1669390400
transform 1 0 4144 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_2
timestamp 1669390400
transform 1 0 784 0 -1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_17
timestamp 1669390400
transform 1 0 1624 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_29
timestamp 1669390400
transform 1 0 2296 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_56
timestamp 1669390400
transform 1 0 3808 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_60
timestamp 1669390400
transform 1 0 4032 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_62
timestamp 1669390400
transform 1 0 4144 0 -1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_2
timestamp 1669390400
transform 1 0 784 0 1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_17
timestamp 1669390400
transform 1 0 1624 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_27
timestamp 1669390400
transform 1 0 2184 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_33
timestamp 1669390400
transform 1 0 2520 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_37 Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 2744 0 1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_53 Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 3640 0 1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_61
timestamp 1669390400
transform 1 0 4088 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_2
timestamp 1669390400
transform 1 0 784 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_4
timestamp 1669390400
transform 1 0 896 0 -1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_9
timestamp 1669390400
transform 1 0 1176 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_25
timestamp 1669390400
transform 1 0 2072 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_34
timestamp 1669390400
transform 1 0 2576 0 -1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_37
timestamp 1669390400
transform 1 0 2744 0 -1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_52
timestamp 1669390400
transform 1 0 3584 0 -1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_60
timestamp 1669390400
transform 1 0 4032 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_62
timestamp 1669390400
transform 1 0 4144 0 -1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_0 Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 672 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_1
timestamp 1669390400
transform -1 0 4312 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_2
timestamp 1669390400
transform 1 0 672 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_3
timestamp 1669390400
transform -1 0 4312 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_4
timestamp 1669390400
transform 1 0 672 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_5
timestamp 1669390400
transform -1 0 4312 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_6
timestamp 1669390400
transform 1 0 672 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_7
timestamp 1669390400
transform -1 0 4312 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_8 Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 2632 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_9
timestamp 1669390400
transform 1 0 2632 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_10
timestamp 1669390400
transform 1 0 2632 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 952 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _3_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 1904 0 1 1568
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _4_
timestamp 1669390400
transform -1 0 2520 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _5_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 1848 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _6_
timestamp 1669390400
transform -1 0 2576 0 -1 3136
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _7_
timestamp 1669390400
transform -1 0 2184 0 1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  input1 Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 3808 0 -1 2352
box -43 -43 1443 435
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input2 Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 896 0 1 1568
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input3
timestamp 1669390400
transform -1 0 3696 0 1 1568
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output4 Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 1624 0 1 2352
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output5
timestamp 1669390400
transform -1 0 1624 0 -1 2352
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output6
timestamp 1669390400
transform 1 0 2800 0 -1 3136
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output7
timestamp 1669390400
transform -1 0 2072 0 -1 3136
box -43 -43 827 435
<< labels >>
flabel metal2 s 2464 0 2520 400 0 FreeSans 224 90 0 0 INmb
port 0 nsew signal input
flabel metal2 s 840 0 896 400 0 FreeSans 224 90 0 0 INpb
port 1 nsew signal input
flabel metal3 s 0 3696 400 3752 0 FreeSans 224 0 0 0 cmnmos
port 2 nsew signal tristate
flabel metal3 s 0 1232 400 1288 0 FreeSans 224 0 0 0 cmpmos
port 3 nsew signal tristate
flabel metal2 s 4088 0 4144 400 0 FreeSans 224 90 0 0 oe
port 4 nsew signal input
flabel metal2 s 3696 4600 3752 5000 0 FreeSans 224 90 0 0 onmos
port 5 nsew signal tristate
flabel metal2 s 1232 4600 1288 5000 0 FreeSans 224 90 0 0 opmos
port 6 nsew signal tristate
flabel metal4 s 1047 1538 1207 3166 0 FreeSans 640 90 0 0 vdd
port 7 nsew power bidirectional
flabel metal4 s 1957 1538 2117 3166 0 FreeSans 640 90 0 0 vdd
port 7 nsew power bidirectional
flabel metal4 s 2867 1538 3027 3166 0 FreeSans 640 90 0 0 vdd
port 7 nsew power bidirectional
flabel metal4 s 3777 1538 3937 3166 0 FreeSans 640 90 0 0 vdd
port 7 nsew power bidirectional
flabel metal4 s 1502 1538 1662 3166 0 FreeSans 640 90 0 0 vss
port 8 nsew ground bidirectional
flabel metal4 s 2412 1538 2572 3166 0 FreeSans 640 90 0 0 vss
port 8 nsew ground bidirectional
flabel metal4 s 3322 1538 3482 3166 0 FreeSans 640 90 0 0 vss
port 8 nsew ground bidirectional
flabel metal4 s 4232 1538 4392 3166 0 FreeSans 640 90 0 0 vss
port 8 nsew ground bidirectional
rlabel metal1 2492 2744 2492 2744 0 vdd
rlabel via1 2532 3136 2532 3136 0 vss
rlabel metal2 3500 2184 3500 2184 0 INmb
rlabel metal2 1036 1400 1036 1400 0 INpb
rlabel metal2 2380 2352 2380 2352 0 _0_
rlabel metal3 1904 2100 1904 2100 0 _1_
rlabel metal3 679 3724 679 3724 0 cmnmos
rlabel metal3 679 1260 679 1260 0 cmpmos
rlabel metal3 2296 2548 2296 2548 0 net1
rlabel metal3 1988 2576 1988 2576 0 net2
rlabel metal2 2436 2688 2436 2688 0 net3
rlabel metal3 1680 2548 1680 2548 0 net4
rlabel metal2 1428 2492 1428 2492 0 net5
rlabel metal3 2520 2100 2520 2100 0 net6
rlabel metal2 2268 2128 2268 2128 0 net7
rlabel metal2 3892 1400 3892 1400 0 oe
rlabel metal3 3584 2996 3584 2996 0 onmos
rlabel metal2 1344 2996 1344 2996 0 opmos
<< properties >>
string FIXED_BBOX 0 0 5000 5000
<< end >>
