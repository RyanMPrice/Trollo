magic
tech gf180mcuC
magscale 1 5
timestamp 1670260476
<< obsm1 >>
rect 672 1538 5400 4342
<< metal2 >>
rect 2968 5600 3024 6000
rect 2968 0 3024 400
<< obsm2 >>
rect 910 5570 2938 5600
rect 3054 5570 5386 5600
rect 910 430 5386 5570
rect 910 400 2938 430
rect 3054 400 5386 430
<< metal3 >>
rect 0 2968 400 3024
<< obsm3 >>
rect 400 3054 5391 4326
rect 430 2938 5391 3054
rect 400 1554 5391 2938
<< metal4 >>
rect 1173 1538 1333 4342
rect 1754 1538 1914 4342
rect 2335 1538 2495 4342
rect 2916 1538 3076 4342
rect 3497 1538 3657 4342
rect 4078 1538 4238 4342
rect 4659 1538 4819 4342
rect 5240 1538 5400 4342
<< labels >>
rlabel metal2 s 2968 0 3024 400 6 clk
port 1 nsew signal input
rlabel metal3 s 0 2968 400 3024 6 gate
port 2 nsew signal input
rlabel metal2 s 2968 5600 3024 6000 6 gclk
port 3 nsew signal output
rlabel metal4 s 1173 1538 1333 4342 6 vdd
port 4 nsew power bidirectional
rlabel metal4 s 2335 1538 2495 4342 6 vdd
port 4 nsew power bidirectional
rlabel metal4 s 3497 1538 3657 4342 6 vdd
port 4 nsew power bidirectional
rlabel metal4 s 4659 1538 4819 4342 6 vdd
port 4 nsew power bidirectional
rlabel metal4 s 1754 1538 1914 4342 6 vss
port 5 nsew ground bidirectional
rlabel metal4 s 2916 1538 3076 4342 6 vss
port 5 nsew ground bidirectional
rlabel metal4 s 4078 1538 4238 4342 6 vss
port 5 nsew ground bidirectional
rlabel metal4 s 5240 1538 5400 4342 6 vss
port 5 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 6000 6000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 106632
string GDS_FILE /mnt/c/Users/rmprice/Documents/Github/Trollo/openlane/user_clkgate/runs/22_12_05_10_13/results/signoff/clkgate.magic.gds
string GDS_START 68482
<< end >>

